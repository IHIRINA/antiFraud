PK                    $ > FIN_seed_148_int_414_head_4/data.pklFB: ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ccollections
OrderedDict
q )Rq(X   conv1.att_srcqctorch._utils
_rebuild_tensor_v2
q((X   storageqctorch
FloatStorage
qX   0qX   cuda:0qM tqQK KKM �q	M M K�q
�h )RqtqRqX   conv1.att_dstqh((hhX   1qX   cuda:0qM tqQK KKM �qM M K�q�h )RqtqRqX
   conv1.biasqh((hhX   2qX   cuda:0qM tqQK M �qK�q�h )RqtqRqX   conv1.lin.weightq h((hhX   3q!X   cuda:0q"J   tq#QK M M �q$M K�q%�h )Rq&tq'Rq(X   conv2.att_srcq)h((hhX   4q*X   cuda:0q+Ktq,QK KKK�q-KKK�q.�h )Rq/tq0Rq1X   conv2.att_dstq2h((hhX   5q3X   cuda:0q4Ktq5QK KKK�q6KKK�q7�h )Rq8tq9Rq:X
   conv2.biasq;h((hhX   6q<X   cuda:0q=Ktq>QK K�q?K�q@�h )RqAtqBRqCX   conv2.lin.weightqDh((hhX   7qEX   cuda:0qFM @tqGQK KM �qHM K�qI�h )RqJtqKRqLX   fc_out.weightqMh((hhX   8qNX   cuda:0qOK@tqPQK KK�qQKK�qR�h )RqStqTRqUX   fc_out.biasqVh((hhX   9qWX   cuda:0qXKtqYQK K�qZK�q[�h )Rq\tq]Rq^u}q_X	   _metadataq`h )Rqa(X    qb}qcX   versionqdKsX   conv1qe}qfhdKsX   conv1.aggr_moduleqg}qhhdKsX	   conv1.linqi}qjhdKsX   conv2qk}qlhdKsX   conv2.aggr_moduleqm}qnhdKsX	   conv2.linqo}qphdKsX   dropoutqq}qrhdKsX   fc_outqs}qthdKsusb.PKa_��  �  PK                    % 0 FIN_seed_148_int_414_head_4/byteorderFB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZlittlePK�=�      PK                    " * FIN_seed_148_int_414_head_4/data/0FB& ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�b�=O@�t{�=�{"�
]�=�F$��� �1^���Eƽ�曽��=�=J�=�>8�b�K� 5��a:}L����d<�	�=���=��=~,޽Y�9=�5O��+�</�u����=��>j�=�g�4-�=�c>�)��1I���>�c�<�,�����=��&�.�%=�������p_d=���2�Z�P�v��!(���J������޸�-|�<n;+=B��/�=��뽸劽ɿ��[����=H�=x�%�`����>:�=3��<#P={U�=��=��g����=�Ϫ=���=��¼�_*>a�$�D�]����.|�=��>y��=���=��뽋�=���<j������=O|�=��۽O��usѽ��8�7��vνݽ役���M ����=o�>\��=����ҽz���Wv>��v�NP�!�=���=�ڇ=��9�	>��%�MK=�w=��Q�� 5�;zo�<G&�:�8���	=y{=�~�=�!q=�PX��|�=O�1<����4��=�<L�U����>�m�ݜc������R=ci>F����%�	M�;����D��aE�=7T=z>pݱ=߂(�ů��E>��	��m`����$)�BY�٫.>"��<]̢�B$=��>�B�=�R'>?ᏽU�==,��a��X��=Qv���}6�$���1��5!�l>^ǽL���:h�Y���&�~��=ع�Ø�=>�\�������!>����p�<\=�۽��>W�=7E$���=cA��G+�M�^�Ľ6B�b�����$&�oڟ=�}�=Aj�"�K��5�<�v=rε���=����ͦ�<�W������Z���4��''>��<Чk=c=��4�;�v⻽�>{���:��ď�=.����t>���=v!��q��B߽ɴ�T>U2�=����]>Z�.<�uz<���<�U��ɥ�-g��m�d���f=�y>Nǽ[;>�0�:>D��<c��=J�*��,<k� ��*���#�����;R�x�;�(>��"�Bv��0����G>j=���<�(��т=3����|��ڡ����x���Ͻ����GW^�7��^�sq=�B�=15�=1%b�,(����t�'�f`�=�a>>�������x\������dJ<痰=|��S�g<R��KH�3�%����=	p����=L�ٽ�������=���=�����ǃ=+F�=�qս�nE�n�=a�>Zp�:�-)���i=��$>M�,=@�㽵��=h�=��м���=��=�ڽ�������_b��q<3��=s��7�>�>��<b��=���="$�R��� *
�]&>�z)�u|<u.�C�x���!>M�>n��<��ѽ��߽6
=U�o�r���#>�*�=����a��<�Ʌ�ʻ	>�D��?�<|'x�cWo��n(>�}�=���,T�=]3����t�:=�����=�b>��;/_��]��,����<[č=�ݵ�!�>]<�='�üY�=^�q=���>����{���47��=�f�=HG���>���=�6����=Q_�<�q��>���Y�>:����n<ȴ��4>˽�����C<����>?v��C<���8?�=�p��!;��R=[��=Tt�=%L��QYy��\�������C>v�=��ǽD��=���=��=���>�`;��Ž/Z�t�v<���<�?�dR�={�g<�߽(Q�<e<�=��=�0T=-|$��B�=�����ֽ
!�&�]= 8ѽ
�����)>�;9;S�>��=_k>���&���$�O:	�3B��Y�=6����k�K=��=���=\�h�7!>�t��n��=A �=�h�И!�&/��!/�<gT�<Jʧ��(��\�a��%�qRȽh���K=�>j���������^���"�=���=5U\�r����<���$@����P>D���>¼�s����>�K����=#�=�3�����
-���>� >ϸ�<���=��R�v�>�B7=���CY=Eeͽ�;! �=s8��m<��=pJ��A=~=Ϲ<4��=\��=�d>E8�=����μ�1y���[�X�߽�;:a�"Z���9<6*J=�D���8� ��ͽ L�=,>��T�=J�*=P�
�Ӹ����K�f>�D=S@���EY=zh�=�[ؽ����Ǒ�=�q�=6$��vo�=G��E̐=�]��_LĽ�X.�>}����=;E�����=�>�φ<�А�1>@�����=f���9�=?Zw=f�=�ݰ=�+̽R��=�>Z���1��Q�<������M�.9ὥ��#m�=+8d��[=&�>���}�Ͻ�g:=��n�������<��=<L"��Nz=|+=T3�=���_�=缐w>Eo�������>����T���0	���:�'=�Y6=W��7;����>�= @�=a6�F	ؽ�C�=O��T�;����*��=���<	��=du�=��]��f2�~>�&���b���f����R�?0�;�Vn=ࣷ=p�>��|=_TA�hvf=z>�̛��1���XO��'��:�̽D��=GB>�c<�b�=l=�>ga�<#{���s�=���_$	�+��c	)=[��R�=X7>�'����=~H#>3�A���[=�O�=r��<��<�!>=�8�%ێ��μAW�s#����J�>:6�����=�%>dn�7�̑��p�=5�`��~�=���=�j	�{{��-�=��>�A*�t	>|Ȓ=�V(��r>�lT<�+����Η���>|@����>�=Ը;j�=3�=���C�>O��|�����Y@�=$[$=�������=��=�Y�<�!�<�K��aʽ@�r=��>u.����,=��i=kl>1���Fn��U���ڣ�Br���쓼#F=<�ٽ�����=7��;?��=��'<P!�=�
Ž�W=������K��,4�=H�ͽ�x���Ʉ�9$��՞⽊�ּ��	��<-�/X���=5iz��;��w�<�c�i�=1F�=d��=�<�=$̥=8Y�=���=�'�2�>��=4�
��=ܛ�=�=�z!>��;Y�����=��b��P��v�Z��M>n��P��<(&�������<�Q�ڽ:=[D�=�?;���>��=q{ѽ�'>*|>*� ����DO����=���={�=7>��p�z>�I�=��ӽ2\>��I�	��=�Ϳ�<4>Sf�g���߽��>}�۽�>!ֹ��r�<�>���=�eH=Ҥ3<p�=-һBr��Q�g=�)��i�>l�"�y6<���=k:>ף�<ն�<�1a=x�/:�����,�3Ӕ��]7>9>��U�����X=�{$�i���q��@�<�s���Of��^����=D�==Iν=�ὀ��=�h>�IM=Io�=�.<%�?����T$���=�Km��x�4�=LUj=]V�<t}ɼ�ɠ�1)��`>�ᴽ�x�=Q�>I�̽(B~�N޽��R=>Ǵ=��>������yt=�&���ۗ=��������=�O97
��=Z;,>����c�M�*���ә�<D��^�=�I}=&\½�R���	�;]�=���;�ڕ���6=-j����>q%������݋>l��u���v��k,V=jB>���;��y�󽾲����%������:=��)�P4���:��G�_g=��=��=�㽇��dr>�D����&>�!;�5�5�A<=�+���	����=X��=(1==���=�!=+�>��[�ӿb=�ʽ�=H�!���=��=�A)��ͺ=e� >c0�-��<��׽8�>�>7ʟ=���,
>Ԫ�<�F>��o��õ=��|��"��X>�P��6>�$�j�=���j~�=~2�=Ů����=�~
>�0��*���(=���˫A�W/�=�����e=����f��c���f�<��#�K��6������� t=��e�=I'޽PK�z�      PK                    " 0 FIN_seed_148_int_414_head_4/data/1FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ1)=�k=G���	�=w�2�?.r����;G�yB���<�6�=xy>�眽��Ƚ4܂=P@��N�=
���%������,�����L���m���	���>�>w ���Ϫ��C�=C5����&�8"���߽�T;�>���?Ӽ��;s��=�']=Y�����@2i=����=ك�4Q�=)�<џ>���!)p���=���N�>�U�=�� 8(��=�W=�"�=�����=��==cD��޷�����mz�=Èf=U�=�+��e1���=�^f@����R�=�_�Y(�<�AE="5���T�=/=�>�s,�5P=6�����齻>�M}=j��VA���f�=�?�]��=t����g�:���B�}���=�6Ž&��^�=��'=�D�=�N�a�=�d�=�4���v���	������[��>�Es=��F��>�?�� D�<�y�=��s<�==鼁2w=��<k~�]��m�=$�ߠƽ���>iw=��ν��<�>=<+=��5���}�j��
H�=��'U<<�>+W�<`�>��������+=ލY���>h�̽A��=[�=(���/S;�����=KG�=l��934>6H�=���=�̼R��_�=!�=���S�=�ܼ�W> U���9��CW=�f���Qr�'�7�$R>M�c=���)���� ����=����)�o�=�^�=nu�=l�*�#��m������
��<�w�;#V��4�<�R�=�=�)
�<7��Q�yd���>�=��Խ/(G=��=��>C_J=����>�~������v%�k��%�U==Ľ��=D��_�׼�=>oD�=��U=�(�<(��#7��=�nɽ6=�35r=�;='�H����f(�=�i���H=#҇�y� =�~="ܽ��K�  |=� >�^>�AY�j-�<��l=�)�=s� �k�=��c�6HŽ�����A����D�=����`�p�<<J��NW;zH�<�D��ʙ��4��=ɿ{��ѽ�O�=��=�b>w	���>&�:�=�9���n�=2���2�ڽ�>[��=A=��- >�2>�򼒈>�Xٽ��=�ӽWM��vH��%n=��н�Rսܦ����<�P���->�ih<��O�YZ��]<h�����-�c����8����<��"<h�>���H��
H�9��ٽI��<�n� Vļ�'�ܽɆ�� �<:����y����A�p����2����=�g=�W�o�<�U��� =��q���ѻ�Dý������"
=�؀=Ξ�<�.y=�L�����P#>���4�<�&/�@ �=�w�<�>���=ڜ=���>������^�ڼZ��;�s�<6Jw��I�m�=b{��>�
�.gພs뽲H��;��; 0>�a>\ҹ�}D=�}{���=��>⼠��=:>l���?��(j�Sj(=������a�:��>��=���=-��=(	�<�Z�=�C=���)ɽyX�=������;��kZ�=Oͽa�\�����=1�=��v�=3>LN�M;��
�=�ۏ�}��Jl<1 1�VvԽ)̽~����=\��Q��p�a���^�=M����<,�8���>LC=4r�˗<=�z��S�=E3�=r�m��=����7���ΰy=�]>���=���=uq>\ۢ�Ċ=z��=d���5V=)
�=�3-:y<��>�q��׈=�=�/��]>����,�=$�>>�Լ�V�2g=�s�=us�sO&=�L���%�=k��C�=�q<��,�O ٽ���|�=G��d��ԏF�]ȱ�B��<���,>�����=EB�<��=���%
ʽ��>�/�=�?>�s>���=����ݽN"�=����"9=0���vh���%��YG%���N<5[�R�ս{�>zn=�w�=�/����=	@�<���}��=�<�<�ˈ>]v�=h��U�=q���7�=�	��bE��[���<ՌF�uiE��b"��k���">���=�,Ͻ� |��%�=KB=�Zƽ��O��dJ��+�;��= v�='�=	��jC뽴&�D��n�>{��My~��-�=BU�=��ۯ�=n�>���<�ɽ�Y���y2X=�4=���V��{U>��Έa��M��;&%=������;f�=�P�$=2A5� t��T�=<�%�=b��<ǜ����>���|���͇���>�k�=�t�=�h=ܗ>s��=Z&Ž����� �=��r�ش�=%T��/> %���v�Xɉ�_�!>��\-�t�>��=zzս+�,�#L�<��*>2����S��{>ҧ�=y�:��=�
�=���=�<>B/��p��V�=<>�=���e�n=�թ��r�=f���罡�����Ѽ�)�ش½�`�=ϛ�=�X#�:�ϽH�<	��@�N+�=��
�k
>�����=�z׽*!�;�ӽ�8��{>��F�=_'��~�=�5�=Qa@�R���/�=vŀ=ia=<h�=P�8��]н|ƭ<4Gy�"N�=�,�=���=���<ق���?��A��]������&����0���B���/��=7��<w�=��>���=}%����ǽ�.���;ͽ�~!�2p>B�P=��>i�=<<�G2u=���=�x�n�=��ĽU2�H >(#>00��&q='"=���1q=��;�T�=O�����޽��?=)�7�MHT=|�bu�����Ya�= .�=D�<)�ڼ���<53ｲ�������n�=�}���t�=�0�=��=8佅�����=�'�k��=�>�U>�.�=F�	=ٛ</��%����>v`b=ɑ#���<d�=|�ü��>ΰ�=���f~=�SӼ*�=n�>���=3��<��潐[��q���T6k=���=@��=ִ���|3���0�=���=�=N�=�;S�W����=�5��t�=(1�*�<녝=�+>���n�*�*��q��;'���,�ͽ�i�<���C�|��e���	��뽻�O�Ek罽�T<��Y��M�e{�Kͽ�>�)�����=��>�N��f𼘴ͼ_��Gҁ�#e��E�>��=?^�;+\�<'��=����ҍB=���o[�=��ڽ�i=Mmb=P��ˇ������Y�=�\�=eA�=�.<>�x���=�#��K�;$���lֲ<!ɽu�:4������>����`�S(!��K���=p��=Չ���D�ǽ��<�1�<�0�=L��<�@��j��A�>�Ù���=��>��;9�<a��:N��u{��N>'-C����=ذ�� ��<�Ԙ=�; >� ������8��i�d��k�t=R�k�����<�����+�8ʽD�=z���X����lJ=�͢�POP��q�W^�=��=�}
���!��
Ҽ�_x��|3=搳=<�>�9�;ī�=,y��Z
=���M��=w�=�5����=��p=�۽��=󧫼�kM=#��=����o��(h�=\4j�K���N>,�q��g�=b�i�L��@j+=~�;E?N� �>��=ˑ�=�Ť�B�߼������>h��=hB:�� }���>?�Խ��y�p�=��ҽ��V<qP�=����m!>/�`���=Z1��1�x�r�B��>�LཥcW�0�м��e^�=��=�[����=�h=�ûa��=e+%�Q��=,=)9�=i�_=r�=�Z����=�q#�:(>�W�=yK>~�>�g�)��7>�V��;|��<@M=��<R��<��`��>X�&>�����=��='����=SS>���=��.=�s(�	�=���"z9��=V�oȽ$V�<�_<y��(�&=�E�<�ʯ�dE�;�/��1�	>~98��L=�e�=��J���ν��ϻ���;���_싽ə=������f��:='����*�=P������<I���)������ ,�PK�y      PK                    " 0 FIN_seed_148_int_414_head_4/data/2FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ,��:�;*EV�y�(; �ںL�<�O`;���;�8�8�J�����-��:xWZ;�s��Q�;LJ�:�To;h��;�g:����]:L�;��;��;;��X;,)�:�]f;�=e�:Jt83G�Jǔ���;ڸ�:�@;��,8���;�S�;3ax;�ۧ;��-:�ߝ:���:pd3���:t��;�!�7�;O:X;�m58��&<c�M:~��:�t<��J;��s�_�:��;�;���:�.;�pT:}�;J�u:�Dκ|N�;L6(;�uX;�♻�A�:B���l)���:��v�p��7�� ��g�:�Z�9'�;Mp$;�ܲ;m�7;����=��N��s��O3:�F'�yI����<;����Y};5Jd9�e9� ;�Y�:���;���:gY�;;��:
��;͞m:c�:/�$;	5�9�І;k��-A���);�C;�N�J�ʷ��*k�9��8�ri;5s�;\:�;��=:nu�y�:z�R:?aR:+/��Q�;�m�:P�;f�<�wՌ;L;���:j�E;e/���:h3�:!�.:b�J;$��;Q�:;rU�:��;j�k���$��(;u�M;�������Ni��.W3;Ks;���;F�M;�DS;ꪔ:��>;���;��:�r�:�%@�68n��:9�	:�sQ;@-�:ŭ�;�к�-;���:s�:��9��%;�6�;L�9�=��*�S;��Ǹ$/<��N:gѓ:ߤ�:���;�;:ٲ';i�Y;�HF�rb*������;)�;�ў;b�A:_\5;�:���:�C�;�ً; i�:pܚ9�]����	:�.�
t�;�е:��:�,;���9]�e:E;P;i���A��x.�:��/;h��7�6�:@h;��N:��:��:Z��;8��:��p9w\�;�RZ;l��;�g�;������;X�9+^K:�A�9nާ;���;��:� :΋;HK����	<L�繧o�:�4	;�\;mρ:L ;;J!�;�o:݇;�|�:[>%;�6[;�E�:�r�:>$5�˽6;�8;��9�6�;SQ(;@x5�L=�:5��;𧓺��t����;��P��;K/�:(�;�ţ;(�9;VkI:|��;��j:	��Jƾ:8�o�L�`;�y=;X�:9ފ;-�"����:�=;��� ��;8(��@ߞ:b��;�f�8�_y:{�;z,F�-�;|/�;a;?6�#��:;�l���i�!dT:li�:�sb8�r�;�wg;w<W{y9��F;#�7�F��:��R;W�:x<��b���P6;�jh���:�
�;�}H;&Y�;nW�;�ᬸpuѺY.;��g;�A9�KϺ���;d��;�mp���:�;];'n�5?�;�L���\w:���:�o�;��;D+�:��ܺ���:Ǎ;%{I;��;�D�;Am�U[;z�8;�z;n��:�g;R��:�7���;��c�.7�9��`;���i��){=9��;U�/;�9;�B;"�8;3�D;���:���9�?�:8 �;���8�9q�:-\�!�;�;���T<;Sl9�;,��9cH���;�Ǌ��;:n��:d�+;�w�[�)�x٧��;F�l;:i;@JǺ�%@;~E�;�u����Z:��99�8;���4�4;��<�Q�:�R;p�:�8�9��ú��;�ޤ:�	�;/�;�cw:�#�9bڌ;	*�;��-;S�d�W��;/_;,��:6�J�|Q;w�;4�;7d�����:� ;%�:�;���h9AW6:S�:�H};R۴��ʗ;ɸt;����ZF;�_;���^�:9պ�$�;�2���n;�ڲ:�В;"�l;׎�;�y]�;;^;Çw;��1;�A;ƣ�;����;^��:���U�����:�#�:��P9�J��:�:�<�F�N6_���9hc<�';J�u;�a� ��H���ٳ:!�$;�[;�z:u)�;7�l;xUm;.Z:�.N;�%;i�C:�(;N��:����:�X;;���;QY�;��I;;��;%��;�	�;���;�W�[��;J�;���/{�;���8�]B;�N�:J.;��;ۊ�;h�¹��;�;/E;?��:[{�7��:CE�;m��7;AC);_��;ID�;��9@��9���:w�;�^:�4;���:��:�-�:0�V;�:3z�:�;``���a�:�:�ڔ:L�Z:�:F�*;R�9P����d��/d!;�~;D����:+4f;�l�:���:�R�:b�:3��;��:C��;��<���;oD�:_��9�*��|:k�3;XCt;A�4;;z?;/���ڔ";W��;_�;p"�"jI�E�1;��:#�;5+;�7;dl�:p�;ñ�;tF>�?::�͛:F�;�JG;����.]����:��;�6<�.��;A�;+�L;1Z9Y��:��;�F{;�d�:��;m�;tg+:sȔ�G�|;�Yc�~����;7;��;�u�;*��:��K���7;�, ;�3��/�9۹/��9�l�:5�/;��ɺ�}:T;dh(��;��<b�<SA\9�(�"S:@�9�g�;��7�o�:&�����;��G�b��;�0!:hT,;���;I��:�A�:,�;���;ő-;㭼�LM�:(<�����壺���9�E!�T	6��.;���;��:ƍ�;ȸ�;���:�+Ⱥe�:��#; �Q���&:��:L�n;Z�I;����s:�������:��J;ds�;@j;ؠ�:�;\�;[7�:��^�	F�:]y�;٦;��:F�/;F5�;a3|��һ(d};E=��]p�:Ad�;�7^::�;��9$!;��9z���;�R;�]�:� e:��Ϲ)��:��;|�ɺΜ"�Z�:�[9�ƃ;ۨ���к~A=;A��:�/;5"�;�ͺ��	;�����:�
��gG�Lx;���;�C����:�E;�7G;�~����;��;�̚:��b;��:Hd����:$В;g4:]�;<�9�:(p�9�D;�bR;v|�;qP;��;a��:�Ԍ:�X�:��w9�w,;��:��:r�:C%�:��]����:�^:�q:��6;v�:;��:��:|�:@��:�&:;(&ֹ�5�:�=�;��$;U|�;��9��9'2;��':���;��ܺ����qb9P=:��L;���:�����S�;z���ɼM:H%f���ѹHc�8{7e:9|K;�m;֐��<�9X<p;q˗:���(�6�{}>�<1];sȟ;��P�z�/;�ꔻ���:��g;����B;�;���㿶:�/�;�W�:7m;4n�2��8K�;wE�:u;��O;�޴9��;���:�=�:�U=;�w;d�;�7;��f;O&-;��I;�A;�<̺�];3F^9jS�;���;s�;��?�N�:;/m<�D7;�W�;�ě�?h�;`B�:m�;�r�:��9�����@;�?	;��;Fs/:<W�;����a��:���:ۅ��Aľ5��:��&���:&�;�g;�Ҁ:�-,<��;�� ;J�:�d�:$po:��~;��~:���:����;� G:'�$;��ۺM��;��M;�Š�d&��_�:(62;�\:�����º�B�;U�<�a���;�kI:d�;Nk����: 맺�;/`�:ۭ�)�O��@:��y:��:��<;�=�;��;��>;����#;v��;�;X|�9:#T���:#�B;a�'�c�;,j��<�:�@;#;=��:@�:�Dx;Iw�:|�X;r�d;H
�:\�:;���9��:�s�;Pţ;0"�:�Dg��E�ZM:�=�;��b:�4]���;���;u�Ǻ6~/;�E;�w�;���F5;�e:	);�]���-;aQ6;���:��/;8az�kĖ;.茺��;�m9;3��;��q�җ�9�	;p�r;�ҧ:1�b9?f;��V:�y;Uxd;ٗ�j��9s�!;��%;�p1;|�Ӻ��?�ά)��O�;­ � n<��:�Lh�`p��������9T޺:�d�<
�e;#�:�T;��;��:���;1� ;��T9�^�:�칣q;�<;��7:�d�:�];� �91�p;>�;���;��(9�Ӗ;�K;�h#;/!;e�!;�<�x�9[���PK(���      PK                    " 0 FIN_seed_148_int_414_head_4/data/3FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZf�>=��;����<�7+�Z3�e���`��<-��; ��<b�1� ��;u}i=�������<o	���=���_ =e�ʼd0"�'�;�o �I �<�="#��s�]=�G�<�"^=���ۻ �Y�<T�<�V��Uc�B����Ӽ�W��d2=���<��2=�e���;�<'���*$�<��C�ld�����}h�Y�M=j����X=��<�ِ�%(p=����X=dT<=)�*�������-=V&�r�h�8�A<�Eh<��R�Q���D=�`��00��<C�W=�p<=Ӻ��	0��C��-C�s��<�=_<�sO�¤S����<W}����;u�=�\&��<���<��:=���0�P�мv�u;��E����;S�����*=�r��&Ke�/����<�}�<*��<�1h��ڹ���;�}=�ȹ�"`���c�3Ʊ<0�V��o%���o��Y=��*=��Q��V�q�_=c�H=f�/<?�/���#��ƺ�O���6]� �Kb=��e=��;��<�݀�J��;kZ�<rf#��(��+`3<�����<��*�^҈<��P �<uh�{�<N���e���ͻ�fo=�pn=ZFG==�j��꼞M����(U=�o�;
��<]̼ɽ��gr/��=4Sݼ�=�{H=�J�;=�o�c\�<qqԼ�旼4�<��b=��<Pc����P;��	�G�T=N�.;���<RN�g�ݼy�U��(�<�a<�r1=��.��E��H�^<�i<���Rt�<]����HU�s�;|^=��F��ic=)1=ʙT���=����U\N;=����`���]9����r�O�U<!a<��Y=�-=󿉼��D�b�Ӽ��4=�ٸ�y�D<�uW�#rX=HA�6d�=����_1B=@�.=�B�;��yl<d81���e=lcg;M�M=�v4=H}��=Ez$������h���-�?�9�lj�<�g���z<��!�giY� ��<8�<jߝ;,=�I�<�r�8���id�`/u�o�����_<�Y4=Ļ������kd;�\b��O|��lQ=��8=f�;��=���a)�b�$�)�Yi"�_U�)L���W��0���e=+0�v-�m�b�#hռ��H=�p:�%8<-��<�w�<��=J���?�;@���"�<�s=$=�<pmV=`�1=~��<�S����)�!�b���<��=�H+�2���Λ=tX=��<P�M=\���*��w�<�l�C#M=�[<�wI�f��q/=%�Z�T���f=��P�-6�<�fV=���^�`��:s�4=
Q��	��-�;(̲;�&)=5�T��Q7���c��KB:�R���)��ᚻ��J��������>�����<��=�V ���T=���;35�N�<%=)=�$="$����+��=U��F=I��<��!�$7�+�H�4%"=%ꪼG�0���=��ļ|j)�X�D�A�B<sͼ�㚼����8���V]�<1!�<�C=7��;�m�<7�=�ت;d����ϼjN�2�X�0<�<s��<�3��>����"=�7:�=�lI�Z�,<�
���K��W�<�L=�v=�j|<A��<�^a�_v_��E"=�=`X�[rM<ޔ���)=9 =��g���/��>=�
�A�<F$L=��c=��;���!�rR1:b�$�7���b?*��P=�CE�K(����<K�f=�F= =jk��v=��'��⤼K�ϼ�DL��W<±=��мrp;��<\|�Lm=�4�=�\<������ٖ���M=g�[�;��<L��;��ؼ�zļ,��<q�.<ߔ����;�/�˶j�����<��|5��9=�O�;�55=�b��u��޽��H<�Z=��<m
ڼ"I<���m:��e�����<ņ����Q=�G=�'�<�,�t���ϗ`=��<\��h"=��\��\��33���3�;={s<�M;=U�}�J�<��=L�>=;��;D���<t��f>==�)6�Η�<���<�w=�;=O��;|�k��@���e�{ԑ<�����#��J9�<��<�t<d��\�N�r�J�8]m���<�NT=�\t�ʰ==&�<�X߸��K=|����a���X��G�o�'O��g&=�d.= j2<-1��M��;��߼�]~=M��9�%=_�=���κ����Ĥ;�������<���;�TC��=��F��M��(��*
=��_=~��
�<�wؼ�]~<a�n=O�<���<�K���q<�?��}�=M�>��'L��3�=��:��˼����
��7�<�e�yTV�bcR<����(5=)�6=�������=���l��<eZ��(p=�=0 T=�1=�1�:O�-=_;���߼�Dd���K���)���)��0b�l(�e�廹��;OK�ݗ��3�<��W��Gv�i�<-x5<�,0=�h��+�a�<�=w�<?�9�C���x<8�'�ܺ����e��<�B�N���,;4��U�/�i;�K=p�˼,�%=��ϼ6Uμ�s=�G��d~5�.���i,=��@��=�=�j�<B|<<�2��'�%=���<���;�(���<-Q�<3�/�Dpf<w�<~/?<��j=z
��jGb;��(<�G�<LU�=�������~�O=��n��~h=o3=��=g��dᐻD0<� �;}�<MZ�)w�=��o����y�<�"=���%�<�V,�c#Q��TK=�(<�E���]�0+,�3�'�p��<N��<��/<��)<w]="�O��K	�&�A�%��<LD=���;O[���Ā=�=�c�^�˼gU2=��=�#m�x@p�!H��~�>�D= 6=wtH= �<FH�<��E<��X����<!B=�`=y`<m��<��(���<��ϼhG:]9�<u���ߘ�U��<��<��<1�;)P�lEȻ��B������Gl�����<�Iܻ��߼s5�<3pt��@=<+�=���<G�<�(k��K���̼$�=�:=sӻǢּ���ڗ[����<�;�Y�m=n�4���ȼ,�<� ���l����<�j=b�=�觺�~S=��6=��=O�]��2}=< =���<��������鵼�t$��'=�g��)E=��߻1B��eXF=�DC<vg/��P�V3��A8(=�ݚ�pF���=,k��<�<?��@ǻ+0��'=���<�^��u�<�+���)؛<�򻔥6=������:asS=I2��)���c4�U�;C�����|�<&E=h	�;k\�H�F=��z3=�,]�:h����H<�s���sOa���J=g�ջ�8�;~�D����<�UA=G{,�#]�Y�;�,漏�J����'L<ڪ�<6�������:�=A4u��=��Y=3��<��\����<�,�;B+=ٍ
=��d��p	=��Z�����=�*=�c	=M�<s-o=��� ��Hɿ��zX=�31=V�8�W���	g=��<d�����;�h�:�����T�Xz=A~��^V9=?��V�<�tl�܉�:��<�G�<ߦ��_S\�0�?=�xS�|.�<7l�<>[�<�	��h =����=Y(�;<<�)ܼ��<���-X!���ؼ������ �=��=��T��Br���j=�S=ȆK<��*=�*6=��\=Ij4���8=&�r=2��f@=�k<��=-�<�.����< ̻��<*z�<�~5=f��<ͫ���$�bDW��r��5A��U�)=%�㼩�e=G6=�R�F��<P�L<���;���eTJ��`3��b��K%=�?A���<I�<�S�⁧�t ���	�<�6�Lk�<�����c��=��(=���;`�k�׼�R3<��q��-C�4�.;ܡx:�an=�ֶ�Hr���(�\��;�𰼋��;c� =��O�-�P<ٞ�:���2GU�:<R�=��[<�;F�R=�>�9G4���<�4�xV&�b߮<
P���V�<T)6=pA㼤}�<�J�<���<DgҼ4�l��[仪m�G�=��D=��6=�#�"��;�i%<�m<���f����!=�P�<^su��=��7��.�!�	�5���>����<y�?=�#/<��<VI=A��<W�D=�
w��t�<�Z�=6;��;�"=��l�H�������%=�u;=��I��ɪ<�ۅ�/R�<�m�<8�l�Ｉ
E�U�4=;�<	kD���<Q==�q��,�"=p(P=Xy<G;��k������k�NQ=ܲ8=�<����L��<��=~w�-��<�^$<�O=<�a=�(=�6��-ܻ��S=��8=����>p��Zռ��k=> <(t~<��^=
��<�{�<�@;��"�;+��9��;�b�<��+=��<�&�<:���"R�S�;�>$�Љ��6΍<��w���=�	�����;H~�<h�Ȼ.��;oh=��V=� ��W"��+=_��X�=�| �5��7�<����<d;Y��o=�=��~<�#��X=���i6=W�;?Oi<2>=;�=2����}=�;����|<�ϒ��ts��E�<9k|<�) =E�&�+�";��,�OU��!����6��MZ��k�!-/<;�ɼ���凣�U�;�+Ȼt#=1�)9Wf
=���å��d��+U=f*�<���<��<ޞ�<d�O��׼k��<�[�;;�����<���;n�����f<,l��2"==M��G�<�U�<-�=�X���?�_u�OJ����`:l�=wiż�f��$=u��P�`�����Aˁ=�=��e�.���E�~��	���
��Cg;�\�<e����>:��E���<�#=��!�M�(;�	��� 6��Lz=��1���,=��><;\=W s<�5�< �:�}h
=f0;�n�;hY�Q�̻���L\�y��<��a� ��<��&�/��߉�d✼��,=.��D��<?�Ҽ���o�b���;=�`C<2�`���<��㼳^���f����������G':�<A����w��qs��a=vݼ�r��x���O[���2=���:�c;`�2��rY�܅V=�D�<ŷE�s�ܼ��Q���)=җ]�H���>=/�뼚? �7=Y[�<e�_�� �%��<7�����;��=��=��9��f��J�<T?h��*�bz;=�K@=~�Ӽ�9�iE�<�=J\������;?̈́=�Y<���f)�����I>=����:���<�`!��2�<�
�<�,�<A�ۼ%����;'�-�l/M=I�;A��<3�~�fl��r=a���_����5��fL�[����1-: �a�_˻��@=�ul=��J=`NK����;�꺼�m=�K:�r�o�b<�< �87�C�=̅I=�+2;���7�ud�<��d=۳=ոc=ޤ��ȟ��е��\,�<s���Z�3;SX�m��<�V� b�<6�f�U$O��pg�v� =���<�z1��;i=��<��[:�T]=��<o�^��C%�<�W�<�üh�<��%���[�/����� �<1�d�� �=���F���ϼ����j^F��߲�)��<2	�=%'<X�;c�y�S�<�.�ܢ=?���>�x�i=ļ��u��

�;@�<������<F�U�`�<��׼�ؑ=Y��<\Z�<ϔJ��q4;��T<�;�E=UC��,o߼�
=��]�I��Z-:\Z
=��<̩E���<�]�_7�<^9=ü�=D��<Xd�<n1���<*��<w~��6=�@=�̼�fs<���z/(����^i8�褼CO�:��;!�g=������C�y���iT<�U9���O��C��l�[��	[��U�;e>=�������+G�<X���DA����f�W=�ˀ����<UEB�*�%�Y�c;7��:��L<D�=��8��VF�q�~��(�U:N=��|���Q<4����l���z<�����=?R�"��7�A�� N�8�;=~zn=��>;韄=��/�X�:='д�u�x=�]`���n������;��i����<��<�$I����<�%6��==ٮr<� =�W =��H=g��<��M=�|���X�P+����<<Ġ<���<�a�)�X�L����$=�S=�k{�E�]���Q�n�ʺ�L=s�t����;�bŻޜ���f=�Ƈ<xJV=�=>掽��=�hZ������=NF<���=L�7���<��2���<�c=�"@=���<�E��`=�Q�G�%��=Rh��hQ<m��=[=�ō���;�������1��=.�P��|�<�%j=^_H<�>�\WӼ;���d:r<�K�qlc=:�J=7.�<G�=i�:�3�"���;�U<GAʼ|~=��9��﷼	\J=���<����4�<�F�^9>=����>u=�m<]�a��=��<^Ɉ=HK=��ʼ�����=�Y�;uK��+W��{�#�1�'����)腼Y=�,��ʈ2�����A=��)��=�<��`��[ :A�<}FH���X=h�Z�]�H=�<5*<����J=��>���<rtw������]���T=S�-���~<��;��O=5#����\=Mlb=��6��
=a�;`��<��I�٭;K�<���;z?Y<�fF�����:=*�N�߻h���-��\���<ˠN��G߼{�<<M�:=���<��㼎�g�֬<�d.�݇�;�&��I7<_�=���<�k���(=+8׼6�a=�%�H�<�eʼ�0�<��E=�6��O��<��J��D��~��<O��Ć4�k��<����[x<��˼a��<�����J=��?!6=��L<�*�#�;�)<���]b�a4�#XJ�YL�;�:$�EJ�9��G=�k>=D��<�M=���~�6=�N�=�mr<P�:˄�<�5D��؆;o4=�;%�"=�/=���=�=�j��A"���	=�؅���໳��R�=�����M=I������[<m��;�Y�<�,%<`�@���4<}p;�,X;*�D=><%��mF����<��:#�D<9���rԆ;�O!�����>��uQ8�
��`Q(��D#=.h��k|���}�o��<Jnr���2�m��C���wz<O�=�q=���
 =ID=��5=U�<�l���=([.���=$�=Ї_���f����=��7��1[<���;�u��V=�,w=8 c=�Ӵ��D/={V@<���<R�T�5����:��J=�ou�ғ����;ymb�w�<qO;?�~o�<p���:�<�~�<�=At_��#F�Kӕ=�y��Ԝ<��<җ=�m<���q�<0�D=O��J:���SU=�8�;�U���f���:�)��}�|=�R'����<ms��Z�k=Z������W��</p$=��?<h]���n�Փ�����Ȼc���<��A��ͼՋ�7ct=']�T��<2�6<HQ0���Q=��(<�|=M��<r�%<��̼�+j�},/��c(=	�P�/���ʼ�=3�D�N���31=�K��>΃<@�¼���=Y�j=O_��*�<�L�C��q �C�b�`��<�$<�'�{.�;p[@<�	U=�dȼ�����<%�;v�l��C�2V6�;��<n��#��wtҼ�%�<��U=�Q=��=�:{<2x=�)0�+�<�ߔ<��\<��;�mѼа�<�\��lӼ6�ټ}�LW==#'<�������"�=1�}<�T=����©=�����[߸<2nf�*i�$f��{��:�	\�5wǻD�<�̋<s��</-�<�7<\@';��O�X�e�����6Ӽu��^㳼�2��)�P��E2���}<'�Y<1v<�&9��J����.<������<�;��=����u4����<���<���6��R)=��<�}><�*T=���<�)^��@�����T��=��;�7］��<���:�ԣ<�w�<|�z����g�+�k58=�ui�>&8=<c�<�"<�=h)=d�*��h�<5[=��<�3=�ZE��Hk=7��<���<���;�))���e=r�ͯf<��H�L�<(�׼l�;\����c`=`E=lԳ<��6���"=B�����<X�
=��=_�<9��;��W���=��#<5�W��=I=/<�)<!���ɼCf��Ge���9���I��#�<KQ��#��?=��;|����,=�+0=�k��C���<����jF=6�:?���=-��;�%��9���<����2�)=��d-�����]d�9�Br<ܼ�:�"<�/=Ŧ&��=.)�<�^7�֐5��] ;K�N�{ϼ�t��<�q�;XS=9N��C���=�0��.;��;=4�;�b+����/6���Ӽ�ƍ<g� =0��;gEͼ�eݼ,�r�����"=�2�-P<KcK=Ub$=�D�<T;�	:w=Q�C���1<)�,��C=���<�Z<�y=́)=a!B�T �����:=�A��8n�֠=+	B:%~(;}$X=;�<��"�e(�<=��<H�L�D:=��Ѽ�tk=.�μVZ.=$$�����;�O���<�绶�����\=^kE=&�Ƽw~=���b<p.�]B�\�M�������^���=�T��wỂ<����I<��;�5Ļi@.=���;�;c��
;ڈܼwP�<�f)=�`�=��=��J=g?=Q�I�嶟�a=��;$�	<T=��ƼT���?���ļ*F��o����� =�K=TWF=�_I=#8=�u�f�2��U���5=�z<��B�<��x�.�<*��%V�<���5� ?��6���Ǽ�Ӽ�މ�")���μ`�5�	�=9q=��-=�¥�F�G:^9
�W�˼/��;X|L=���<,�*=ͧ�<�[<�3!<��<��Q=�����*�<�ټc�&;)N�<}�
�R��:���<�Q���G�<k����;=�8!��=�ػ _��'1=7[���ư<�dw<Q�<��h=�㻰7_�� �<-肼>�r<�L-��T]<�A_������x=4�k�5��;+g2���όd=D��<[��<�f������_:=K$B=��J�Cy#��}>=U�`<�I�:P��5`�%�7�B��F�!<U�/��<W��{vw�|=R<�<6=�<G=���<� �<��#=����=�b"�Ğ�<����
6���B<�a�9vҬ<t�=A�b�?�,=@0=miܼPo-�;o�<�<[���<��y<"7�'Q(=C	+=�i)=���<����<g;1BR���,�`k�;��{=嗁�q&�_�<��`�B�.��# =gbo��<�=��F<B�=���(��_��`h���w=� <r=-��{�\=׼Tf�����=�&�=�g=ǘ�;�[�<y�#=v��<T��k'(<�)=%�2Tļ�{<�x^�I�h�!4�<^�&<�ܔ�I�����<|X���I$<t�M<K�м(� ��<�;rfT=Z�0=g�!�E�<�7ۼ�$�<^��<6mg��c��RP��!`��m=12�;=�;WBa��h;!��`���� 	=)�6��>o=�yT=9눼��й�	���ǕF=H��M����r��q�=�_�;H�:��
�<i)�=����r�(=w��;� ��}�N����,����ո1=�X��Hֻ��I�����c�����=D:����2�3��<�}伹�<h�A=��I<,6Y�D�'�k��<l�g=��;A� =�<�<��!m��7b.�ΓZ<����<�= <�QM= y�<�[�*�=#�����S�Sg=������<��i���X=�ļR?��Ҏ^�><��u��5���x<|��<�<�\����</z����;�-:��@!�=��J�<�������9�=U=��<{=���<�
=����f	<-��<pu�^̵��I�{l�<�=��#���*=\(2=c���q��]��,�=~��<a.�;,��nba�F=�.�<�g;=�v�<j�<vFZ;�|"=�Cu=[/n=�=�܋;�|<W�ż���j�G=)�;��ؼ.F��07G<P���˥�;/G==��<�мˋ�< /=��:=�#=.��;|!���D��i�Mj6=y�=g칺�mR��\=`=�?=CG�i�L��}<o�˼��D=�{���o&��d5�U�:=Hꂼ����<�����d��s�:V�=+�t9}8=�<�m꼫�>�����m��eC��ME=_e�<��G��J��f=���<�oB=bit=�R��|�;�a���=����B�3�Ty=(�=�c�;��f���`	��H@��r���F;�4;�G����e<DVo�S�5���μs8�P�b�r-=䡆= �Ƽ=H����<�=��;�+�6�U�v�<J�;?�I=����h:[�6"B=<�/=.*���<��T<D㽼��2=Vj�<�=ļ,7��6��;���$ּ��7=C�/;��Y��-=}~D=V.��Ha��~��`=�u$��43=f	=����=�S��>����N�7����H9��9��k[��u<<U�;@L�;-&�;"zټp�<O]<�r��"� �ʹ���n�<��<d"�g�<FAq�E�"=&9�<�n�<b5O�}A)���"=��<-���� �<^��|�<��-���P=�?=m
Ѽ��w��R=~w�N8��`=G�f��mR<5}�;�i-�DlB�����'��ϼ����G6=�!H<=�=�~L=ܺ7�	E��M=���eot�M�q=g�����)R^���v���>U�p?=���4����'ъ<�_��l��9Żv!뼏���)⼤��<��� ���r��.�=%xռ"�`�=B�u�1v�:oD=�����x�;{[9�@R���=K6�<�����/����2!u�Jg=��<}{=c"�;�E�8�:=k �;0�߻k� ��;.�<��%=I%�<i`*= �Ko¼.&<�����=��<u�D=�ʲ<��2��\;�V���!j�˚ü!��:�M>���ּ�@m=Ȩb�*���8=eC@=�V|�����+��B��Ύp��	\�▏��~���(�<���<��;B$+�������<w���`;�\�<��<)��<��%<t(�ʍ���=���Y��U�ռ��<ޮ�+i�����r�;x��<�y�9RhJ�R8};<:o=� �;�iV��kI���<?'��z��+�Q���k�<����dx�<t4���I���;a��<�ۨ��`6=�MG=����:�|�<{b =���:r)=��R9��#=�lN<�4=[�]��:G3[=uF���4<�t=���óc��=K
ں{�=�)��2�,��ո���w=�&�<���<���|L�٦�ZႻ�<=d�<��m�򮵼g���a*,��}U�T�)�LE��'�<&<y�w��S�;L��()�#�a<��!=���<���;���,<	gx=�� =�Ş��Y���2��f9����<�s=��<��:� >=�]��I%;��<8=�.�<eB�9��w�RϜ<�<4KD��]��T���p[�b8=;*w=�C�S��<I4���M������};���q*=�K��V��>�=�=0�=��1=�i�<�\=c��'F=X�K���<��ȼ�rB��О�8��î�=��=�e5=yr[���9�?����l��X	��w�FC��w���E=+ �<%�[��Kټ��G�Wvɼ�������=�p=T/1=L�<�мQU�<��#<~��`I<s�)��w=����RH��"�<��L=gx���M��������<�߭�D���=����]��v�;���ʪ=�(�x/H���1<�:8PL�.�A��^���[�O	�;
×<:]%�b�A;(g߻�/x=�I�<}������<����/���<�|���#�,>ͼ_�6��m�@?�<X �<��I���=���h#=}�мQ��D'�>��tO=~�=���f�&=`��=�����1=�==;�MW�FII=���I���j�&��=ze=�a=�|7=`�!��?*=��.<<�f�ޣ��ڜ><|��<GѴ�+�żgI<00=̣,=��+�����S�R=>�&�{L�[@;��)�X�"���;y���N-=Y�=m��<��1<�=�o�;����I=�z�;?�<H
=��ڼ{sk��݃<��3�(=_u�/ ��I}�<hN�<;��G5�<6�H=(�D<ёp��z*=w��<��j��ն;�1�<�q2=��h�
�<Ҕ<�<-)�ay�<�(�;>����!�&p�<�4��=,�<���<3��
X=e��<�3=��O�K�
=14�<�?=���֝[;�H��B�;�6���<e��V�3EI��:A=j�;�{�	=l�<ݘ=�˧� }H�`�<Õ#����&�	�<=���<b�>=��˼��I<��漽U�< �c�3t=s�����[��<����ʻ�"�;f��;��:=��<[@��|<��D=xv�<��%�:�(�m�=�&��դ<�D�<��<�Q�[�:0��c�dwm�W=��)&A�O��<�W�<l�2���!��G_��7r;:�b=~��<��=�̜�<�!=W;��J�cO�<��%�[�����<����¹�U��I=�&`�� =��=	�u��H'=��˼�M���D=�IX<� <^�>�Lh�<�q�<Ⱥd<p=<e��Y��G=/�a=y� =S}�<
9D�ǭ�<�ZZ����+�^<�<�O&;��<�y)<S�<Fʄ=���P<R4�J` �ō0��fA<�Ě<�<��$=�+8�]��<~2ͻ�@���0=���<���;S[Ϻ{9=�==�X�=����@*=T�	�]I!=Y����"V�/`���["=R��<T<@x'���<�O����T�%"���M�|���_<R�"��1���[<b2��Ұ;Ӎ�<������,�;����2;[#�< �<�kA����kA =�ۻ1�ۼZ=`7���x=e��<U�=� �9Hw��J�<�.�id=J͘<識V����"�<�W
�u�h�%��iú�;�;�N;�O��C<A��<�X��(1�T/�@�\��X�<�<��;����^ƼfX	=�<H���a�?=4��g�4=^K;��ۻ��x�r�(=��=d��=B�b����<�Ӽ =��O��a߼ó����<"Rz=�4��1=*ۼ}�<�2.�����0�G�	����1=�6���)N��c�<�W�	�1=��=22:(�R:PV>=�M��m�z=w�ük�b��a��<-y_�w���T�<��<)s=e��kP=��Z�iR��ʻ��)=�`���YA��N=�b�;���=�⨼Y�ݻ�;��[=^���1=���=�m�<�2̼���a�<s��:}�<z�X=@��,5f���<����=��H�g��I��}<�L�{���Fa伡sμr�=�	=w|o<>��μ;4@��໣�N�j=��;�냽?� �I��ä�;�XH��d<[=�W�<�])=�����u�<�0$=�����6~��Ƽ�T3=9ܼ����=�ӖJ�޸/��g=^q�<����i�r�^=r/=��L�����	��Sq��GZ��=��� 0N=WOh��N=�̑���,<��]�u��,�<�z��<�D�=��`�H�^J�G�<��R_����<�H#<��D=��I=&}p<|�)=�v����=��̼Q�<nm+=����j�\���w=��<��":�^�<��<�R%�}�Q=v�B=�Q	=@��<"�;)7�qpQ�D<�Ԓ�<��-<<%��Ah��W�<�b�<)%�;��<wF=�	7�]��<�f=;�P=	(=Q01���:<-)`=C�<�Mt< �N��<����"r�=��#=>��<�=Л=��.=�"V=�CC��W�rGo<b�I�^�r<�ڪ<�=����3#<��U� ��<�=�`�<��<��7=���*G(==�P<M���\�1=��<�Z!=�I@�,�:�Y=-[�<�� =��G<R��<�XǼ�E=[/!;y�=i��<��g=� ��Rpx=+�ټ$N����<8ٌ<*��<8^P=��s��]A�H��<;�F=x*�X�M�(�<8��<���;׆�<��<y
 ��r#���7<�`<���h��<�@�O���9�;1NK���I�����;��;@ żU2B��mD���[�NyS=��L=�|9�t�û�]
=�҈<F=�
B=��8��e.�dۛ��Nǻ
��<�CF=;����<wu��aUe<��L;��R��
��)�<��H�S���<���<kك<�䋻@*��#��#ۼ�]O=���<?�>��T�;�F��q����<��:��4=5�i��5��W�	�l�k��><��F=1���0�ۼ4�e�$9i�hA_=�q=4<O�AA�<P��=�}�<��<�)���y:<I�=jQw=)?j=�]=��Y�^Z<�M�<�r�</V=��l���	���=C�
��PT=�Ѡ<y
��2+����-k=��@=�:=�Z���<M�8�`츻N�R�p��<�᪼���yV =[ �b�=��<I\���=�;6�Ɠ�:d���J�=��W�p�Y=�sz��}ٺ��E�bS=����*T�<��<|�-�
)+<%E�=�ў:WCu���;�+�����0e;%8�7�9��h�<i���=�O�o���\���< �e�Q"6�6�R��i*=9G��.��1��<��ѼR�;�-�=R�:�zZK=b�k;��<'脽Q�����м�\�<c�J�EPN<g�L=�%#=/�/;��n����<1�L�u�Yl��<�H���E�l�	<�4�JWY�� =���YL<9cU;n�=~y>��>;<�=�;	�C���;5�<�8�<u�<�B��Y��bi��"�Ub=�밼��<�&=m�Ẓ=��A =��Z=�d�	����B=ńF=������<~�Ļ]=����<$�,�	!=)ߕ��C��R=���<�g(�='%<�I=7Je;8>7=�ׅ�;~D=%�����E��8�^���-M:=�f�8𼧜e�wG<���
n�<�=��);�����j�?��\AC��?=��i=�P��!ȼk.6;t���v��r��x�U=���j1"=�~g=�O���>N�� (=]�X��b=$��:�i��\�&��1��;R��<C�W=�$L� kE=��ȼ�?̼�%���e=�V"�^�v;�q/=��=�;��=y,����k<C�<?�ݼɷF��M�=��T<�?'����<��<4� ��6��uX=�.)<]�Ǽ;Fq�\�<u+�^ּU��<��4�������:��^�Rӌ<�,�fcݼR�뼞��A�=��;Z���8=���;F��<t2�U�v�+Y=6]�}�kM�u=G%Q<����%�=��=s�<�x=:�;�*��o�8;�(�ej��?�<��H=7��<�c�<kQ"<��Լ6�9�`<��a�=y$=�-�;���;N�9=�=aF=�������N��
=��Z�l?�;(��<k.'=m_=1x��g�;R=C�p��^/<��a�%$����༜R�;�le��/��.';å�=m<��>�L=Ei��y=���e�����Z�Y=��=E��� =�߅;�jּP�̼'���S�?�|�<ӬV=G=�J�Dv
;~O=�����E�ʼ>ʸ<��<=�K��T=�	��{}���e=��x=rIl����<�(F=�¾<8&�<�=7�s]l�ʪ�<�赼�K��X�<V7s�t�{��'����=�j�~k�9U�����y����:�{��Aƃ�V��8-=7�<�LU=˛]=���`���b/=���<U�=�;-����<u7I=Z<'=�<���<���<|Wn�T@=��;I�ܼ�JW<�I(=�@x=�B:>���-�l�j������}/�<�ZX�y�O�S�m�e�p<��p=�;4=��X��<G�����fL�[����#�<���<�%1����9=�@3�.���u������=�m���m�������p�*ѓ<��	�,��7C#�F��9֔�o���;��l=7_\<��;�q�<[y=Z�=��ż��ݺ"8��\=�=�/=u0˻J"��c�=�;.<��<��v=�^��j"�/t�;�"�;��伳%���y<Z��#d��+#��Y�=����H=i�}=����(:;u��<8��;l@��ǐ<�"�;���<�d�=N��<#k{�G�9=�a��<�Gi�,A=����;m�<��6<��<��E��Z�<=:�:��+=��=D�M���p�MK=	/=��y=8�׼]�<׻h:��F���`����U���G��r=ns/=���<m����<��<���;�=���;�ο���X=c�;G����<5�=����<��$��q�<��^�i�*�y+�;�Nl���w��[�0AV<�����=���4��U<=��b�W�=~d�<\@=b="��b�;���<��~�f<�ƻ��K<��]��'w;'�!=���G=Ub����<�H��Hã����;�; B<fS��=�.�Lnu=�I�<~6�4��<_@b�����=̶A��F��:9�;�˼�M����<��?=�r<
�R��>"�� *�l�%=-�-=��)�� ����IY��0s���<���9J�6=f����(��������H<��g< B���|G=���q��v��|=�0�<X�л&=5��U�=��=�w�<��q�Ꮹ���<���<foм'Ef<�Լ�����M��}�E=T���^���Ѽa<��<�n��Q�=A�������:�b
=��;�e<f.�<ߗ��1-<��)=Fʔ;�3&�W�B��op��
=㮕<_��<T���(Q8�����ʆ�<	tp�[;�;���C�F��<?N<R�x���<�����Q��3��i<7e�<��;���e��F=�=}����}ܼ�C���<�()=�5���N= ��<��<&�=yG�:�2><bGN=�-4=�����v��eX=:4�=���|cD�ˇ�=��V�Y����;����p���46=`�?���F=,=�r(���=�(=�3�7�}=ܼD��0�<����Q�������P�T4�9n=����#~<��=�Ɵ�7�Y�h�}=�M�;�{�<" e<��t=�E5<��=㷎�3�2<��Ӽs7<x�� �i�dP����	V(=�b=�����T=l[Z�O������R�<bώ���(<sZ��Y�;%�ټ�Z{=&[���k�<���;����Q����=o�R=��l<u����<�H�>*����2���R�O����:�Q<��v=��=EY9=��<UX=����7⻯��<����[P=pK[�3�<��=�{\�Z_;=q0$��G=W�
<���<$�F=7k�R��@��<\G7�����H���c=I=99:s�����<{�YK�<2F�Pkp<vK=%V=��[n�����z�<<%Ѽ�Ä<c�;���<�R���(=4 ��&��=�-]�#�O=�L�<� �����;v�4�ʲ0=�b�;+&��;���W�����]�U�Z<LԼ�-�V���5x�I�FR�@���E~����	2�9gt<+��<<6
===k�<�=�F�;� =~2�.8^=-4���궼�^߼-��[���hC��X�;C�i�61>��3~<�I<t?�<�*N��(<Cs;���U���2��P=�4b=�YC=!{��R�<�� �*�Ǽ ��<�IQ��mg��S;���k<4Њ<'�ȼ��W�op��	~<�>�����Ҭh=�|;n��C����<��<*�C�f"q��^��!�;t�3=thl=�.C�3<oy3=5AJ�����n�7�h=�+�<id伩����Ѽ�H��T+=����<�8o��Ӝ<Y@=�V뺋�.==��<U˼tJмOW&=�4O�ع;����<s��<���<A���t-����<r�O��f��X̻���;�61= � �R�-=F�=Au�;</��Z�J�B�#�j<��=�s+��]D=�͉�����=��2��<�r�<NL�;���m~�����w&�E�V�)]n=�ȼ<k�Q��]v�/l��� <��M;�D=�+:<_�$<W=*]=$
=������<�lF=��<Ѓ�=i��D����d�=�!�X�#�y�8<�����u��m+�����鞼5��;'J3��n���3� ؃<0��<��*� ��<��<��P�0�����#�J��'�:
)޼�@�<��<,�<a�[=I�<�	<�¿;���=� =�4H�L�N�~C�S�;K�^�%=[�8�d�����Q79�E�@�;�!缜�="�-=/ݚ<����&�E=�E=pd�������;�１�+=@=h=�-�K���LM�'h���Z�^��l{U��'=�d_�}�j�ձy�|Q�;�R�;PH�W�v<X�<n�9YVd=�Ul=|�ü6䏻��@��K$��.z:�#O=>� �u�=	�:=�����B�;@�5����:�%=�a=�L%��}-<��v�a1<sW�;U�v��_��]���3<��H=�K=���;l`���K=�q��2=���0�'=��r�V�==�����F<�7�)�:�<�=S�^����<��%�Ԓ�<ǻ�<o�W���>V)<�J�-_�=�S��Xb���<CJ�G����a<���f��n���S��J���#�򬼟b<���1����;�^+=�����۬2=r�q�s��<�f�;�c���i�<���9��t<H�=;Z.<���;z[<c<��<4�`�����oQ���D<�O�;Q�1�v��<����3�z;~�O�=�GǼ\���:/�/y�<S�O�ԉ<�=��D%;}eϺ*3 �W��;�z'=����O���}<�^�W��P(e;0�=���~]L��F��Y�I+�<�%L=�O��!�<8�������:=�GM�o�'=D��o4ͼ�4;���<�k���'�d�=�)K=�-�� #=F����Y=~�§4��D��I�h�ܥ�x���Z=-@��&~-=��gH�9�B=��^�)��;\~<�)�=#M<F"����)� ���b��/���c�;�yE=�fϼ>�@���U����k;� \�	h�y�0�+]V=�O,<HoǼPs���f�<%��<�� ��<E�q��5<`�*�)���� =O��;ƃ�=U#^��5�@Ś�6�<F�j���m�=���2=5*k���R�����nw��AS;f}=��<�(�<�ȓ��8���j;u�@YQ<-�:7褼1pE=��;mM�Xhi�'�K=��T�'Z=��AqB���<śu=��D<�1=� +�,E=R�<�-���I��`���b�.ZԼPc8=,=l�A=��]�ƺp=m��<�-����<�?�K��.�;�EW<���<�� =����l��<��_�6�="�@=�t�;�F	=�tO==�_=fͼ�/:�/=ѭ#��aj�!�A<EU� s=�����c<�=G��m=	t#=\��tbz����a�����	�h=X
��J���q=�3�q-"��M0��仸pv���<P� =�K�<��<(�ڼp55��:#��uP��/F=pW�K&=�U��J��<�#<����`i�%�o=�)�;p��<yS�;{��u�=��F<�
������j�)0,<�k=�R=ǜ�л0��5����;5��ꍫ<TI�;�_b=��Q�0=�߁�i� �逽d���|=KR�;ڻ2�9�S=?�+=�	P=5^�<଼S�	��Y�H<�<�I?<��(�w�$=ޓF=8U<�6)=>*��d�Y<�yU�� a=�.����<}s�<M:�;�b<˗[�. �<
�u;{aM��}r��8a<�Y=��^=e��<�!<�kL��79<uf�"��<��C���)=X�G��;<D�6�:;�<�g�)���];�=�@�<�輰ߒ;IV¼��%�;�+=�,��Q��<����C����U=�<���4���4<�u=IK̼�;U<@�f����yF;s5<��<��H=�*�<J�H=�QS��i<<�=�=�*�'���g�"'���;;�]�<݈�<!������λS�=FBo�aJ�<����T$���S�R=�����=��=��=k����C��B�B�f���u<KL=��<a���<��g=�I@=xh� �<��.Q=4�0=�DJ��h=��;�??����L����<��	=�[=H��<�.9�==�X��q�o��<*`�<��F=P�=���D=x]ϼ�6�['�<�%��4?=����ʻ�=J'����;��V=��X�>}=+m�b�0=}(�<��0=y#=93G=�ռ������<��:���<�Ty=�M<�[=������C���<�k�2K�<�`=$�}=�ج;4��<YD�<�����<���<YI<O.���U=$|�<- V=#DY�>���sN?<cOm=��.�u1G=7�@<��V���(=�����?��}<͆;���<�pU�����%=�<���g�������e!=�])��Yp=�v�=L#*<Kfռ%�<�6����X��o��7Fg�3�*�З)�S��;�]�<"(���[�(L��Ay��<%Kd��O�<sMd=�!R�����+=�c?=i�D<&�x���)=��/����G=<�;���#=)�<���=R�=5����i#=�2*=D�=��:ڼ�z;tM��ۼ��ü�8/=0�%���)=�jʼ��\���y;��=�PT<FA=yQ4��!�3��;�>����E��<l�D<,=��"���&=��ջ�s�l�Z=�+�<;G1��[�g<�q2��l׼֟/�P/R����WiG<}� �Q7��O1=��><�%];#�!�O�M���J�ں��|�,�:D��G=�p\=�~���x��6���[A��K����/={��<w0��t�<���<�B��3=缘Y�;=�=�vU�a���8y=���A���~�)�L��>��1���'S=�9���_���ʻ�8��*��3�J;�l���.U= �2�<[k���g=�0Y=,v�<��׺���<�	���d�9*<;u��<�J=~�=���3&��2�e=""=g�a=n/�;+�<�흺W��gЕ;v��<q]���1ӻD�M��_�;TGn=��#<ٓ���4���<h(=�n��)�=��c=S���hk<�|�������B��J�=�*l��D�;�6[=u
�����<��<�$ü���<�٬��@ټ�%=`y`=�T;��`���4=۷�<��S������EE�h{¼���<�����<t�<r�<�
�<7�s=B<$�����e����}��j���6�7�s�6�]=U�\�B��^�<k=;����1�$_;��=#�==�r,=%2]�6-V<�!<��Q��N=;�<��<�´�d�d�4ƙ�hB��AN7=��ݻ �w=&3ּ�Ԙ<{A꼗'���P;T����l1�T�ּ�24=B��0v���H���T<�1����<nJ���=��(=�K=���'4ʻR�y�~�E=ڠ,=�Ʀ��!0�2D=�k=$�=�w���K��kҼ�>4=	vE�-�;=�)�l�X���=��<�<�UT���<��(�7�y�Ļ��B=�}����=dL�����<s߼ZSi:i�Q�&1/���G=�<��8�U�<.�g�۸�<<|v1=g�<=�SL�+�
�/Tf=���~�z=�k	=_( ������<Y������<�<иm�ʒ0�Q�n=�����Qw��o=��"�]�<�����<4�/�b�:GwƼy0<�;=ȹ����x�=|P���<��<�ַ#����(��C9������W��A���\=<�/��T]=Q���ҼJ��y�@=�;G=��M�­�����<�_�=��(�;�=�=�?�<;�S=�2�<��˼����9sx=�������<&�<U8�ȑ=�)=Y�_;�2��6"E<�1�;��_=e�L��6=7�,=d�
���D�/�!=m =6�V�Gv@��2��꿼�8�)zռ�s弑5l<{n$��GQ��=�}=^��˝�<�=^=���;�~Q����<��r���;��Q��msS<@X<���<̵�<�� =��{��灼0N�����<�'g:� �<��M=N���&����Gl���q=I	Ѽ��z�tt:=Tl���T�1�<ʿY=�Ђ��.=�󒻫?�<�`�<�Q�<�&m=`۪<�΃�,����;Be�E�0=���<r�H����<yL=�M�5y=�ڠ��u�<m�=����Ǜ<��K��(�<��5<�d�<^ѱ;N�<����ǔg=���ΚI=��<��A=��m�߻]؉<T�#<*ݼU
5��*"�\=�2��|=g�<�f�<�ۖ�R+B<��q�����'�<S��</�Ӂk�:;F=f�u<`�;0(;����wv�<�3��q�<�P�< �e<�d�:oO�;yH=��<��=O҂<�;�<�80<<6J�+~P<(�l{������C�;����r=�O���<�^=�M<���<ϳ=�����g�<��<w�)�P 6���=Ҵ�<�TE=�G�<��<���<�s��H
<�,�<�
<Ȓi=��=�Wn�=��=�H����z:�4{���5���/�*�g�z~z��E�;���<S���},��2�L=�Ƽ�<�M�=�$�<!Ҽ{�`�b�[=��X��� �==�=nȔ<R<IQ̼0�����<L=8�H=W9��J�H5��ͱ�<&���t4=7��9�xX��<�«=��/='9�<Y����h<a��<P��T��<�B�<�&M�b����b�:x~�xsd�����߼� g=$U'��R����><
�����~9=�Y�:�K��t�Ȣ�<xv���{����*=p��=�O���ō<�R=��Z<�'�i��G~�<�=�� =Y]7�����4�M��3<EM#��\=3��<.\?=B�������#�<m���d=P��'&�B��<��`=D7N<j��<$����<�4��Xc��0&=b�=�X=H�a<:9���=*,(��G�:��Ǻ�FC=}S_=X
輰*6<y^ʺG�ɼ�H9<!�<(>=�|6�T�=��+�w��<���=���<��P=r����e=�H!��u�~��=t�<H�/���;��'c=�c �	5=�ː;"j:�۠�9�<
,�;i�V=TJ��*ü�Y��]����=_*�;|dR�r*�"�üq�=h�J��"E=��=<��\�œ&=?��<񌛼�·�&���T��8Є= F=HD�Ծ<79�<6��<�Y��ӵ�<	�I=� R=��%�ͨ�<4�5��IL=ၽ��=Ǧ񼩩0=[���=���t_=�"U��Ia�c1=,�>���<]�h;Ȉ�<a^�!�L�=.&*�B�J=JYx�x\U=������/=�6�N�<2��|f�8O���2��0��=�:ߌ�)_=� ����<��;E6!�hx�<3�L<cg�<Mb=9	<��=�L�<��^��5F&�ZN;g��<)�=��ɼ��5=ض�諮���)<�<c�K�G�(��� <�ͦ<<[Z=����&��/�<CU�<yO����<���<�!�<��/=�d$=+H<��j;���;,"<�ݩ���mq�<g�j= O=��W=�vg�c���mx�)���v=�4�n λ�#G�:sF=���=}㔼���>z�������|u=��˼��5=|��:.:"=�<�\�1�=K�Y���=�ώ���	�7'ż�8�0���J�[��������f1�#PL������S��U'�A��<XZ�U�~�G?Q=�P�_��D��"G=T�<��N=��ϻɲ,�eE&��Yn�x?��B� ���_9�<u<�����!�?�0)<�
6���*x���1=���<#�:=���<�췼�ͳ�+GC=��;=<9*��Q<�rE����S!�;��+=7�=@�@��=�-�%�b2=�>=or=�[=^�=:��;��?=N�<ς�<�c�<3?=d�<HHW=��0<]��h�:�v==м�<�W�,�<X\<�:��i���]���5�_Us<T~ʻ/��D�;!�����<�'b���B<F`��F����X�<l̂:RI�C�-=O�<�?Z=�:�R�S��8;�9%�M�^=ጃ���Ӽޥ=�=3E���<g���rOr��Һ�R=E|��U+�Ӵw�˒�<� 1<S�l=�2W=�]_���<�)M�Qּ�k���'2�Dh�;Hg�����2�l=�ԝ<ʐ���U�G0=��U��_�<�P���o���;ʣd<�$����:.mE=��a=��<A$<%YR=�_̼s> ��Ǽ.A=����ߴ�0�-�ᡢ<<�/<�{#=�u�<��a=�s*=wx:<�f4=�4�<SC�<��=�c=�i=k���;���<���<��x�/[��̾g=� j�� ���='^�<���<PCV�D�R�:���{���=������;���<�N= �Q����;��V�d�<J�<M����i�=��eG��O=����S,<�E=����$�<�ߡ=[�Q=��=�Id=t�w<�m�;���<KUB=�"g��6���9Ӑ�<6�=v=e�K�aĞ�$�=.���U����<���<�<S$1=-���;�κ��;u��<6$���=ɵ�<BH=}M�zX���꠼������!�	��0��<���Iغ���:􊽺{1=�w�<52	;�1���F=��9H2��Յ���9=X#��CC���o=����1q�,m�"XP=���<3l���_�ū]<#.t=��|����>�;�%x=��<��0=�|c��v����>��e��/<�����,<�YO<�4�u+�;p��<Ђ�<d'A=�<�<��.�Z��a���
T=�y�D�=ؿ���`��}2<x���=}�)=)HR�����+���V`��K={�0=U����r+=�Ȅ�2����<����Z؆<H^=��H=���<hC=3@����<�~��n��;��<%=;��_��qE=~ǿ<�RH=�=���<M'���[q��!����E��zM����<Y$��,�<t��t��;�&���u���9��^��.T���)<�[�<��I���!�զ(���S瓼u���O%�<(Pr��+�;�?üv!��t��<C�껙�J���<�B��*#�n�<ڔ�<3w@�#�<�}���`=��:=�S�<vi�;ګ<[j!�Q�;nf��1�`�=&�ϼ�`<f��<yi�)�μ"���<%la=Vj��[+=��<�4�������;<M�;'�����;<�=⫯�B�Jc�^?=P���(=U.=� Q=~#���0��1=��=V���E4^=��<�E��#� �9�r�?����J�=�x5�����i@�x���J=�l|<�K�<Ty����;�Q�:Y3�0����:���;��!�$*��{�#�������&<�U�;- �;e ]�}�k=i�'���<�(r�%�v=�X�=B��^Ҩ;D��<�{$=����B�P����<����Q�K�L�=�64=�K����<��d�W�����!�lm�$~����"���M��[O=�n���0�a�)� 2=�B�:�f���&=����D�'
=�ȹX�F�����P=�0�����vǀ<K1���*�����rȼ$μ����bm�<��l=^(麞��<x�ʼּwv<r`�=��[���w�f�K��d�28B�üռ��=F��1'=rߜ<#�B��{��%֥<�}<�D��-�=��ϼ��z�� �<�^ ������-<Zb��U9�ND�<7=$X)���&�I0]=U�{��c=21=
E*�"�Ƽh c��X�i�t��(�����BU��q=(.�<2P�<T��<N.8��NU��� �6f��&K;h�ϼ�R�<����pS,<�@��k1��A=�*�<+�1�AY;����7ϼ�삽�פ<k�t=pq[��� ��t�<�9�=�><S!�<^V�<o.=�^P���E�?���Œ�:R�Sb�;]�"�gW��w���<=��<��s=>=w�Q=����p�<x��=�40<���<��z�������;"oz<P�R=�nJ�7w,<H��t)X=�/P=Bq@=	Q������M<O�,=B��;,O漪���v���,H<ڊ=�⽼\�<$(�:��<�A�<���<P��~�B�{���Y0�<D鏽�=���=j�=�aE�[^=D!=���<�LH���;|�=��=��<%�.�UQ��iq�Y|<�p�6�=�=������8=�=�<��=�]��Z�X=����< �M=&����E�_�Ǽ��z=���֭/<&�*=��;w�`�'��uc0�����!+��6:=���<�ǡ=�f=!�������9=�0:�x2� �<�F��m�=i��c��!�=z��<�V��"�;��u�1=�ʼ��<��A�觩;�%=
C=�*P=�E<?=ks�H`#=�Iq=��T=�i�<0��z���%=��X=�=8L��[K8=�<�SA=���偈;�B='�-*=M0�<��=�3P��=b=j	<��/�.�<�=[��<[��>B<&���w%]���W��Z=9Z	�~T�c��^J�6(���=m��<�G�����	3<�$B��^9=��4�`@C�?���6��R7<��ȼ\-=o�d=��ܼsg"=��=�;"RY��6ռ��[<Vu��Y~<*7��b��;"�;eC�;o`���ᴼ��<4���ݽ��y��<K5��� ���= ��L�N��n�<�h�]ߺ�̎���׼�u6��B�;NLB�-I=��h�uL�;�r#=g�ż��=WD���=1�;q^T��8=k+�:Q{<�R�W@�;��M;ijٻ��r��B����D��l�h�k<	�85�=�ƫ<�36=��4<��Ҽ�X$��;'�>����y�;.������������w��)�<�=�O"=be���4Z=���=R��p���v�<�e�<T2=�7x=���<��t�{=��=)3�<C�R;���:�إ:�Ӽ`G&�w�*=R���|5��d:�VA2����(�Yr�<�I�<�ZF�
&S������<�}X������t��֛���[=Yf<��:=1or=��F�>s
=�g	��e�;P��<��3;�����$=Z�B=g:�ZFS=�k��3<��4<��j<��=�fZ=�$=�ۤ<1F���&{�a.Z�+���KWR�(�c=|��;������<�W�'�,��>%=*P=�P�;h�=���<��W='@_;��=��;�f�<�5�;��)�������	�V�K=�Q�'�ȼ_��<J4�3�S����=)nS=m�<S�G<K�ּ��;�&�><=���g%!<��Q=	P=u�~=YG�<�F��@�<O$ ��ռ9�=?��a�|��~[�p��<h5y�~"D�y��Z�<JU�DҪ�BP=���\�4�ܻA�$v���d=ڶ=C�¼�3=j��,4�*a{��|�(�;���M=?}X< � ��=��o-=>ܮ<���<��U=��м�2�=�����<k��g8k�VP^=J��������9<t���:M��a�<?�lU&=��=n��<�T<��<�b�<��<��a���G� �%�=߁�<]�<S�I��C!=8�=���������<@g<��м��8��VD<�F��y�<Fd5��D��O!=W�
<T����V��+�X�S��;{P�<A�ݼ���_�i�|̻'��O�X'��͞<-�8���;�6�x�=�5�໸��d=�"ڼƬ+=��м��Z<N���5<E��;
k;\[=�2�"7�P�<S>�4���58<;�Km<�v=>�W�ռ�\&��!�I3i��V�;�u�<D��<z%7��;
���;��d<��⼠�R�a�+=�˼~�1����s�q���=���<�/�	��.�R=��=�� �<�)=`_�aJ;���6=��="�N����<�����<7�:���<��K;!��fM�<ῢ�o�=gd�=��<�V�<.t<��>�;�*c(��!;[Ac=�(��Z��)�n�%a=>�"=��=no=��2=�u<[H=�lƺ�9�=�3<��;�HL=[�˼�'�<�;��7��	=��<��;)�L�j�^=Vr`;��}��v=�*��)=EU	�R��r��</<% =��a=���<ӵ�<���6s|=D�+�G~�<��;����T�����W< %�o뉼ۻ� ������lӻ����)��мz
C=��<�72=V�G<��=^�J�
8��q	<��l=�Gk<?��;���<.�<��ټC�<;�*=�8���7=\/= S�׵���z��Y��;�Y�S���i<� ��,=E�>=�$<�a2=!��:/��9���<j��<a��v��*=8%λ�o=� j=qZx<p>!�F�f<E�9<�IM���Ǽ*OU��(�<��9=�z�FiB=����V�=�7�=�J=E������[�PM�����<�û�Fi:8�>=�07=�'�ZR��-=t����K��}�<Ps�;�Lh<i[P;ίP�	"=��;"��;8�;y������I�O�ۿ�<>&�<o�\�~��Ɋ|<q(��~1�<*�=�?�<Ԃ��A��ܱI��@=>q�i&d��+��H(�;���^S��Qƻ��U�9{<��}�C���kW�8�;��<�j0=&��<٫�<w	�<�C�<WH#=�V ��~�<��=y{�L�	��..=�|2�~q=����_�&��	�=��<���� �3��j��V���A��<m`�<��M������X=�Q�=��a=��X�i����8��K��а���%=�4��Kf�=���<j�=^K�<'��<��<�����	<^����ؼ件:�<��%�'b�C���V=��<���<'��� ��i=��Q�ƣ:i�y:��<��6<~��L*<�(���6��%���{<!�d=BI˼�(5=�9=-��XX=BC��+��<&�K<��ʼ2���ʃ���c����<|'ټ���~��c�<�e*+�j�<=ȡ��9x��@���/�
@�c�<���=<X���R�0�O85�,=��E�H�u=o���}�;���<�A��Ɇ=��<Y�k=�{�<���<Sv`��4U�1%<�8}<A��;�/;D�?�/������n�c|j�#�=l^�gx=�%����Eq<7eT;B!=O@b=�	��b<S�<�<e X�v�M<nH���=�`<E�T<�pj�����o=���҃Y��h��䒼t�!�f^��c=�Hϼ�[=�E���o�<$M=�b��
)�N[=�=���<�~3=��+���;_mp�aH=�q,��-=!�<y�4�i(�<7����<�cR���<�Y=�Cݼn�=<�<,�><��=�i.���q=}�<'�;$wļ��K=B6C=�'<4��<p�G���8=➹�r���M�"=�g��vp2�0�6�<�=�>� �]<Rl��)���=mp���
=�R=b�(=�Ǽ�"���
;f&�=o z=mz=Ww�;�T�:�iN=���".E={�;��><K�<�����6��L��*=�	!;}�j���<"OD=�j���<u<���r�<��<���<i=�,�G-;=�x)��8=--��h��σ�<�uL<��ڻ���<�a��^�]=�=�TQ��Nȼ�g�< �<+wE��Y�V�k=/ҁ���8�a,h=,���Pp��"==Cļ��g;0� =�d�<�P��\�;�C.�uK^������*�s��<J�	��94�v[;=�z6����:>��M����&���yS=6*R�f/輯%��F�<Zʻ�t��,,<z�4=l���α;��0=4_b:�<8�h�YN�<��:=��T=b����(���{�;�,(<z�;����ѭ��&���=&�,��C=IC=~=:����	<6m�Wm�<FJ���R=�#=��<�&g���I�T�0��Y9���~<���V��S�v=�ℼ��%M�?ԫ<)����<��=0�߻ў�<,�e=�ڻ�Y=��Z=/2:��)��%3�<ǝ�Lpj�b�)=A7=�����;��ػ���Or"=0~�;��R�q�<�j0=C!��oI��+���<ؕ�<	<���o2G=тf��G�<���� <pBX��+=�M��q9=#˼a�f���==���<�h�<É ���
=�=n|�B��<B/�<P�Ǽ�T<�T*<�'t=D�|�|"=�=��<�n����':Ĉ�<��<8EƼ��m�=陦�X�2=NL|�͑s<��f�eCC��oF<�ة�_	�;�Ύ<%�I=I�I�ٽM�5=/��� =�3A=# =�;:y%�;l]</-���=���a�S��0�<	 �<��;�;3�����<��=� ���<�M��{`=�N9�X�<=Z �x,�<O!g�8�`�nV�<�
���Nڼ�L7=��ʼ�;~��<�f=I�%���8�W=��=�J|����<[k�s9d��{=J^ӼM>�<o�B����<W�<�y�;B��5xl<!��X�=�=m"%=G��M(=�0= ���@�� ���=�]=`��ςӻ�m"�����"��֜<e���Ȇ�?k���S��Z5=�Q��t]Y�E�G={��<�H6=��X=߫;� ��������<�+���M <�#*���=�uQ=*t���������:��R=��<�=;gm<�q�<b�f<��?���0��A��_o�eμ�pѼ�d��R�>����<���<�*����;�v���Ƽς��)� ڦ<v{<��$�� μ�y׼��=q^�, 9�i�=o? ��*��*�<z�'�����:u=�j�<m���a<�X=)�Ni�<`�<�}k<{���S�=��m��m=�฼��;��/�n��<M?�<ܯe=a�=��w/8�r�{�o$%=3fj=h�<R�6�V�<����	=�<==�D��<hO=��_���s7�\�;�h�:EmҼ=��<�^ۼ&�A�M?H=���;u=ʥ����1�0&5=A�=X�T�@�<=G�<\��q �tV�as;�!'A=g�/=k�)����<�#2=�Ҽn�!�{����:=�F��i���`��1�>�[TR�5��<�H;=�߁�4�\=��w���A=�M� �=O���4�N��(M�]m=� P<�uz��ҙ;�J�<�w=�L��"1���c��j/=J��sh���l
=x�b<�.;]��0=��O<��P��Y��}<�m��A���j�༔��<WN�<3 ��t�<l߁=z<�"=���<߉��}jm�A�t�m��;�{��we-�w���f��E�s�=��/�q�4<���<6��7��-b=D-�<=E =Z�:�'Z��;<�m��LM<=A=q�<)���l �qN<��=��=/�j��]y���9�c4A�7.=	=�	�L����:�/�a�/�ܣ/=�tI�0������R��51=�#=%̩:�=
��+*=-M�;⺔���b<�����%2�<t���8*=st0����V7i��웻�#��#A�~��!!��<0=�u�<�-份�!=wK=�|�<�Q<�TC=�5=��&���1�� �c<:< �<��c=ЩP=�`�|_�$C?=��"=��<o��<�4O��,T<�@��7=i��������Ͻ��&ч<m���</zS��N�����;�at��Ѐ<Z�;��1=8��
��<=%�;7�<W.�٧:�'��h���L
=����S�<�4i=$� =~�3�-X���.��Z��(<a?T=M֬<�5=l&�<l�W;�<";9��<�΄:����Ӽ��7=�Qm����<Q1`����<Jޤ<G=<��E= ��'=�b�<�&����<^��T�d<
����dN=,�=��1=����J�;ΏӺ��=�m�;m(�<��C<=�<��g��R���-��`�<�*F���&<�� �1��<V�μ��N�_�<�+
=n�
����<;�w<�q�<<���m�G=�|���ټ�U�̄�,�P=DH=OK
���=�*j=�"�ȶ\=�c8<�<�j��<�1=�-@=������<?�<������<�'��rR���K�4w�;\�<��_;��V<�G��2o= ,�;�9Q<��0<5�����Ἔ1��� <��3��˼�&=�բ� <ȧf���
=�|��z�<�c�i=�:�`#I���<�g<����4�T4^=��#�h���+d�<R��;mD�<���;�4���x�q�-���v�W]�-	�FV�<{�G==�v���b��X6� x���;���,<�a6=�y������<��+=F�=�i�<>�ļ�r�Y�O=��}�K��<2R[=�!�XM=��<�p�U�;�1=&�ּ�\L:9l=P�Q<㽻�I=�V���D���r5�Փ�<��E�<�4n��	��*���Q��o<=I�g�&. �!A�[�Z��A�<`<���#<W(Q=�Ԯ��,9��c�<ʆK<W/���v���<p:1�y|:���=�(=�c��u�V��G�.�=�༖�=�⵼���T�k<
��<V�C�d� =�ۺ<�9��LH���e��e0=kǩ<�c���K�wJP�S����:�<��R���D=��K<�o7=�J�;pg����
=` �<*����A=,�!="2;Gz='�Q=("-<Z�!��F=dͼn�L��Pb�<	b���ۼI����6��2�m�
�N�+<�D����<ʠR����ѝ=��a= ^��Mq�D��������J��Ȭ�R6J<:ӻ���<>$�͟ü�A���}S�4��L<1�<��	���<��;o�=Tg�䢇=����<ql���i��������2���)��e^=}y/=�.�<=��<Y�����V=�<� �� �;~��<F�<z%��KvH=-.k;��<��c=J�I=��f������}*�͘�B�d��􆱻}U���,\=������V��M�K<�<^Zq=����Nz�;"D�<%��<���c�O<�9˼�����ǼLv5���<��<�<�=qF=��|�cr#=��N<�O�<�̻��ż�[༆�ƻ��<]��;��3;%6<�{�<�H!<�m<��I��(=G����WS����<Վn�~��;픰�L�)=|��1�!=�j,�����
��<)]M�⍼j�S<�+�ض=���)����<��z��Y��aM��6��e�;����e�C<�`�<��=2��:E=	�P=%�c�4s&=fc�+�g<�5����$����U:����<��]���=�M�)��<��0=f+�<.���ךּ<�b=^�����+=&1=&_"=�f=�
=��d=�^=96S���#��A�8�^=�^0�te�ؽ1=��<S <kk�D���ݼ�Hm=3����?��ϫ<]a=�ʼ$D��:���4�<t٢�>y=��<�0�<�fR<=YZ�������&<^7+=$h=�!,�lA���T��`n��xE��wR=�G=[��P�B�ڬ�<H�t��=X��<Ҍc���v���_;qd�JǙ���<��� �/X=�&�<�a<!'�Z���_b���A=Fv=b����<�.��n3������g=��ּ۔<Jɢ<<z�l��;�����<P`�=w˧���=��"=��|<ŀL�p��<q7�_r�<��=�[����;=�ރ���=	=��@=l��<(�߼�^ �7/<MϬ��E:�����Z���@<�]H��=&��<�=)�_=p���ʈU=��/=�:J=�b�<2٭��5o=�lP�=��;VZ <��w�sA@<d1�_ !=WlQ�cF��>:��Ǽ:��<�Ӽ��<3NE���'���U��i�<���;��+=zi=��<�H=�e��J��� �<���<�"��iL=��b;vr=���<�=]�c<�=T:�<�=�+�֎<� �D��9��;$�ռg`x;Lb�3����<��`=�	���%=Ze=@Q���S���N<���<���5x%=�t��'<���<=�o=��Z<�/e�z�><>�@�^'��AU�a`=�ƍ<�h:= q?=����°<�:$��l�Έ���/?�t�2=+3�< �@<W2Z��~�<"i2�� �<)|���?<SG<���<|]�<��Y=�*S���E���8<����n�;�����p`�f��<I�=���<fW(=�~N�������*=���^;�����+�;C�d<�2=cW=��t%�g�"=��!��$�\ !=P輄ު��|:����b �<��2��b�<d惽�E#��hʼ)�(=����2�?�L�]��fP=�� �O�/=��_;I�b��U <��-;�%����<.�=cA�e�X=�`y�HZ=�[C�f���2=�=�7��:=f��<��<���<��8=1O";�>����<IX=�T,<��=����B��@�%SA=C�4���!=#QC���h=��=��F���m���l�;�)<�=Hr��5=��H�V�� {=�,���P=jH=hy�<*P=Z����Q�<< ͢<T��<v��<�7�ݐQ��B�:!9	=����.����@= �h�A��:�*�>&Ⱥ�"�<�=��<|�w���;��9�8e����;Z=@J!�'((<|=p�м�#�<�!��dԼ�&=��<� �0=p<�l�~=^j��r���g<��.=�,=��=ϖy<0C��7�}=̙��^�n<1b_��.<q�=�M�1V�e:���B=�A��&��<?��<��!�g��;�H=��x��o������W=���<Z���iP;=�=��7�dVq�|Η<�Ȣ<�a[=��(=¹�<{ <[�<yJ�;�h�<������vmG�Y ��5��<�<śû��<c�������=�;`�?���m�����@Y�=p�T�ks����6��7=2�\=�|h<�@������'���;v9-=8��<f�=w�t<�j=5
�S�6�-�=��?=�K�1UN=��8������=7e?<p�<���;�CF�i�<5���ٲ	=:���A��()p=��h=7=U=$�<=�6=�==�x���rO=��߅<M���2<?P;�F,=��<"0��2��י<+�%���b�7=��<=�����L��B\�A��=�ҫ<��:u��*=?�ü�8�2+;�o�%= �߼���<�#�<J��<4 /�%�e����"�<qm��/<��A�x�)�oѼVw��� �<3G�����	<�#5���y�Kő=0�һn/�k`=�by�3��-Q>���=x��<7ڿ��xl=5��<�<r���������<�i�k���d\=�����>�B���#��`,=�=k�v<{Z�<z�ݼ�+<=�� =-�R�)�(=H�E<��E��������1<�.=,�0��6�;��=%���ڐ;�_Y=�]\<�zA=�^��KI�a�=���<<֬�%�7=:k=X?<���<�==���tC���S=�9=ߤ�;��<�,�RF�u����i.=+��Q�˼{��9�����r<�@�<������<���%
�;�v�:x��n���g=K]1��dE<@�]�5-�L��j�<Ӣ]�8��<��=�%E�L�¸���������<pK�^�ԻF�C<Сg=��=�Q�˾a=�6��Q�=��<}1�I7�z_üҶ=Ǥ=3�)=�.6�j0�������.�ﴒ�o�;=�8=���;�FYl=uTn�A�t=�<�-=�T=��;*�0='?=��<:׷<*	���; ��@����5=y^#=�g}<�"���^�,K<�qҼ��*=���<�a=m�=U��<S�1;�h=����|5�3T���=@��c��96��ؕ�<���=6�<F{\��Q=�!\=6�Z��d4=��k����<��<I�o[�XV0�T+(���i=��k=��=T����t�֙<���<��N=��a=�<T�=ƪ���X=�9r�L���=�D��Ƽ��!<ÿ%�4Q=aX���p�);=��<_g�;#����ӵ�<<je=IP�<��=�=�U:;֣��S�������o=��+�c�t�b�$=�%f=�-�#K=GLT=�14�X#ѻf������?��;?��Q�i<ys��
� y&=��=Ȱ�:"����h�/8������M=������[�I�X�����<Mt;�8�=��T=�/��)7=,���=�F	<��_=2��K=[I<=�=!4�{�?="�<��W�d<&�u�R\~=߇R�&��1L�<j=�U;�x�<�,߼F��<E����-k��42=�4�3�=�G<�H=4$��[7�;w�<9aܼ��=�^�;
�x<c9B=_�?�p3�<?Y����F���*=S����ܼ!<�<���;f�L=�C=Z1�;��==�i=�.������x8��a=�۾<��)=ķf��d�<N<��=�7]�����Fj�!2=������?<��<��=L���Y8�h�<Ʒ�<M��pD=\��<?MH=��4<�v�;1����"=����|�<�MF=�QƼ����=β�<"�j=��=U^�,�ͼ&�,=ғP��B-�R��u�;&(���&=��!=�f.=�� �v�i�sr==b6O=��:�â<��<*M=��:�����<r��}�=��>�8�<>eͻ.X�LY��(E���%�tb�W��;��9���(�#c�r5=ow[<~���\<=��P���<��K=���;(��<x�d=(lB=q�<?�=Q�#����;N�!=�/�b�:�e?�ۺ�<�"@=�߹�m�<�W�ޛ�9$�<�q(=�f��Aa������4{�$/�<yl�<	�z�<n�
=5��٪�<96y=��)=0��<-O�<�=߼�<Xc���W��M�<s6���	����)��8�c��<�]�<���<�M���I����=��1ڼYM"�4��<ĉ�8������<j�=�'��)[�sO���+�(6O��&�<j�=���< �{�<L{�<�F=8��<�$=|f+�A�/�"��'�=��b=��<[�[=��I=�ɻ�_<�ڼ|[�?;��<�	[<ȟf<(�?<Մ@=���<�Ad=<=�<;<?ϻRa;��P�UJC���*=����
|=e�s<��.=K�8�����ӻm��<���<s����H9���=���<�|=�}c��'�=�en�y�$<��~�$�'=Msֻ�W��!tƼah���%=7a<�=XH=�0��0��X!�<3
^��=9���:�My<�$r��E���[��A�(=�"=��̼A�Ļ\%=��4=6��<k1@�6�W�6��W<�o��	N�>	�<�������<�,M=_�Y���x=�˼L]��.u��=Pἱ�7=�A��^�<��=�&=)Z6<����F<�ƽ<1̼<�x���=GѠ�s�0=F/��s�א<�O=�Mi��B2�|@��Uu-�"�#=�,<�(�FfǼ�,<�?A���4<�L��?ȼ�ti=ب��j=�	N�%	���_=)<�<1��<�3F=�%=�=m��QF���=�s@�(|�����e=�@�<䃼�V�<��"���^�F��p�n�@���?t��� 2[�ko=H�%<�=��zm�;�t�<�7]=-pp���;IR`�L�X<Y7��y�<n���<(�Ѱ0���)=^Ǽ��N=n�0�	G=�<p�=�5=��̼�B�<A!P�Q2�����R>�[9(=�I��C�Ȳ=�C>1=������<�=����8f�� �=�<�==��������<�^�_�/<h�|=�_�l
��%I=<N2�r4�<�G�S3H=�a���3��Ο���j�)�%�ռ�識l:���0�e&�<k ;<��Q"o�����0=p9"=��<Cv3=VQG<�b�3\�͙�����B~<����=�c=��5�c87=(��<Ź�<xD=��D=l���1��Z�*�Z����<f�<%��;6cl<�TN�^=�*�:_qZ�V��<U^�<m��<�[�^/=�N�<C����eS<;<=�v<?-"�������:�ܸ�b��<$A�<f؜<x/�<!�9v5[�ͩʼ[T=�&�T����,�E[09�����C=w��|���T���4�x<�(=3=s%��ٺ\��
a�y��d���tV�<L��==�O"�Ӣ̻�"H<&�t=J��/�=����,�99�<���<s�<�	<[�;�GN=�����g=sS�&V<��	��d�=�õ<�K_=�%�<#��`��d>=W�=��	� �<8�u<ꍁ<珞��U�;*�%�<�!.=�S,�R���~�G�ټ!�o�f�d=7
�:C�Ӽay4�{;���� =y�<9�=�xE='�	=�=���<��b��o�;��뼃�ʼ*u=2�;=�>E=�Լ1Hk��}Z���^��T!93���?A=�=�F8���:�f�<͡K�n��<���<�x;�n={��<�e=ia�;�<jCL=㴻<́=Mo<

S�gҸ���c=��<mk�o	�`�d= �]��
=�Z�<?��s\�<�ڼ�� =E>˼Q�u=�u=��<;6�򼢘�<
�<�˼;��I;�=%=���~��<BaP�P�5=Q��<���6�C=S)=��/��AO=��<����&�%=�ǝ�<
�<��)�ɋ�b�t�Ŀ�y�<hƼ�k=�-����D�GD;��<�����n ;4�l=��/� <!�Լ �==�5=!A�;X�<#B=�*i��-ټ�6���N=%���Q=� 6=������3=�=ʰ�<N���td�8;=Iۼ�L=\r�n�;�(V���<œ=Y	=��R=ƛK�Gh8�1�%�=N3C�J	���V�rÜ�̇|���=v$�<6=g=o��zv�<�)p=��e$��8=w��L�/=�5�<��E��� �%"伽��BԼ���C7=Sh1�i��<>�<�E�7O;<�)�;
+K�d�g��Oe<U07�4�#�N�%:�K�<,��
K�<j@= =��=�ݖ<˓c��ͻU���ņ�cO�;�O=	����='�:�<����X=]��:�X`��/�k�=E���zï<ȅ�<�$=2�@�ҥC=�A�<g�¼�����<�A�<h	D�����Q=�:�7��<ʎx�[D��\�����;6�G�u�>;�E��a_<��м�����i5�g>=Rg-=k/����>�܊9��IY���ռS>�H�H���<�C�<���<��/=L�`�AU*=��A=�{�<B���O=w=��<�`&��P=+�ټA�m=�S�����ʓ(�9�=�H�<)ݖ<��<�}��Ը<O�ѻ�����<��U�@����?=~�(�=+�<͇����U��H���`ȼ���`�-=b]�����sh<1��<��i=9�I<Ns�<aWV=�?T=�O�<
帻�3�=��.<Дʼ̃��4\4<.�;^�<��輶�n=��=��	��0={#�sO�:�d&=1�Ļ��<�ϫ<Ե�S �>����3=�����м�N��>����?��(����=�6�:����|�:TdM��
��Ḽ��t�<��J�'=xQh8��$=��J<��S��H��A����;G���x������v��	��<�r+� �!��������<�h=��<\&Z�)K��]ar������񼦶#��p=�<��'R=ؽ�<��<'6J<
�0�ټ��t=��&��̼�����f�Իmx��fֻ<&l=�i��z���g@��i�=���;�e=�5�<$�K��M�;I�=[�M�Y�����$<(�?<���i|�x<j�<��U=��8���s=��𼾯~����@2=-z/�0)@=��`��;�<�=��=E�<���<*=�v�w����Vżʐ"=�~�<�`�����!��_�=�x�;�=�)/��ļ�_+���;���%�E��'�<@*�����<K�zM=&K�B�`�#	���m)�;<c=�I�����<��ɼ�7��i�*�#�/峼�b#�1�������'�-���'ûѺ8����h＜�<�yK��^^�ge<����#�;�����<Z�<6��;�I����3= =d=�;�m<�<I��=�b缌)8�U����<����|m!��FY�C2Y<�=~�`o=��]�/D;���0!M��)��)K�<�7������3=��=df5=�&����=y�й{D6=���<w��<�k�<vq�<�R"<��м]�R��L��;y�<���,U�<Bb�<�R4����<82=�܏<�c�Z�0�<|F�os^���l�8R�<l�9=T��9�@��(���J�XtT=�ZF=T�=Y�<W�{<�V=�7�R�_=��M=������N�Iڵ�LT6�Z��<�0ܼ_<�>�=�}��"�xv߼�)\=��E<p�:���<OY�\Kػ���<�K<-�<	?=y#�=�0��ȼ|�=Rjn��"��uZ<<��N��<�[��#�}�)W�<\z��T=�.=����c�<��i<4��1=��.�L\-;�> =vg%<�	B<��<���V�:g�6=�;m�&L�<ѳ��B�׻�3���c�:9�K
�<��m����B��;ɪ�<ch@=?j=7�=z<V��(�����<��<S���>�u�q�d=TL:�;Al�N�N��yn=�Q)��&�=J['�6;=2A=��>=�~�:�/�<�Q[;�༵���7�C=W�=�/#=7W&=�=!=�7z�E��;m�s��U@=[��$<�0�J�b=���t��h�!=+C��v�<V�ܼﵬ�Պ����m�8��M���<u��e*=�X�/I�<�o=���;�[g;*P�����Lv����<n�>� �I=� +=^f#<�<��=�o=ĳb����������<���<��<3�����q�>���R=x $�,���kA=� 5���`����p�oe=U.=�~�<��/=�[�:�g�	��*� =&�P;�g9�-	��<�-b���,��e)=��T=0����=�E=�H�<{X���;�<fFj;�X ��@ ���^��G�<���<��t;��<��<Ѕ����<�_r=ۛ�%�@��xN�<��6�� U��o#=���=�/m<�޼Jc��g�h�V�j�tRo=>�����^�<��5=��#=�9<�8C�Ů�~�ټa+�;�^9=�Q�-Ɓ�q&e=ևB=���J=��F���=��㻾陼$>��=����<�����&I�7o�I,�����	�p<��-=�<�,\���=�dA�
��~�cN:=1�<��k��J��*)���<�%żl��<��d=���(:1=�;=|s�<�ɖ��>8��}(��aѼ"p=�a��A=U�;͛�<�E�<���;&=8��<��4=f5��4��<�i������F��$=��F=��}<��t:���=�.f�A�,= ���n�(��4v�f�<�_=���<��<t��<#H�=���:d�[����<�=A_��$4=^Z�`���t2=\��;�E�=��#���H�<���Ĝ����;˙����;S��<,���e���m6�8B!=	 ��r���ƞ<��<�wj���<���߰;=��I=;�_=�=-w@�!�׼�nj�W7'=��<x��<J�[��o�f@M=D�	<�P=w����YC����<�VŻ�3��Z!��&����=�r==��=���;j�O�{����Ɯ���:����l=Y��r{�!�<Z��<z�=l����<m2=ÿݻ�1�;�B���m;��<9�p�='.<�6�h0�=�<.>�����<=	����<�v�<D����»�ʦ�˚�<:�W�L�=��=|��`�\s*=7���B��:��/<y�;��ֻ�͊���8���S=�hX�%�;�T�<�X/;kc.=��ϼ�s*��>�<'(J=�*1��)�<Z�?�'�]��9�����<�<FUH=���;�3�٨<��Q�U��<cp���A�A�3=�M�<���p��G�<)q��dvǼ�1y=H����K���@<�r�h�o;��<�h=fZ=��L=D7�<���;�XJ���<��뫻�l����1�	ǋ���i��,O�R�L��|o�gk��tV=*[��ƻ�B�<p$[���a;�;��8=��t��h*=ꀅ=w+_=� o�3|�<^ ���G��������|U�<�x�s�9=ye==�H�P�=Nų�T��Q�<�-=[)=$�G=���x0=[a$�\�%=��<@�N����<� X���u���<־����U/Ƽ����G/��M_�� �l�@=+��q�H;��<�k�7�w<�e������ޱ<���;PE�3�ü h�
'V;l�����ݝB�T}]�+l�şo�5�F�p�c��]�lt]�I���S%>=u�[=�������1.=)�v=t*ؼ��=:?=�k�<���<� �<��Q�ׁL��e��X4= %�<�_0<�$)=g��<��J=�лH���߾��>w=l<@]%��R�,�c�<;s=;�=j��;��¼�E��k=��0==2@�;(��<��<ט��ѓ<x=li���c
a=�r(=�$R=ۓ�،V=D�4=���Z�e=��4��=qm�Ԅ����-���c���<	=ק���_�<]lP��=8�I����R�2�<�⻛s���/7=3�:+��<�>=��,=�<��~Zc<{¨�*�Ҽ8 =���<D�������U�<Z�<~�<��/=�<c=ɘ=>;A��'�P�+<J��1�Ѽn�"�\1�'�M<ZW����<u��;8<\3�<�|z<�����n��
�<��*�V�=NO=)w�`�*==�.:w*=��=�g�<h�=�aF�%�L="�<=([�<��;��(���W�\I���t=C���"/<D����"v���»�.j�^�Ҽ��ʼ�K1;��6<`.<��"�,�V<y�:��͈;^�%��E=. �~I�P%#=Ħ��;޻xIX=B�3=�{����<D'G=⧽<@���1����{m:u\H=�:��=tT����[;��=�'�wp��נ/��/=��b��P3=_��<�S5�$�Ӽ] ��*?=��V�6���t(��}j=��<��\=T�g�]��<��C=���:w��;���T�*=1N6=
T�<Z�<!Ij�*��(�,<_]=E����;���<�ӟ� ��;c�̼�K�;܇��.A�1����X����6?�����H�aw�;+��r4n���<dv��Y�;�y�=Uo�Kb��#H�<��߻	m���1��=�aR���U=�g�:ȁ=VI��OڼEe���Ǽ�7Z���=k0��R��<�N�<T_=�cżqߎ=Q6�;�D�;��]�۟o<�i0=�G"=�D��aZ�J6��+
��_I<������3=6��&B	���[==��hH�nP{�h=��Y=b�=�"�;+���R�g=�e��D��<CA�����}<���<�J����w=o6�y�$���'=��=�E�����1��:�_�<�*��kD�<�nL==�<!�����;�T7��A��J��iB��,��O���R�؁�:p��;<X=x,�;�\d=�݀=2=�*;���Rlb��-�
��<��&=G퀽��̺��HJe�<�9�<�㼑b��x�`={�Ӽ�=��p����������<�R弈�=�:�w�l:���<\˷��K��3<q� <�6��=Y=O	�Q/p���;�r=Ҥ��`�<�-�)�\��;	��<�d'=���;u�<���<�	�<Ec9=�a�<���A������K�����Z<�Ԅ�� I��H]��oP=��=S}��Y<()G���@���@=L[�<AC��� =m����I�'=: ׻��u���K�<?�t=�����c�#��<�O�<�F�����;�~=W8�<p/x<ò]��2�<1i���J��T�Y�W w�E;=��`��)=��-�@��<?�j��E=�D޼�VH�⒲�C�1�O�Ƽ*v[�ݧ0=/�M<�E8���<&*-<�K��J5=�$@��~ڼ�p=Σ=�.�<׋�3���4t����=���<v^K=
^���T���ּ�ί<"�7=U�M<�� �b֜�#bb=�<=)�^�&�={��:rt�p��<��3��X=m�D�V�I=��A�_�&�?�<���&i�<|	.����<&iM�Ѫ*=&~�<��=�������c�<zA�$9�گ_<g6;�*�v=���:g�+=,�d�ni<��J��p���ƒ��z$=����k�<�|a=L�p�#��<:�F<��>��<�,>���ڼi��Q{h�_��0{�<[)��?>��3=u�>�NLh���D<�= Aļ�C�<e���¥�Q���I�����<ٱ<=�-�<):%�/�g�����.����<�ջP�K�$=%QJ�b�=8o=��^�	�y�������)=�4M=�WE=H; �~����������<��ׂB��=9�<�a���F=L�����>����̣%<���<�}�:���Ɔ=Q�D��T=@8o<r�=�=�����7�1�=��*=���OdW���_�ż2q7=!1�C��<�������;/p��<B=+'�<��R�`k==TX�;輮�
�ٌ=�>� �b�=?<=�D=%\`�������p<��+=��<0��w@<2�]<b�G=5��=�z�<R�i=���"��N��ȱh��d�[�(=�����A�< �v<�ҧ��y�9������=�	=��J���
��s"=u�=F�d��M��w�ʼ��
����׸1�~�����<�7:�:�\�&	=�k=o:u<S=�5b��n�<1[���=�<��:�J����<�=ۅ�<ɿǼ�C=�����7żK'��..ϼͼ�-G< #{=��!�A��<:�;,�]=��	='�������z�:��D:lh=�5�<?U=��4=�lm;C������#���ѧ��Q{<�N <�T�<�)=���<�6=	�;�L�;��=7(������n$A��G9=��� �=6V=
���~7<��?�LZ��N�ɼd^��zȼ9�;h@�]c=�����-=��;���=<���<oY�;�+U�KYy��W��_���z�<��;�^;�'{A=9h�<v����#	<v�5<���pb�< ~�9��N=������ ���?=��<M F�L���G>s���T=J�&�X���'�1���<��<�}�<�jE;�NH�D|�<h�d�]H;+�u��'7<��K�!X<�br��8����P�=9	�%�5��q�;{+=��<�<��P.���+���=�s�;䞀�Ȏ	=���)��:M!=�=Z:2��B<:71<�VD�S�<w7s�'1'�{���� =�-=��;����l��<*=�g�<Z���b�ms�:.�#�8����<Z���^o���4=xD���l�:ʤ<s��r���C�'�T
1�~�<B�:����i��]v`=��;�N��2�<;�]=<��Ә�.�(����,JH911~;P�����;@�=yI=Hzl=��<~}����>=Nȓ�)}�<qѐ�
/�p�`<�p����;�f�� �<9�D=��t=�⼌i�<M�;�%=� ==a��C���F���!=i��<������<��� �H=~�]�3�=�e�_�,��3�=� ��\=`pg��MT�n	��x>�=��<��>�+ߖ�ItV=�ف=�@;]=g�ͼ�'ͼ�;t�fu_<�<�s=�C=�5<{��;�ֈ<�$>�U�h=`h=\sk=� =�q�<@I=��<��	��6���=� U�eS=��@<�	�<� 7=-�:��=�ט;�~��T����\�3���ڛ�Ǽ1���=�S���6='c߼�`�8���ּ~S_;�Ad�M%�v]&=M�>�V�7<�k��<��=?8Z�5 �fO,=>X����;��;��q�M��<Z����{Q�e$�<i�=؛b=���<ʺA�Zq�<~�)<�\�<ʖ<,f�<޳"=a�J��5W�.Mm�l��!�I�����u�׼↡��Dn=��;�v[=�B�)(���h��)�<Re�<+`��iCD��M��oi��rw�~�b�F�<�1���p=5��<r�G=���<�==,���e����[��ɼ�3�� ��<�h]�'�2=a�'��舼�~=g=.C�9�)�;
C���<����M�ں3J=4B޼��T<3�;t��M9O��ힺ�v/;�g<_~'�kA�!��<��;�я<q{%=j-�;��@�J'?<��5<���<̀��~�<U}�<6c)�H�<0�k��b@=��;�=Bc=[��<�P=�}}�Mf<=�'�<tM�;�6��Y�Q�����E� =S�5���$��6=�t=�!:���!��<|V+����J3I=.�7=��r�S[=1�f�8�3=E=Pg'��=���<';U�WB�3��y�*=�~��X� P^=m겻w.ۼR�== �,��u��vWH�jP�<A��Fb�<(�*�Ca3=U�(���<�<	�=T+Y�
��	��;osA�7ݺ� �*B"=�x'���'=�@��`W<�Z��X�=q}=��&=3�8Þ=�[l=�)�;jBϼ�jռ�1=����!�3�n�r��<�.=�M=��\=�	����;��6-=|�<���<��ϼ.*=�^=��<<�B��t�<kp1=9M��S,#<zf=��=Y�`=/�:��3�<���o��<�dҼ`�ٻ���;.�㺮�^�J�Z=�%�c(=B}��o�<��/b��2�����=�ȼ��=ʩ�����!�H��ϣ^�
̐;ξ�I\�<,1e=[>@;H��:;(�,�\�
��<��=H"=LZ�=����J��X߼kl�#�;��!���<J	><���"ٻD2j<������<����_=c'�5f���%�<pd<	v=��a���\9V=�\J<�܎��<�L�<����i?�<H�=�Z?=��=Ώ"�"�2=iü9���2l9=�����)=���;�[k:��'��|@=_��<_���K�<��H=3U=��޼�1
=��abW���<ۉ�<^���Z���=դe�W=�}&=łǼ;m&=ѧ	=B�;=�w���] �3 �5�L�<[-_=�h����sH¼I�������<�G��� <�Ғ�Zs��pÌ����v#�<�/I������0c<n"��x��<�ph��bڼd�������u��y����3�H]w�	�n=cF=� >�V��<T�=���<���<k�=�Ui��N&=H;�<vK�<Bs$;������!<��7=��0�D�;oO=!�5�Li3���S��.r;�e<�r�ؒ9�s�=�{�:9�i��
��`Q8�t�E=�,��wP=�!��^n:��s䄽m�?�D)��8`��z<ꔼ�L�=xa��6?���E�0�o<���;(꣼�dE�nm,=/F=�=�B����;n�����<�q0=���;�is;�r��+B=${J=A]�<``��导��L=͋9=O�R=&\�<�+=d��<d�<�Z�O��Ko�U��<�>��ȼ<H&��9�E�������<7��<|�[�P�<��͎��!�R=
��=��];��t��[<���D=��'���<�"L;������û��}<"�Y�*U=w1��?�r	1<g7�<k�=U
�C
<t��<*�V���:�W=~'�<͆1����.��)���m=_�
=./�����w1�^�h=�
u����<'�	=�+~��6���:����6=�
�<�񝼕j7�9q��0.���f��跼.��$B�<��=�9�<Ӿm�ͷ<�C�!Ծ<i�<�bY�F^���0=��S=���<	=�<�{=�q�<����i��w̆<�^=X�_<`@~=�=M<�[=/��h"��'�<��2���(��U�hѼ~��:�z�<~z%��<g=��6=�<�����&=���
e>�&��� ��tR����.<�e���Y����M��z<m@�kqܼ2�:�ޭ\����<g�׼�L�<C��W%O�#���S�F<hB��jr�Ŧr���ԼWb,���_<4#�<Iph=�9D�h	><��<������<j^��Ữ<ܴ���;2@=A=̹+�$�=�c�<�,�F�ż��Ѽ��$=��F�e{o=]-�<b�]��L}��&1=I��=Tx��F<�	%��3=�`1�ax��	:�UT6=p|0��z$==��bq����=��j=���O<7��D���23�<G��<:�J��<V=\C�<>�0=���B;q��l��'mӺ�2'������D=���<�:d=K<a<U#��r���?=6�׼�u`=�[�<y�\���N�U��<�1�:d���)�Ba���	�<�í��[R=\+q��X=i��<E�&<���<�$�����5�<����G0�<�G�������;�H6�ƍ)=r*��,�<�2��j:����хv=��ʼ'� ���;�	)�&4U���0=���<��Լm��<>�<!�6<���ٞ�<�}<��<Q-м��*=&�I� �<�'=�*�	��p��<8Rٻ�+7��0���$�;�gѼRe��`�a:=}p�����H�<�
Y�5#=��4�=�t<*���K��\�����f^��x=TK�<����6� <g�#=G�<o��;��߼���<�=�g��揁=�=�&��_;�p;�h�<-��b����@=�����_��{J=���<� .=���Gv<���;�V'=�_G�T ���=yW��=�)=��Y<�K<)7�<��Q=�z��*��=ʂ<0��ĩ�<Wt�h�:=G�<Hs;��o���x={�/=�te�1��<��ۻ�0���Y�#����0L��]5=�?=i�%�Gܼ.*p�g�����=�Z���!=��s<!�I=�e��/�=�
<F<�:�<h�!<�K㻸@d��1d�qѻ��C����q�����<G���`=��<��+;V�f=��!<z�|=:໗*H=��t<��P<�	<��<�L�N�=ȅY=��.������<�l�<nG
��D=�C'�x�]��x�k�@<>"=�Y�o�\��T�=ȃQ�d9#=Ja
����<���L�=68=w�<�%�Hػ饔�9{=9��=���;BKK<PR��=�<��=�K<�k<���<O��<ZG=������=����X=�Ǽ�p���tE=sZn���¼]�B=2J�<� �5;�*A�W� �
Z�<������HG=v���X�<�[ڼE�.�{%=~�]�M0��	3޹��l=~=��P;�O'=�M7<�Bk=��K=�!��hw�;+<�b<>��}�4���Y=��=��O��I|�̆=|WL�?��<�-l<�4�(�b=�8"�Q~�<��]���=*�ϼ0�<��Z=o��;c	����$=��Լƨ�w�w��(�<�q<��n���N�ة[�����k+=LFL��ި<���<g˰<�Y�<�D��E8�*���e"�dW�����<�W�;%����; �x�>6=ĸ�<w<~ͫ<�ve8]�8=X|	=q�<Eǿ�es�;��;�Һ�)=&K�� ���h�<+�|����<r!���S=��mK@<
ʼo��<��{=�`D�->��R�]�ļ#'��B��?��<���9��S��<t	�;"%h�s�=�q~=�fļ݇c<�����,<�[�:��b<�"Ӽ��Q�<��4=��<K��<:O=.>N=��@
h=]�F=lHƼ����<��	=�¼�&/�MĊ=��g��'<�=������<B��p\ؼXɑ�j�=>ё�D���F�W��f=�;�����}o����<u�T������6�<Z��<�&t�Gq =!G�;-AE=��<���k=��a��F�<��h�t�ϻ���i��p`Z=df��Iw#�M�`�^c'=pD<�=��-<��=@'��FS*=���#`껔J�<��o=��9;ºg���� =)�<��<���<F>=�tĻLr�<�a��Ԃ��;U=�m޼j�]��2���]�<�:��R�����<���HP@��*�<$#��Y��̼k�<��=��=��C�[u]����<��V�VG=U9=�=mm-=� L����;�\��u�:�\L=ֽ<ة[=ݾ�<̋�<��x�G<XG���������-7��
��b)���p=�I=�5�<T�^��ʞ�}i_�ݟ��y�y�s4';
X��C7=�Y���b��&=�h6=�[=~DM�������|׺�m��<a���=�<��׼�t�;���s{�}�<d�L��=A�������]=�0�;G�=���8<����w�<}od=6# ��e<��i�>�<�a�k���*<|��<>\
=��<&Q=�ͮ<��=,��:-�ټ.��<��3>%�jl���+B=/>��o�;���:lR;d����[=�AO=�2�<�V=,6=a��|���<E�=Ŏܼ�)��9���f=�@��o�9v�Ѽb�W��=?
E��'=T��<��=X�k=�n����2�	D*���=�ɚ���<�P��(���Z.�zE,��������9�=��;��j=�9�<��N��7h9��(��ı��P9=�>=����]<<v�O���X�<�� �!�H<�6���Np=�W�a2�<_҆���?���<��;��=SPR��J�;����W��<	��.�7=�䓼ځ���ּ���I��a�j�u՞<��ؼ���}&�8���FV�<�X����<�ě<�<�)��	�r��YC=Y�T=bڼ��:�{7=�����7<�\`��0�;�w�;H�9����<��E�������,3�<e�<{�5:�M9��Q{�B|�<���<�6��v���>��0X�J������RJ:=P}$<7�=� ;�	x=3��8����:�#��+�J��;�=�v<2�:<m1!=�	=nE=g������;<�~���F<0���t�2=�����c=-iG=��A����<X'�+�Ѽ�t�;�EB�@Q����1=Ϲn=���<��#�����߆���yB=h��<��N�fs=��=�eJ��;���6�<8�<�N=?��<$�+<��/����<z�"�p�?<�G2����<��T���ɋL<t�켆`��d������mS0=��-��?6�!i9���Q<&��<��;q���(����<���;�X���=�2���u<�J=�<���z�=��"=�u�<9hG=�=��=��9��=π2<�f=�3���G�|ʠ<7uŻ:�=p�ڼ�����<�<"P��o�z�:]���Ƽ99����� *=�J�<6J=���<�7=&Q���|=R�����U�A=rZ�<V�=�|<m3<3;=��<��1�z; �G@=�S=��<�hh���;�v��� �������<�B��L=���<tFz<�R�ꢻ��=��;�Zm=�κ���<�8��\�5�&�=�|ۼwcҼ�I<pH�;#8H<S%<$��<����%�7���`<��i=�p�<M�����^�l��'�>�=������L�NR��~��;eW��甽$d��1���?�<]��^*=�zʻB��x�<K�=��;�O����<}�˼�^�\B��ֱ�;nv-��a(<rv����=���d��9v�=_�><��4�B�w�-� =Jq<��H=Iu=>��;����=�b����`�<MP=IH=��,=���g��=t��<Fh���x��q<�W=}�3=�hy�2\*=�?�<>��9Ķ��˔�<�ǿ<4M�����c��<�G<x� �*�
����<)��d�B=|�l�JT�K��|"n�7�4�'�<X7=�>�	1c��G ���+<u9=h�U�*�"�</A=���;P������a=d =��^;��I=�@��8�$�E���	`�"BV;�==��=���u���=d=�r�;���;F靼fR4=;��;�
�<U4O��8=��"<yL=��<�f,�ܞ+=z���<��ټ�Z=��5=@��"�d=�JL���);��;=f��s�r�qn��E-�HN<,�=�����<�B<�^=T�5<�r�uG;��5�<������w��2T�l�=�7�P=��=��	=*[����t<?�I��d=����t=4�Ǽ���7�k;;	U=)�0=9^=�;Y�ic�;fj/=���<��B==������E<{Z-�����3�mV�<�pP=��
���߼х=1�@���<& I�1I�z�<�=a����<<��6<�\�=��>=B����+��<�<�K[;�f��v��"�ޣ<{�~<o��<�Cv�r�����<B�2���<ߎ�<������84�l�߼���<��N���W<���<C�:��4=&�*��?�<�š;%���0���;�*��e#<��ȼ�|I�ԁ�;��;���4<�Cz=��<k�_����\X=�X=О<�tM<u
=CJL�3���ڴ�k =E��;��={O��3����<E�<�/���\�Z]��r�<���<���:�U�����=�;����ⴼ�7#=�<`�Ƽ�"��x<f\&=���uY��Ԣ�3�.���n<==A4"=��<�Td��@�;>�<��,=B��:m��<��Ǽ����02��?}#=�e!=�t��4���!�-�=�H��2=;�JTm���e��7Ӽ�����:�O�<�?��x=���z7�e���D��$�<G� =��<��V�����`�TO=��YL��i�5<)�@<�:�|}�IԼ؁��\���<��<��:�닽	jڼ�p���<��N�?�3���$��t�y��;��<#-f=b��<�Rf<e�����<t��ҿ���ҼH[)�`.���=�]h�JT=<��:��y�FK�����{A�،<�&_Q�˖���#V=��S����<��f=i���E�v��1�<�� =g�l��.Yo<Z�i=d��<v"��Zf%<R����Cr=K�<�L=�e	=|��;���<�U=��j� ;\>Լ��<a��Z����<p�,=
#:�<uw��ţ�<ËW=���<�B���.<�:=��#�<Ҡ<=���1P�=ut�S\F��2�Tqt����K	���S�,���	J���Q=� �:"��]i�"c�zsI=y|�<��=aq\<��K���c<�0=�H>�j��<�y5=�0�_������7/	�Q�9<�%ټ��T���s���� "�< E7=�`j�S��5����漃u+=fY��p�����*\Y=���<nļMr4=�K`=��<L&0;���<�6�<F<�<}	ȼ�TF=���ӡ����Q=�e,=�K» �!���>�ى[�`�˼��$� ��<}Na��w���9Lpd=Z/P=�"=\����O=V����.=��<*1A=p6[=��<���<Xʡ�1��M=�l���D�L��'���!���_N=��r��qW=��&=�*I���2����<��=�:�"/��$�]��cX�qK=��\�&�]�.��<���Q���4񺼇=��9���<��T�f�=��<xݼ�C����
���1=Z�;~�J=g�=��;�j<V�H<n�:���� �F=�=�<?<��<D�.�R7�:�~H�_S�Y�¼�=�J<h�(��u<n�b����#h=��G=�������	�ָ�E�=8Va�o�<=�}+��m���j<tӾ<
�L=
��^�;= !�X_Q=hr<��<�oh4�3�`%r�G�/=m�p���<�*�7�<��<%�<��'�5��<$+��T*�f�˼%�<�P�\2��|V=&�6�(Г<јP=�g=o���J�w��<�.=w��Z�<�⍼�@�<Ñ��E�Z�D�鼔�J=�W>��Տ<M�<=�r�m�j��û�W��q(=��ļ*�ѼW�^�&a�=r�?=l�>=/j���6=r�<�a<E|�-=���I�<�N<��Հ弥l߼<��<d�=rY�<�;�0[J=����d2=�r弌\�<&��<J�F=��R&=%�<"+�;q|�<�'=����\<���,=�Y?=<T<��(D�}�A=w�����I=�.��9��<�׼�}����#��$�� �<��<I���uo�9U¼�^�;>I���;=��� Y�ЧJ�r��;x�<�fq�|�!�]��S�n=(r�/C�����<�fk�}�E�h3��)$�F�����<Ű?=���<�+����l �h���)&�;�My��PR<��"<��x<��4�wC=g�ؼ)x=Pϼ2�F=�	�&���`�b=2��<v��<�9D�ʭO<�����#�� ���#=)�j<Uo�!�����r<T��;XM�<-�<���TN��g�9LuI=3�<S+�;�E���g=�e�uټ���9��E�j���<��<�1>���ڻ��=��f=�&�����:^���  �ip��.�C��@��5�,=��@;��<�����P�	s#=�=����<*	�Ee�=�:=E��;fٹ�]n�<��=�y�5�����;(z=��Q=�R�<�ָ��
=�s��|,���|<&�<' =_��𕻖� ��Z=��<����1=�{!=Ŏ��}�<��.���<@^���ndO=�[�<�탼|�<��O��`�*V�<�?=��K=1wz=��b� ����༲�����¬�<]J<�q�L<x�=�M��K1�n�i���<}�A�i
0��e=�!<�7�����-�O�=��<{�-=�;P=~�k�r,߻V�<�kf=6��;Y=;5�3�Ga8=�i`<�i���=&h���R<8�ͼ7_߼��K��Ɣ�F�=X��>�<��Ȼ?&��_P�ķܼ�鼵�V����<�N��&=��E=V���_�JS�%=��2<%B=b �<c�!=e�1=��)<ݜ�<�9=��߹$=�$=c�{=�9D;��c��n2����<�ͅ��e<�Y׼����)�7���b='�=�=F�<_'��?�<
=1�̼��A���Y�R�/<�-μ�k<�Mb���;��<�,j��><�*|K��i��aY<BS=</��^ZP;dY����c=0N�|�6���v<Wu�<��<�=g��<�p=��<y�[���"�H=$d�n� ���<�f��oYs���?=���<�sy�#O <�I���<���CJ�;��� 5�<1�N�$�<M��;��t��=_��m�=|;=qp뻫M�;�}�=�A=���<������=p�(='b,=@%���:��"�ĺA�<�C��٪�M�<:�<r<໗�_��/��.;T��D=��H��u�$5I��\�<�r����\��X=��5���<M���&=ݙ%:T���E�弗�9=H��U�<�5�t=�:<�=�d;=�-�Х=��X<
�;�f<ԜB<�Mj�e��P(����ἡ�%��i�;�[���x��G��h�*=�,������o�o�p���1�e=�z:=Y�L����R����<}����B=��=�:��>H�n���{	���L��A���6�;��<T�z<ͩ-=0��K�Z��<^����^=2�"=�꼞q��G�H�#����A��r/���)=~ �<�ٻ�T�!���c=��<9֐<T��<"�<<����w!�j09�/s��H$6���M�=���V�5=����g�:��=kR=�I=*�9=�x�<0�=�",=��<��S#�Y˦<¥n��ad<�^f���ϼN��;���ʙ漙uf9�ɭ�q=p^��?s�p�_�6=ϼ��"���������<uq���<�ɢ�ahz:�g=u =�I9�2�=�cI�,�9�UW����<O�>�b��;�$Z<�O$=�1=���'Ri�n�ɼx�c�?}�<�q�>W�<��=��@=@�ڼ��[=ĭu<����'�6=@�d���(�w�=���(�ʻʊs���P=1� �g�9��<Qu.����<��9<w=�O=�z<L��̓�;lq=c��=�#�2=�W༬�@�=��9Lv�vF=\��I�,=ǑA=ƫ;=w&��9�<k!w=Cg���^��};N�}�x<�ʼ쪜<��	=��1=�ש<�=�l�<>�<�=�q=�N=�X����2$�<��<<���<C[������6=�a<hY�	ߺ<��?2�̾��f�;Ps <T��OC�58�ߜغ�?���cP<�����s�:�L;���<X�=��[=v�\��x�=ߚ���<=qv=$�"�{=�r=N���NK�	TL�ڊ'�j��<#��;V�=����_2=�ϝ���={B!�S�/�R�$=z�g��
B�]��>o;�.��$<#�@!�������;Vr��2O=����(����<@J0�VH�;w�=ڹ����7���c�S��a�r<U�k<�ah��W@��j8�5dd�=�u=��μ�&�<�D<TӢ�9=�Cn�������U�r��<��.<KGm=g[D=Π;���v�-�	<���;�A��P�26���r�<���<'s��á���G�uF�~Yu��؉��Dl<��I��0��(2���B=��%=��j=[1�K�=�"�;S$=�oH=hqh9<:�<�{�;���<��<Wg2<�OK=� �� �a��:�JO���z=~��v+=ac�qD�;�)�#v<�/�<AF=Ty<X�<����~ٻf�m��Z�V�)��C=6�ռ�F{<���<�V׻?�6�>�<e	��k
�_�<*� =w�<R��<��<3/�<]����&�<��ݼ��W�r��<~��.zS�<Z=wL�:� =�T=a��OV�;z��<���FW�<�X�<S��=*i�N�z=�&i���I:��~=b��v ��RQ=Z�= '�<��݀��Τ<z���n����=��=מ*=�(@=Y�8�yx*=$�2�':=���<��^����Es��fj<�p*=�]���W��ޫh=1�=���dӼ��A�ю̼L	缰�.��hH=�{.=������<2D�qe�<�6�~�u���!�¢\=��6=;��g\���=�_`�N
޼8��B���C&żH���+vo=3o0�c��0(i����7<���	 a� �2�����R=�==?&d=<�l�!�=���<��J=�U0=�{��Ho,�у'=�'=����<��I=$�I=��2��U<%�ü�켡:Y=�8A=:�i=uZ���w#=U=*;����?�YŘ�J�P=;�����"=g�<T.^���\��}�a�p��s��F����=9Ư�#�;Z\'�'�;z�1�%yc<	j
=o�#��5��@�g<=B0�/+���Vڼ��-�c�=��<�."=R3 ����<��o�}�A�؀�����<ud7=O=�hR=n�K=�=�C=@5�͜߼��!����<�`=7^��Ǜ<qX=��<7K���ɻqi5���W;�=��������I=ho';�m�_!=�u��zq<�����[=�Y9�HVl=Z6=����ƻ�x=��=���<W�4=�,=�K߼c94=��+=��"=wq<v+;rX=���<����<RU+�3r\=-p����<|ӏ;��a�%=;KZ�Z5=i1ټ��ŻY=�==��;[;�#@�;�w5<�y��^P=b�>�WGD�(~=�V�,��=�,�<}��<zsa<l�ϻϏ$�;��<����;��;=����,���	"��K=X;=v�9�&��u�4���R��($��< =Y�<	3=�Pu;+,d<�3=lW���h�;�O��@`=����m=*Z�=�3ջ��=II��(=э�<�r��������$<k?ռ�
��#˼^�U<.�=bÀ��'Y=T绒�i�"�0�ω�Ä�<��=���<�ɀ�o3�<�Qǻ��<|�=&F=xQ=�8����Ѽ�=�6�e���ü�NW=�ʫ<u�ټ��-<Ŵ6���<f�V=�g�Im<�F5=�ٶѼiY�OA������>�,Q2�i�<�E&<��-����<cm�_�b<~���t��;��=]�ؼ)&i����<�J��ƭ����<�o�;j�l=RLU=Q=kF'=��!<@�<���q�M=�	��k0=�q`<gC�=&�;=���=@����~W��D,<i!K=g�)=��=���;� B�Ŵ����;����������'=�==�==���<��<��]���=�=�<�]=C�4�H�&$P< z��*0<h��<�=~��sPk=l��W���"��(@<B[��Zܲ<7�����:��<��=�Y/=��<���=��<�1z����~z]�����t��`����t����h<�M=��n�Q�J��q��=.����.��$=q�v�/eU��PE��0м���<fF+=��)==Of��(�-W�<N�<ᐤ:�_1<ߤ<��N�yk��fi&=P��<�&���y���<�%7��ao��4$=���<�f&<�r��8=z	8=�ؼW�D=`�U=� ?=�M�����k*��PJ= ��=| >�ӂ5����Y'�������R�_h��ז<�t%<y�<bg[=|�]�p=�<'�=�K=Ȗ��!;�f�<��~;W�⼀M=��M<+���/��`�8װ��G4�<d�0�����H���=wӼ;=�.5���M=�=�*�?𲻖z��D����=U=������"�$�����S���ºa�����Q��i8<K�=��H�e<MXe��!����k<�7+�0(
=#������=z�(�&���n�酧�B����oc:������\�*=m!J=��'��"=�5C�e�<A�<.�,���q<MT˼������NƼ�n�:�Cr<lZ=ی=����wx<�Qk=�u]���*=��~��ea�tB=/�,=�g=�w=�q���;/���fo��l�0�d�4�2��<��wx��UMh�K+�71���A=�3X;�=(<�
���6=��m<]"���=��ټK�'=�4��z_=K8E=�J�<�	P=�������<�(==�Iڼ���<1��<˵����X�,3��$=�T�[�b��"P��+5<S�N=������nE��.�)�@��<X��;Ǟ*��x ���o=��"��'����v�/=���<����;ؼ�dü؀#=�}9�,��^�%<\G��Оq=L�ȼ5��b�@=�yd=Y'�}�L;�O9=�켠��K�B��U=\n�x
�<0���4�m=pM��@'��T	=�~,�I2�;ā������<�Dƻ�2s�Q,B=}¯�G�R�� �<�lZ=�	��{o@��"�;��h0E=:<�|�ؼ$��Z&���c�R��ڈ<MiO<w�7�#��<}�O=�!��L��8���?=
)޼�)V��.B��B��S=�<N������[=U�Y= �<�Rv�����^�=��=~AP=N=r���,�<W�<��<��o�i���`�A�<U�<mC�;�R���"�;�<c��{��<2�<ӌB��Q���W=_2ϻ�?`=va���m������	�3�<���~(<�C	�<cW���V=t�<aV}�5��b,��m��:<����*��	J(=	#�עe=���Y�G��P:����r�� ��<MV;<P=;H�<k�"<4�<B9W��=$��;��
=�s =@!B������;�~�˼��N=y�C=���<Q��;$�7�	�N=\4���J��k7غ�!���:�Ax<
�ϯ(=	%�<J����u�<�,�<2]�.ĩ<]"�<��><�=���lϻ@�F�B֋=#�<����gG�T=a�=`�H��-(�;�̼c�R�:r��5�<6"B=���<�W��??����=�%"���~�F�2�����R���5=�I�\�<U���n�O��ڟ;�D^=�i"=5���r�<r5�-~μ�$X<1EH=J�9<�i(��C�ߟ�?>z=qԆ<�HL=>�G�B�*���=�=_�H+=R�e���=H�G��c/�gw��D�]��U��q��<@�]��uüe�ƸR����4=,&ļ�o�\�;��Iӹ�Z�@��=�;��8v\_���s<�hR=��t<������I=7/��Xu�T�D��Ｙ�S��K���l3;-��<?�K���(��a���� =�sA��=�n��i�o=�2ڻɀ�<������b=֯d���9=�}|��LS�_?<��P=0�;`(=c�@P�!�<D�O=�1�<h\��� �d!���c)�b&����i�<�	�Q�	=�8='s����58����5��*�<R^�<Ðh=��=�g���-=�^�� �7<��<���3=���Fo��m�7�c�8ٻ�J�V�Y=��Q<�*=���Z9��聽d"����k�^~��j����9C�T<
�=)Me=��=c���1�;�l�;�ּ�]�>6u=YF��@g�G>�<M�=Z�-�V�<�O����<2㘼�C��:3j���ڼfo2�\"�<�j"���<fD�<�i�;Ց!��|=��-��|<��-��	�<��G=���<��$<8k<���~�<���;��/=��W�V	���K�;��=�������#�<̓<^f(��=DP�)�:��zK��q2�t�=��<��%=�,9�8i����&6=��`��=[����Ѽ!����O��tT=&�!��m�<"�g=_�!IA��l�?���w#=��5=�d=~!6�h��:�=ѷ=g�< =@�<��=�E�;5D�<ㅍ<��8=�Z;�h<y�;px����:��;����c��m�;��Q����5'Q�J=ڂ޼0�P=�J�$K�;��<�(伭D�~j)�(8�
���N�<>�===��B=+�U����<�9=��<���;&;x<֙���;�m4,<��~=CZ �<=�+o=$���c_�s�H=��^��K�,/=D��5E!�9������=?㦺S��<�r<���)<ɇS�v���< 
�<�{�;�(=;8o�=?�=�S;�L�<�˂<��߼��L�M�q<p��<X�m��w��`�=���,<P�=<�� ��S=�E�<���;�[=�[�����P�=V�7�Ŋ?��G��z��<
lN�vT�;Hw麏��9u�f�f�H=�=�:���<.����AE=� {<�=91��<�z}�<�r�x"= Z]�~0���t#���<%�;��M=6�<��<��R�#v]���%�]=�a�=�c�<u���p<+#�^��<Q�<&�3���,���
U�=��<�gp=`�b�9�<���;=cl�KK=��ȗX��{6=�R�H�˼QN-=��3;�m�;�Q)��[U��X8�+�9=:d{=��=�<��O�G	�;�MK=�X�<ܖC=�ͯ�&)�<�>=!��<l��<��������+=�y����=��(���=��-;!H�<qO�[CM=m#@94�޼����^r=��99�u7��<��<������f��o�<�y#�9N��g=K��i�_=�]:��<.>=>t=��P=9�P��Mm;Dy*=���:
�4<������ƼCt^=�[x=s�I=��hh/=U^2=�=<\Y=��Y;֛����S=k�i;�݈���=�={I�<.���fW<`|F�XQ��ڦ�f]�<��A=4~�<L�>��B������li�A�;#���6�"�S�[�˚�=��<��U�|�ڼ�I �4=%�<�.@=�X.<��=⡽<��Z=������?A�<��4�P�=�y����:�
2=��=��`=�<�E�;��A����<u�S�c������rEG=�����<A����'�����
�_=����X=�:<3�������'%���;d��<�<t*F;��
�3�C<�u�<�3?��?I<.��=굀=|{@�=�-���:��=u��<�L�;��=��N<4==AE=�=��Ҽ�=���<����'=�� ���l� �Nmg�wM����%=|2м�@<{�¼�l'�p�={��<�����<ǛI=�����M=�C�J�]�� o��Dü�f�Lo���<M ��,�<�	���&Q����'���5�S�ļ�fP�'�=߼W��|�z= _c�f�.���F��'�<�����2�H�ּdp��>�����,;�LR=��~��}=k�Q=�P�<����Ъ���B</[I��~<��=�b=���<��<]�߼ӱ���;#=292=��I���<kb=ȷI= ��ܼ~��F�<�>���=��u�A��<�(<��@������<��z��S�1� =����}挼A��Hxp��=���<r�2�g(49͆�=ƪ��p��<X��
�<=$�<�L=��<�/¼Y�=v�{<�,Q�z�>=�����pV=6�;Z��<+X*=NVм>K%=�`�u�h�	3�<�����l�;7*<���81�y��<ԝ6�e=�+�:OM	�O?���b=y�i=�$6=V���/������=�<���˙m=�F:,>H=��A�UN����=�Y;Ԏf<�3ڼߡ&=�9�<��D=c��<�X�QB	�DeV=:��<�m;@:$����<�=kr=�cT<�*�:b(@����aH5�//=<H?���R=SA��ۋ<��C����<��V=��H=F [� z`=z�i�j�7��Z-��Z��uDd�fB�<p?�_���C
�]f�т�<�L:0��;�;<�JK��W =�μ��<�������=D��uO=BY�<h��<S�<��f<k���X�<d-=�@6=zo.=��=�=�����9�<A��<��üj�P&=�
�;�L�<|����������q߼�_^<�\>=�(=��ü��==j���Sro�Ǝ=���<P{<�􁺻�=����Ȼ�U�\�<hkO;�6�gg_;���;/_�<�)�<�j��k�<��-=��<���<�n�
�^���I=�i8=|���⽻�b�<S�<�sX���}�!:*��<ϭ�;�*��������v.��:=�W-�$!l����}>=
#�O�ʄ�;�{�S��sP����3�<i���<q��<C�����LZ̼[�<�N�<g�6��7<�nһ,�	�Q=>�C=N�Y=�Վ����;2�v=0x�<�$G�<��üg8<=q�;Y�,='�3���F=�g��p�������<8'�<D��<�O;�����<��}���;�}=����M(
=��=�E<�Ya��.=�b�<���;-$�<;�7==�E��
#�V{�Ӗ�<�;\�=���9l1�= ~=$ =����<?Q�8��=��2<��y;��=:.�<:��<��<��;�L�<�G"�M��;��W����v!���4=��B<I��<D��<�m<�̀=B�X���ܻ/���H����.=��=�e��s<=��Ҽ������<�=��<�=�?+�;3�'=4�V��9R�@�L=�	=�o!=Ls�������<��7�}&~��5F���;��%�=�(=�伖�N=��e���X�<��A��S=6�n��#�;gȯ<~^��q<=F�#�We ���Y��8�4�j=�m��l�r<����z����J�=2��<�P�Ux����;���<��G=4�7����<h#;k�<�[=�Z�����;�}���3=�+T=tj�;��弯�λ/y:=IJ3= �;�cC=��5����<2
�c�;������ߠZ���"<1{=z.|��LѼ/8�r�4<c~�;�嬼ȻH��8��X=˽�;HaU���<���tB%���*�v�7;P=��٘�;��<{��<C\-=		��g�;�r(=M���N�䳮<��=~�D=��6=�=��.=s[=���&�1=��i<��M��OP��r =�S=E;<�5?=��<���<�dl=9�<�m2��<@�)t��0�;��<�e;��r
�����<�㯺�V�<ث=��`��M�<I;��9���`��=�,u�G뼆��;�e�?�L=�n6����:��=&�d<s�:`��<��r����{��;h.�<ݾC=Co���M�QY�;�+=�뱼B�������/��Y��<c�=�:=uv�<�h�<�G=�6<�:h��
�;�(�<kH)=�=F="
E�
3���A;��%�������1�YT=P'E<V�弻WJ�'3L='��̐=��=;�[��cl�;��'�.[=�w<�OG��4	�;�+<�T�H= C=��<=�Q$��N<t��6�<�$=-ū��kZ9X�*=ğ�����<৽��U=�L<?�<�o =�K�&lͼF	
��0=�+��ٜ�;nh�� �<�;<=6#�<��=<�$<ʯ����<nj �-=r鋼������(��Ī��#����=�m�<W��<��4=�����V��6{G�&S;�t�;�K�=vb6��c�;_�<�3=��:W�!�*$�L�==��=Ki��A�=��t��<�:�Jy=)�z=�ꊼ*Q$�'��o�����r���˨�7l��o�y=�4�<N�ü�M@=v�I�':"�"��ƌ����7�=�y��_�)PN=��(<��*=Վ=��1���ϔ�|<="�P=ԁ:�b��y�V�K>"<?o=��ἅ֒�f_�+S��K=p|g<��{����<�*�2@D�M~���`<�/V�_?��b�=��2=h!��ˀ;�:�һ����[��M��L=�<� f=RK�<J�¼�=���KP���E=OeT=��j<N�ܺ�k3��
=�R��(=����/�:;<���I�;^�!���A=�Y7�׷�3�`�$��<6-=#l�;�N�[1�����;_�<�*��+��̬�HO<������Ҽ�	��/�K�"=?��J�N<E�߻�J�H]O<�ܯ<��6�� ���-�rY��D��QX�@��<��L���<_
�>8r<��4=�陼�	�5/����G=(4O�ER=�)M<7"=��=���M��wr=�5=�3o<�@=�#p:^�2���k����<*IG=Ny���Z�og���Ǐ��TX=�4���lܼD}����?����;I(=t C<�5�;Ͷh��'=���r��<!��<�g��N0<�P&���2���<�
J=�8/=4V�<}��sv�%=� ==ԡ0�:M'<��i<W���H<���;�I&���
=� ��҈U=f����n=��2�%v<U�=�u=�3=l�e��Q���_�s��<��j=�mԼ~���#K�_#�<��*���<W�J<=��<�&�(�=̊��=\;�W�;w�<N>���Y�.� ��"�N*=�E=���<*���8�Ϸ-<'U����=Uz1��{�<]�O<:Da<Y�T9��]=j<N8l�A�ûT�o<��E=��<�E��T} =)'=l*�<`�z;��@��l��?��<�=�T;=��;�V=���<�@=�h�9#1����� �<��U�=�r=E㨼qy����B��.=I^\��	��h�#1{�K�=��S���'=L�=��_������0���v<RJ�>�j=�W�<;)�;"�:.�	�H�n�v�z=;$	���5�vI��/ɿ<��<�������[<=�~9���<�#=�SQ;�(��B���]k�<!(��&��$�iᚸ�'������A=�ڬ;��ջ�n=���;�G���k=g�M�ϽP�qL>=&v���<m�*=�=��R����G��\l=��,=06����;���i��<�ml���ߝJ=��-�h�u9nv�<@�|��w"��q(=�z�����<��=��l=�4ݼ (Z����M�=Ϙ��D=1���޼�$P��Au;}i��}D�<o
=G�k�gE��#*�<�ѵ<�zx<��=:��=�Y�<�]=!=n<��	�|�<Q�<��;M��:�g�<�l�<{t/=�(����޻Y��?������<��z=��B=��X�������<�y�<�&=��A5��=�Ǽ�#.<2a0=�^N=��BL�<Yyi=�?=��C��SF=�i��L�9���;=��;D��te�<���U��@�A� �]k�nw�<������ ���P�B[���O=��q�g�S�������h��}��ϼ~�=��=<�� <����Bռ�R���=~jm=ﻗ=I4=~1]���Լ���=T�=�f�<��W������;��4��h�=� ��8}<�&�<DJP��%"���;����y����;���;8%
=�,��Y=PF7=
@G���=h�U=��2�q��<S�̼-0d��	�/�X=ehB�����ߨ<\��/͒<��^=Wt�<�B9����i�]��)5�gḼ��<BO�:E5<��+��=��g=�x[=,�Q��=I�n;A�,�� ļ�]=��o�3��<�<�a�:	#���W�s�����=<\���=�	0��_�� I�;3�`=�"�%*H��u5� �o�º*<uRG����]�<��i<�)�%�]=V=�&�a軲��k�v�#L<��$�\6����:��Z=��<M����N=�I�<��n;&�G=?�V=��R=�뼼�A�=�`�<����zj?=4�@�������nk�<r�(=�0=T�@�¥�;öS����;�Q�����g�)=��%�ۿf<�Yu;s�/��o���N<I��U�<�][����<L"�;L��چ�<gT<��L=�a=���;�P2��+ =ڷ}���!=�A6�0���=H�G���g^�ؕ3=J�=� �G~/�\�7���G�J�2�z�H=�8R��+�
r�<�C=<�|ͼ�7�;��z=,�.=Rnh�J�1<�����<K_&=i��~��9x=�``�<��F;<��;��ۼٟ<��=T4	�>�1=�NU=�q<	�<}=�*���q<���<���i#���Z=9ͺZ]<{(9�y��؉M��h�<3Kb��6q<Y=�� ��%ļ	b��+�<V2��{���LŻ��+�:��?�k<�{#=l��U��=��9[�<��A� �ߒ=�j�<U�<����޳�?b=����(� 8p�W��>�<�pü:�<-r�<qWG�s�[��@�<�L�^�=��ͼ��/8a��<�f=��:h�;1�n�G8�<_3�=�9�o�B=���FK�FA�� =�X\<f�A�2xƼ�b��v>=
��<�1�	4M�V� =`�#���<Gԥ< �m�<s^$�%�`�)�g�|���=���;$�<�2�<�OѼo���b���
L���ջ}�;f��� �^�|�V����S=Qm=���Caؼ�����^�~{=�w�d�<�"�ϷD�}H=��;�z��;�;2D� ��<ϓ������Ʒ��mμ�F[��D�=����=�90=�)=Ov�d�;kr>���V==Z�G*t�I�C<�J�|��w�=�����\=ۊ�;�`+=?d=�\�y�
��A���v���:���<��=�l:�V�<ג�G�D=n�S�u3;u9����<�����ʼ���;_|= =5=������;0&=n������]��<��ʼ�����<0�&��t������;��=�/=7��;Y��:��==���������]��8��9�j�,+ռ?���=M7=���<�;0���¤)=d�T=Ֆ;<��<�7l��|Z=�����/=���<��J���-�w�0<{�n=O'^�g�<� =�Cy<<��<"=�㜻�ՙ;��\��m#<Ui�=�;�Bo=�'=�HL�I��<P���T�;cC�<8�w�C��J�E\�<��M=�/=�`�<��=:R�;�_=��<���<y3=�i�;{=�_=l����<��j<U��<
�V��#Z�C�<�^=N=C�<��h�{�=>(�܈"=Ly���B���QS�x��)�<2��<�K=/�<7�=n�����m�أܼ5�=k���G��h�<�`t��2�<D��G&�։��_<^���μz"V=9`�5�<�Ҡ<��[�X��vlڼ���4�x���$��.<�x�z1�+���0ɼ���|��<e*�<��<��;���8�X��<>���fp�r/�;V`�<Q@<l�:NN<SѼF��;'���Gt�"�F��n=w"?=�/��{V<�B<ϔ!=��{��z<�A;�c�E=�]6=H2�6U#�ܪ%=R!�<|o�<w�JV�=�
D��SG�g��U�-��xr<(}<
�PCQ<j]K��	=����*=@V�<S�uo��=�����!&=��=�5i��I=��a�ǼU-��a��������<�����ÊI<�jV<С�<�bݼyQD=�<��R^���$<��<�0�Z\���0�y����t��k��VO=+� =��Ǽr��>?�o�ּ��=�Z��*<=6y[�I�)�]����"�,�ۼ =�� s��Y=:I<�E=���<p�=��"��$!=)��<ި��L=�p=��3=�: ��V?�y\@���w=Mƫ<�Ə<x�=P��<"M,��G'���F=,�.��M<�����&��"W=p"̼��U����<�o=��==���'�;�c��1y=�G�2������4᳻w���S�˻]<��Z<[-;�(��+�;�� =����#m<2W��=�A=Q�����%�}�[<M�
=��b=�/�њ��"����<�{B��mؼ�T<h�I����<�Ԗ��z�<�f%�n�z�t\��N<�V<�#=��])�g�=15=)w�<0I(�R�5��(�N?<��<qj&=]%=�����L=���<�
N������M/=;�o=��0= K=p</��>=6�;n��<<$��d3<\�=EN�<�m��<=j�u�*���^˼j?���u'=����#��<�F�E�d=~�;=9�W��+:�ɤ��f��:ǘ"�q&=��7=�b2��H&��O�<�&ֻ^5U<z�S�z�2�l��<��]=�P�F�3��-���5��OƼz�X�p/=/��;��C��M<��-=�"<,=�3=�0T=�H
=�j=(&�<��<��"<���<E�x=j_A;mo���2�9X�-L<ڢU���ۼ���<s'==�-�<�J=LR��[<= �=�o=^,�]hM<���<͉����+�W�<�j�<ǲ-�A��<��<�8��_9Q<�]�<���u��;N�;��ٳ���H�=���/;�;50H=}H'=����e� =+_(��
�<��@��񰻌�N���C�ؐ<4��b�<5=��T�=״[���i�ּ�산���D���H���'�j�F�}��Gn;�G�<> �ք� ��<��o<�J�Ӈw<��6=՘� G��i���<�)��F�<��ټ���Q��<�=ϼ:��<ZR&=�Qr��}���:A�=��e�J�I�zpg���� =���<��
=�ii�┕�:{��(�X�_8�~�ݼs&Q�&ŗ�CA��-a�7����[	Ļ��;��8�0q;��3=d�G=.����XD��i=����S�c@�S'%� "B=��=��)u��������m=]�W���a-��M�<��-�Yy=ZI?=�i/=V�<	$C=�"��K�?=j=Qۦ�&k=�ad�<�y��7���%��"<��="�;tӼ���;g�F�`J����h��'g=z����E='�<��=�=���	=�Vb=eC�2�=)�G����2��<��=��8�.�<�%�--���N�w#���~`=��2=��'=1��$^_='r��b��#�;_�<��T=6�A�Z���j[E;�V��FÒ���6���<pM���P��;\�)�9<+Ҫ;٬�;"��;�l=�jV��S:��N��&Y�l!<8��c�=�A�#�;1g�<��h��i���D�ZC3=��-��L�A�1�Lq@�m%�<b����a=�ƃ�4��N%�<��<��ɼ8�|=J[	<}�< ����v�I=��L�"���Cg��}M�^�%�z��<tX���'=�ݙ��<-=zf=�ɼr�x=5��:��]=������=��u�����#ԉ=�d�N=�q�ӼK�	��/�=�;Qj<��<����jR��f,���B'='�+<�J=zQ1<�M�:=�&�6��Y��<�X�p����sn=���g�v-=�w<}=N�W=۾<8��<d�>�f[3=L�=�F�;hU�:�ߍ<��Q��|�<#���q�g:i��RQ<FY�<kW����I=��<	�h:��/�Yd�<�h=(�	<|�_=�D�<�k;<��<=�	�tR��ؠ��W=�D��o�<�X3��͘<+#=a�X���r��X=Mf�<�$���蒻\�/�8�ʼo2�;)Fi�%�=B�9�jH�<P�K=�9c�n�5=�-��2E�	��;�IY=����P�7�uT�8�d=��!=>��<�f���޼>�����=a�����;`�h�o <�&=���<�W6�Rۨ�o����-�'����l� '��E6����<���Mj)<�Գ�*[=�t=�H7�!h>=r>�������� �%=/�1=>�7<*�0;s�<�x<����V��q��c=M�,=�B���t3=�j�TI!�V&���;A�<d��<4�N��p*��l���6�r=�vZ=4�,=��<��0=�?���4=�A=Vb��=���<dl=<W=b�B=��B�8Q=={��<�����=�/���L=+#�B�<��<������X�F�@:[p�:��Ἲ���
WW�'�ͼ��9=�<�>b�h�<�Ǹ<�!=�-�$��X��*=�7=Đ-�<N%=3
��/Q�;���<�K�<v�<��y= �O=����`c*�>���C꼮��:�G=il8<ZN=��/�Ĵ�:`�-�!�ļ�,�lW0�N�C=�Q<�#�!	���kA=Kv!=������U<���<.0�<��=j?��?�'<Zo��?μ8C�;_h+<Ⱥ���C<������!;�쐽+Y<<,��<.�8���S=v�L���D�����<[iS��+<�n��ݛ(�-�^=�'g=�h�:�;cA=�p=��ﺲ�)�QnS=.�:Oc����.�'�s�%;��E�������:�h�3�P=p_N���7��t�<q{��,={��ٗ�<�<�i=ߚ2�N��=�ߦ<���<�r@��?�<��(=IA�����]=EL�2�"=�<��	���=���;��~Y\����Qμ��)�u��<�A=��n����<ο��C.:=�`	<6{}��+=�V�x�=�"��Ǖ6���f�U�X�hi�o�E=Tp�f�0;{NT�Mz����?�{s�<c3Y��0��T}�<��<^��<���<ZQ�<���US�@"����=�P��h��<B�=���g^
=MN�)�a��5�<��ͻIB�ћ(<Iʅ=��l�<w=^��<��f=G^=�l�< $@<��һ���<w�8=�u�y$V���0���'�XZe��_=�]<�Fȼ�#��3=�Q=p},=��(=��;;=�J�-;��-!=�'��"-F=�'m��ż�T���;c����Q����KJ�1�����:��M��v=?ϫ<�m<�r�%�8�� =w�<x�=���<���<�w�����$�LL�<$��=uF=	����N�z�1��==���μȺ�=��h��UC�+R#=�<�a0V=*B��Y8=0��<��=:�=�|��O�<�_���H�<ۆ��T�<s���a�W���b�;^W�;x!E�+s�<�!�<�eX=��<ߣ���/=���_�����v����;���;%�_��O<{=u�I<��꼉�R���=��R=2%I=h8(��5�� �;���<�͝�����خ<@)��ߥ<P�\=oy"���ϻ�<{4�<�`=j^����?����<p�;5\��&��5̊���S=�\=»:���(;-�(=��<.�U��4��ki�i )����[
�;�i������Fl�<��%=�rK���|<_���m���I���0=(�E�.�#=*ܓ=�/��0߼�3���V;;�@=w��C-=E:=访�T�=�=̔=��z='��<�[�<�Dl;�^���q�h�<�����E�ɨF=�pL����%�d��SD��K�<?m���/=!ZX� mƼ�f�=�=��<A�=<轼<7e=
vS�5;N�	����$Y<f�t;i�i�rI��d1=VP����<�NL<��m=��<x�a��ٔ��5=��0=��<lQ��q�7=7�!�T�W�L�5=��a=�c�<��n=��<�)���$��k�=��.����R���^�����K=KZ]��;�;ӻ,=r�-;C]=b�<��NXa<�<��l����X�<^ �:co��Գ���/=�=_W<��˼"�F=ٱN�v���w=N�;�:��b=�N=­˻��<v��<&*"�X�<p3��Б�ᬤ��t�.�J<L�<�q=�s^��Z7���<�7�K�C��B=�=�B%�y,���$�O�ڻ�w =�j���W���.=�<�}��]iZ���5�/���3�(�=�F��)pP=���=���<W������]�Ҽ0�$�x��BZ=z���6=�W�<��<U"�<���<3�=�����'=R2��K��׼�_�<��#=�ꌽT[��S3��\� ���<��R�7@=9bG��A$=�<��<=L��͆}�>��<ĎM=�u;���k=���L=��y�M1���<=zĄ���Ƽ E;� �O<Ѽ*<I$=p�<>�"�rІ=��/���P=u��<�&�PJ��&�<өS=�G=�]H=��P�ԯ�;%<���<P����<�[}���N���G�+WL�N?<b�U�A�;Wt�5�m<.67��1�W=��D�*�;?$Y�:fl=� F=�dz�Q�;.
<C�� ��3F��YX=��D=��?�����	CO��^�<I�=b��<�|=�P<w-�򬧼��<�2���:=�-;<"�L���(�b	n;N�=ŋc<�'��H'���n�5kM=ʤ"=��E=��y�`@7=�p]=?�
=P�=?vݼ��1�J�E=|�'<z���b�<R�g=<솼�T�;|��6�r<ҕt<
�S<��z�<=z�3K��%�1�+��"�<ٵ���X�y}=˒M=�$=P��;hm���E��=��C?�<|A/���<�{I���<58=l�<4y={"ּ6�==����0������#h)��k|���,<z�=���<�k�<ν<Ԛ�����8c<VBm��ټ&������l�����=��o=7~�<џ�<�hm=*�u�!n�<���v����3=/����{�؋6;�o���������w�����!�B��D��1D8���<@�;��=���*�G�/=�N��	"	���<�컟�L=;��<1l����6<\���N�;�=,��'�<�wc<
��=_�=��k=� I�~��<��`�D=��D=QQ�����B�:e�f�"==<컼o�;לN�hi< ��+�)����<'�<#��g����8��z%=Ot�=38�<_4�<�<�>)��W�<�ڂ�.�L=�Ż��X=y�h�l��<���<��<�*0��g=͘)�6�%=�݁<G�~�P�#v=��%�i�9=��w�
���s.�v�!��K�1Br���<ËǼ~��<�>����<	�$1M�^p�<�w	�s�<?PK=O�.�n�����	=���"�$=*�;�OT�[_����<?Q�<m�=4A���=Q�+����<��=R���ʨ����<>�=x
�<T�=�w�F�:׭�<1[�;�#���B��4��1�=㾃�o�'=�N�<M7�#�={+�1P~���0<�`*=�t�������t=�e
=H��;�!L<4D�<�/�Rl�dd�c��2�:���4��#�8��ۻ��u<>=�y�B:�Wj<��k�P&e�%\�3�5�zh�<�KC<ˌ�G=��n;H;�����<�?�<�9=��<�Lo,�]����P�3�a<��;U����Gy��oƼ���������m������H%������=�w=gK=��`���2��Ǟ�t��;�{L���4�Xͬ��v�9r޼���:0V=�5<�8M���<Z�<z�6�B=�.;GU[=ED3=0=d�l�Ƽ�TкXZ¼�<�~J=x.=@�}=OG�� /���<&�a �<#��N�:=���<�=�:=�#=5>��ۼ�1�znK<�:��l����v2=��H���D�u��:k��<q0<�kɼ��=S@�<!-R�	�<�@ݼ�E=��}<�]_=q"H=��=J-��V=;�ܼՎ<	&$=���tr�!�I=�����:�x�~=�H<ը�	8���G�<6=�&�<9�D=O拼eS�����ؼW	�8t���	<�a=	�<�i����=H%K��b�ӵ���O=��D�2|2=�c=e=�G*=]O�r�!�K�:=�A�1����>�`�\=�_=U-&�e�����_<)e$��8!�8dQ��x;���<��h=Aa,=���`��<��=��A=I�"���μ%<���Bk��UR���^=�F����;����~��Wͼ����#t;6�м:���U<�%(�s��<tUt���H��=�=[�c}�=]Y���$��rĺ���<��= �<=��;�#��Y�'=/�ZN���	=��O='1���ˈM�j�=�������2�<)�5�r���3�;�P�0U�;B�9�y#o<�$<m�j�X�v<�N�<+�>�Oa�:A�"��4=���[;��<�����#=ӝ��)��;^="5��S]����<��<�=�`A=�?=m�k���6;K�e�Q^�����!�=w����t=�2���K=�{;=\'f=6-�=J5��LĻ��R=�_&=뀂=Ƭ�;� �<�	ļ ��<B:;m<c)�<Q����,0=�����ļG�'=k2C��Uf<J�ɼrlR�*�=��J���@��y�<|����IK=M�<�7<�z=�@�:jo�!�F=U={�w롼DD�<9�*�pT��>��=�+N<[i<I>q��Oɼ�� <�R��H�<�>��P��J=�e�<�Mͼ-�S<U�ݼE�Z��{�.uk;���y.G��e^<�nL��ɜ�f+�<ň����<*�޼"k�=�I�;�������r=�a���0x<�=�*<�\��n��'k���L=Iy8��{
�j�e=�8{=��6���F�q�=�R�Gϒ��޼�&�)��;�5S=����*��G.��ۗ��8Q�Uxd=!�=1��a��<�pG��'F�{��;��f<V�6=��
��{���&��n�;K7�<��ݻsߟ��H�b3X�;f<�B�R�<��=������c���<�-0�C]-�И��X=h��w�;�L����	=%�<*Yh=z=��4���%=��v��� =�	��;�2=���;�yC=��ܼ�z����"=R�<D䉼�n��1��2�I=��!����<v��<�!_�yM������%��	<�mL=�j�<��7=Aq=��<}o�<�pq��Ix�(��<�H�_=D4ȼ��g=��b���ܼ�'���<���<tS��m�=diP=/(R�8��<�y��˼b��� i8����:'.�;�6f=	�W��U��:༒�;\>_�ym�<���}�=���[�ݺ���<��t����<cO�<��f��C=�ض<��=솖<��<J<=�ѝ<��g�MuP����U�ټa�f��!ּ�`�ʉ���Z�<~�s�#���$�;/f=�0��B=vg���K��q�H�* ����&�,W8�g?T=%xZ= O0�MXU�%B"=�=�t=-� �)q:=�k�;�\<�;X=H:8��D*�u(���E4�E���ou�� ����:�=�����l�<:3o���g��b<�\0���B��y<=CY��~=ӨS�@�J<,R��a =��;�3�r=8�<L0��JR��H����2�z{<��a<����t��M�����<s���q �<W0�Q�n=�L��^<� ��\_;5���(��T=v�a=b=�Q=/�J����;IJ�<K�
���*�~۔���=�w=��Ӽ.$==�z�-NQ=|��t��͋�<�;�<�陼ٸx<"��<��|�-���v=��z�N��x==�~#=��:6,��_���©<�]�����;���;h��읺EzY� <&����<�W���5�j9�m�<�
�<`C���&�<�����U=���Q��v�"��<�/=�O����<dv�������˰<c�h�(6�D�	=�(�ޠ�=_\[���h=g�Ѽ���=���<��	H�S���N�<��I=�%2;�����;n�L=u(�=o{�:�»?.;�.߼��<��o;���x�<h�=<����<V<�<zV�&F�<��;����1����D=��ֺ_��>-=��S��;<.SA=J˺�<�[<mV�W����=t*���O=Q��D�%<�j9=zmɼ�1�<�'n<�g�<��:u_= �]=��<��U����<3�P�x�Y���#��c��51�b� �Q;�a�<���=v��3Z	<���<=iF;��|<���#�V����=gsS�� =-|9��0���7��Aː�`O�<�=Z�Y�[l���<]T=��ݺ^7�������h�;�s=�Q@����<Ж���ټ�ۥ;}��N+�A���G�<�[�%uV<��=<�;���f��}��e=�oD�?6=��=?QS�l=j
<�}<Ŗ���߼�k2=h׺;�?b<��	�d�g<��L=����R+���Y=�[=�Gl���=��0�
-M=s��;��<������#*�.�^���g=�P���<rC���=\��:�*�=�V���۵��P=��6��GP���F��aD=�1����<xμ�<�ٲ_�+N*�Rэ:֕W���=7�-=aN<�>:t+��R�����A���=)���Ef=s?���:�<p�Ӽ��`�-�^֘<�$����<2�<����P�?��	�<�5��T4<6�g=��K��<@�<ă��i�^�ԺϼI��<���;Š���n2<V$Y����w"=�0.���Ul�W�[=E�?����%!�:�.�R�=�U���1=�˅�7;=o=^�W�s��`3;�9�զ��<&=�O=�G=
�=K���Y�=+�m=�� �<��4���=�
=\�v;�zY=��~=I�V=�(c����Fn�ָ�<D`��ʯ<B'�<�p�:�%V<-D��+��� �КӼ������<�6�<�l<��������.�ɞ*�X�2��O=1���v"��G�y������@�C��W���k%�U�[�<��s�;���Wp=	r��M�G9&�i����@�<�E�T�>�α��_ͼ�6�:��#k���y��D&=��<DmI=�H;=O��;�>ʺ#[��E�+s�����<5�"��3��F^�4��<�$W;ǻ<E̼;��<��9&�R�4=���;�Y�;z��;=ʈ�* e<-&s�QgN�M�=��:�=�̼�^�<I�<���t�:<7E�<��w��ZJ<��=LR`<(q���U;��D=��=]�I���,��<S���$0���=�4�&lʼ�9)=^�<��=���?�<=k.���)=ٖ=�λ���+�;��S=Ϛ��`��;�<��0���
<�`X=��~w��k�=>#�S�� �\��=�S�:=W�a�yJ =��<=G�]ן<�SB=�5h=c{1=zRx�d0޼�"�9qռ�==��<�tO=��<"�u��6��A9���W�;�\]��;=0i[=I�%��,v<-�d:��X=��<=*�*<�<��:B�\��7޼x�<0��;0!�����z=�=�T����<�n��^W=�w{�� S��0�����"A�1�׼0<��;�qK<mͻL�<�H^�+"�<ˤs�����g�
�=w�����F<�<V=Kf=_�$�1c=R�8���<�8�<��q�d�8<_�u����<��=V.+�F���w��v���g2�m\w�4a���gM��L��]b=P%D==�&=5:n=)�-= ��.~="�/�Z�G=�~��l�[	�i��<%f�����p��h�<�.qX�,i߻󨠼w<�,���3=�}<���3"=�5o=l֏�T�[n=��B�8�u��' =���-�W;S+�H*.�K�Z=��7=qq�<�:=��S=�m�X���?=)=]����nȺIY�:5���;��<F���t��);�H�0,���`I=��<2f�%J=Ćx�eF=?����U=��<J�2=U���_�<s"=69f���#�7<qn=�*��a+��g%=�� �<L<<%3�<_�N;�ἃy�<�;�<5�<����p<n���/��5Y�=�G�=���{C=��=d�&�%y��)��Tc�<:�i=Զ"=���<|�+=�F�<��=!�)�Nd�<�Hk�0�6��S��M=��Q��Ha=0�I��"P=:�f=�0F=U�G=�R=R<�=��l��<�+<��;�B��.Bs=���<<-=W=�'�h��pN��(���V��by<��]�w��^��!��<��;?<���� =��K����q<�՜��'<
g$�|�^�k�E=7��.��<��z=�A=Y#Q=��=1��e69�U+d<�һ�-��s޼I��<�)1��=p��m�<HG��9�!��]��f#�Bz~���;�^=XRG�UI}=a�-<�i�;`*=��=��<DvG�089���R��=;Q�;6��Ý<��0�~���
�`��<?��;�y=�{9�N-=�z�A2=u���<�n'��"=b��<O9=�ς�S�)@=y��]��XeK=�E=Z�׻�E0�M�=�G����C;�����=@����<+���yA=:<�dƻ�y;9�<ӷ��xf=+�=�Ϋ<��=bk���<Pv_�P��@ <���<�=,Ŋ<B�C���
=0,���c��8���W=ܠ�V��;��i=A~=}��"S��H���p<���<��=��_i=�>=D11=���=A=�;�"�;r���I8�yʺ<M
=S7��m=$W;=��!=_͐;�!=��T��s�D<z\���L<�?�&S=_?5����<�t=���<���<OHҼ�3=��=��]<Gu,���Q<�fG=��=v��}��<t�<�=e�=��=@'/=�&���_�;�{�yj=:�f;�7?=B=��'m���=��Y������GD=�r���T�C�+<�N�H�U=>����z�N	=��>=|^�<ư=r@�)�<ϒܺvg2�%�H=X��<(ļ<2�<�����2�8�Z=��=g��<���)�\vT��}<mo��R2=m��~�f�Q;/=�4)�V%q�產�4��u��<��G<�R}9T�;���<|Wz=�o�<7�l��� �>�U=XI㼔Ì:f@u���R���TL\<q�5��۷<ѡZ<�G�<�r=c �e�/�y;��`�� *�u%�<�y��jS<��<�M=7�V�u�A=���;:'�j��<zR�>=�R,=l-3;�żiI�<xB`=���ɸ'=��C�e�*=Y�:=��=A�T�S@b�YѼ��g��+�wpa<�N�~�>�����Y=�&B��u�7*����4����<�SF�ZF<�{==�z<��=.'<Ji=N�<�f6=�;���=�Ic���=��D��ݼ&Tg;~�(�]�N�}����y=w<=t1v=*2����6�=��<ab~�Fܣ�p��&���ɚ;�AA<Uk�<��<K�#�����=�P�����اA=ca�d�'=;`f<�;�<�Cü+%��*0=��3<�_A=���;Jyܼc|�(�N=q;0=�]��k�=Ӭ=p/=�(='J��˴/=-A��z<�y��lG����G���Eü�3=\���l�`u���k=�'�t�m�xp������\�;s(=�I/��S=5�<�{��4f�:��:My3=	K[<�E�T�=XK�FM�<p�=l�T=��P=�
�<C܂=e�<a�<�Fd���<��L���\��IV=e�9=G�<=\��<S�+=���<�xP=n�L���<�f"����Z����	=������=��M�5D��2�.='���񇼸�Լ���<�3�ވ<����M'	= ��"yR;��b<ZЗ�"I��^=0w`��<���:�$�<sI�L�=����qE���<c���2��}�6;�]����:���V�F�^�=.����~?�@Qc�����A�\<������"=ƣD=�r�����\�<)�*�H�F=*`�<�Q�<غ�<Ϥ�<)�7=��1=��S<���<���\n <�o��b��"$<����kP�<�������!g=���$J������q�L�=�ؿ��%�<f�3=���=tE�<��:=�;<�Y�����.=�h���{��[�<��=t�G<��]=�N=�Q�<�������Y=�*.��\!�b�MN<�p=�o�<e��\�ټ=pC=�<�'Ҽ��Q=b�<�!==ֈ^���H;����#�[�7�k<Le�����g�S�h<�~��������j��M=͉,=b�v���<�U���S�|&;�%y���<��;n�@=x�=^T=��h�����<V��z�ԕC���8��'�YS�8�=�<���={/�;}�o�e�����P�%���όϼ��z��u=z�U��bb=���<):<��Q�t�m�F��1==Z¼-��R�d=�li���<7�H�6��p*���D=�b��U������5�<~:;<��ǻ5��ˤ	={ǿ�����Kh��V���<:l=W[b���F=Z�=�C=ӌ���:�T��v�?<�=��f����<���������7g�(�:b���i��~�<2-�<#!=����<t�O��<c�B��߆���<X�V=�	߼П*��:U=ϙ���3=)SV=��q��.!����<�f�@����l�_
:S_��I��>�9Wm�<��<m`7��M�1�~<j�,=匭<v�<Z��<LA;��<1�_<�G=&qe<��<�;��G��Y����<ӨZ�EwP�xt
=G*�9�B��=Z(ѻ�Ǽ?�;9�2=�9(=��v���r�B�-�'wܼl�;=o�,=�WU<�@={k�����ơp<Š0=T+N���t=
��OmU=I�U��[8��x�= ��<˹˼D� ;�s�<L���:c���B�Ѽ�i�X��:z�=�z=T�
=.2��<�r�B:�e��xn� � �&�-����<�,=Xl�6s?<��B�;��< n$���E=��<z��n�<��8�%���f�J=�Ѫ���s��<{)G<T|T�q�/�@0�ͅ��?"=�ڼ���z-z=2,$=U;_�j:�ᨼ^A��=��A:#S�ײ�<i>�<Ԁ�:>=O��<�;ѻ\<�GA��z�P��=��5=�u2<"R���:]=���<���"v]=�<:=�;+�08�<�i=_F�˿=��>�Gg��J�U�i�9�w�	=w�)�K���u�;|Wӻ��ռL�j��<�B=j���N<S	������i��O"<��9�\_d�gP��وN=Q���`;�Q)�$h�#�%=X^C�h���MH=ǋ�*��
뼟s��l�<��<^-��cB#=�B=�T<\�:��1=zu���\����+�z=9�T���!�Z;�<~=���<x�\�!��:&�2=O=��<z<�V+���	�)e����;��H���<a��6ȻJ='\	=�2�<Bv<g�6;�$}��-�A�伉=ә�;-�꼇�<�j�'8�� �<�}1=��ݼ�2�楂�ӄ2����;a"��;�:�C=��J�����7������K��<0v<V=$C���u��ݵ�:kM��N�<6j=���g��E���k�,���v=��o���f�U}�<|S�U|+=�j=D1=X�<6,=�=L5]=�0�<�Ɗ�h�G=��(=�ļ�D���=���;֦����S���K;�0��<0^�<�O�;]���=�|�<3�'E'�.+
�#���I��Pt;~��:�:��1<��F�D=���������pG����<��ܼ�ɶ���мD��oޮ<�鼖�x=��$���<.`�<��jC|�Q[R��q>�������8=��<���<q͹<���;�9�/�<�t�h�w��<���<Yin���;�=�똼x�V=m�ٺIE]��=�8<=����^O�B��<�k� ���0��;&>=fU��C!�1�%=�\-�P�=0ܼ�K��Z%;�ȋ���R����<~�=��1<�ZQ<�E��'W=���9|����|8=n�����;�4J��r�:�N=�%ڼ�=��=��Ƽ�{�;v��<N��<XT��69�a�+Y�<x��|ӭ;1E�<��m�2=h�5<�	'� ������<�'���ܼԒ3=-Ҽ��<�#����7վ���#=��<�I�_��;�|=Ti[<Pƶ<S����S��\¼@r����<7i=��v�U�ۼ)z���?���ϼr-=�ë<˗�[C=�<W2�<����q�;�*=ΤS�e0�������q����R�(�nZH=�=�Y=��>��7=$��<���ܶ�<�BD;A��<x��c}޹>1=��,=�<��E�<\j�sW ��_��5��*ռ�3����=1�+��u5���<7�n�C�A����<M?<(��<U���"=�2L<s�ϼ�=s�"=厎�¶�cg�;el�l%g<W���%X��o
<%^պ�g=����뛆;���'��cJ=T�;ՙ#��,g=�E�;�q ;\�>=�R�<Z	�J�i=���<#%d����<��໾�T=��<��)=��.=U5���ٻ}bs�B{�;*UX�dBj�=�<s�=,	p��Y����f;]��=W3O=�3=�z1�T#��~������.�f=�(�|�8;"�=�0=�mμّ<=�<Y�=��ּ(3=�,=b?����,=^�<��������9�<(o`=l=�=�Q��� <���<
G�<*Q�<e拽�z?�0����<|�=����$l�<!@n��2?=5fW��,��%Ӽ�"<�4��$e=��=��2=X�=� =��	&�N�<b3u�gwU=������Ի�g<�a!=x�˼0�W=���<��̼*�!�Q�h=��μ��<� ���/�J�I����<�x���L���� %�	ڮ<���<�F��/�;O�;�5�<���:�ٻjL-��E�< c�����O���s���=�W���I�6�ں�}=��K���R���N<�O���D=(����z�lr=<�G����J=#�F=�=��;Af<��<�X����D=ca�I�<������wpe���&=��^=��^=��C=�!�y]F;tL�<�?X�9%:g9O;-����k=Z���F ,���$=}E��hUb�X+!=9��� R7��}={ؼ�W�ּ�Oۼ�(�7~[�d���i�<��ElE��y[<U8�<�qPc���=+�<T��K�=+�;uMK�/<=�̫�a�O=k�]<Ҧ>=���0��{��(�d�c滔6˼#O����X;�
=Fo<� �Y=��a=u��:9�%��żep��0��lK�;m���n����/�̰��,�9�mo�r�s�hQ=Jo^=�ļp�]=��j��bD=3�P=Z�=\[ =0[e���*������6�=�j7=$=3Y�<�8�B�$�9� �ݯ�:�g=�xS�d��<�켬���F�2=ǿ/���I�+駼��<����g������<�����|���is=d���C3��T�j�=��c;�r*�}F�<Ģ!=���9��X=6iP=�
H=	f���"?���d%=BZ��E�i9%�Y'$��{<���<�+S=�6)�M�*<C��;��=�����%�(�v�=΀ ���M����:�(�<����
=�yX=�8<��L�S&���`=@I�;� ݺ_�����N8��Ȏ<���<a=^쓻��<��<���:��Y<�g����=Om޼&6���#�\ <����$���O=+�V� ��<1n ��5G������7.�'-�.!=8AW�r<�<�L��`!=���,]���m&=�y�<S�Y=�
U=��w<��c��7;=!c�;l;�<.��<[�]�3����<�KM=�6%=�f��Y83�	��;
)�=j 7��_�<6�<�h�<4�(<��J�7b;��d<�Y���V=!0��e�mF��}����a<kq�<��"�$�e��T��Nռi�D=x�:����Ms=�2 =���t��:޽�=�x	�����ۼ��<��]�Q\��'�	��R�<\�E��Q=�W%���������Isp=����=\P⼐�<�>��:|�X=�o�;�p(=>D0=6$�Y�(=�2�<��.��������<�Y��H�A;��]=)==��j�<��< [<��(�C��L��<N`Z=ŀ�;Wn�9U=��:�=�޼�7��;�B=���<�]9��%z=��V�e[���'�	�l<_�<�)�:Kî�p���hb�H�m=]�<����!��OlJ����<1�;��V=oO=o���ZF�=�=~F����=��>��R<�`��V��<��<�d���<Q��<>e�� ����<U(�<�~h��V1=�n=o!I<�磼5m==`���<��+���A����<o���m=X��E���ش|��<(�ּM��9�;�<�b<q�<<-�=Қ�;���<�W;k1.�j�X������V��5"=o.�&�@���0���B��'�W9�9���;�V=��K;�eǼ�m�<�"�V6�$�)=��]=S�Q��鷼��D�E2*=�=d]���:=���
�����<��x<>�+<� =0rn��{-��v���	S<"&�8%C���$�(+��Դ�:w9��e�<W=�.�<��;��G�ߒͼ�͘��B=�Wu;�?�<�8@;�ڻo�>�{�;��=T�=��.;�A2��fE�=/�YvM<k��<�����<L��:O�(�!�
=m3E=+�F=��<%}м�ڥ;�09���I��{��ޞK=��_�D'"�Eۉ�&]=[�����"�<��Լ6�t�-6�<�3<o�=��O=������<=�ל�Hl$����<gkܼ|� �Fj=��<���;�I>9.?==k�<�W�ˣa<�����2n�>����
�/a���<;�����@O�=�ޣ�e���7�	=�h}��#��2�<k����d�E��F�=��<�ڋ-�qO��'6P���&����tL=qV�co>�,^�<� ���3������=�(=��$�r^h��hB=�q4=]'L�$�f<����:��p1���G5�ਟ�SR��c=<�v<X�7=v;�gt��}��� � ��Yɽ����?#�Rd#=�����Z�<�i`<�Y��Y��<v��:��?���%<�V0=�0�ag=�T;Dc6=��6C=����Q���%�9Pv��Mp=�0мE�μ�g(����<߻r<rZI��b!�'n/<�<1k�Qg�<��ļđl�[�R�z>��5�r=ON�<8.���.=�Y���0b=�z�;�C�<_t|<nK=Ŭ����)�oC��6R=3�=�Y�<i���cǼ����=F��<=vI�=��=<�r^��p�	��;��ļN=��7�	�4�k2�{��;�����;�p�v���z�3<e�s�kQ���D=v�<��D<[$s=���*X�I<��@M;B<
���<�O8=g�T��,=+�=&���ɶV�kVa<<�;{(#�~/:<���:bQƼq=�����Qּl��<�r<'��<<'|�r�uda<�>=�2������-��V�{<�38;o
�+-O< 닼������;�6k��R/�<���M]��&=?0Q�W�5=2O�<+j=�Fb���<�LH=�O�<�z����P<d>⼇��<��c�=�=���<�������K��;4<����!�9<�V� ��< l'���<.����<���<�[��5���Ӽ�r������q=���;�%�����qp�h�L<$��<r�/=��<-O�<��x<��	��=]�9�[�A�ix��H�U=��P�
M�����9�qD=��(=or+��)��颼fc+=Kp��G��U+<<�ּ|�<@;�'<GC���{�Mf�<̻��I=��N��8��tS=�ـ=��<2?2�/c�<xv&���9��;�H;+?ûm	�TԼ4[ռ L���==�Jx��F=�n�<ډN��V���4b= w�fD=�p<�e=?J=ܙA=�!H����<��=td<�7�<m@b��j,����<�8J=�9Ѽ/X@=�zx=�i=�4ɼ�x��n�s��< ()=��<���<""�L��O���R;"Ѽc�w�v{�<Z�����<���<��r��6����;-���Z�<S�Լ'|�<�1=�䆽͆�=VX���%�LGK����<�]����kZ��=p<KE鼦}=�:Ｕ�=� f=�3|=P�=����A'!<?l=@�ż���;XrE�b恽�}�<r��:��$�=��"=6l<0v���/�ʼ"��=���	��/=�+=����=N&�<���<�U���=$��<�Y����<��J��:F����<Q/�v1��F<uWf��5=0T�<2!=gh<?�<�=1'<�ݺ)k���=��[����мO��<]=j��;�>߼�W�=\��<�mR=�UB��M�	��;�\<n��<��2��2t<zzs<��2<(s漾<�: e�;���<�V= ���R���S�6��;ˣ=imżϼ�)G��R�<�x1=��߼^���o�+r,�%�Ѻ��l<\���H�y�����]�l=�=]�?=r�����0�Y~��y�=)��< T���4<�	��h�	��<"��<#�,���4�H>�<$9�j�<��u��<���<\G=V6�<��=K����<2����G=�0�;D5�yh����<lL�<�b�y�D���'�>i_<q�=��\=��<!D=����ر`<K�=�Ί���^f��wT=.=�=H�O|4=�ʼ�>�n��<~>!=	`=�J4�*=ȵ=:ځ<��]=b,�;�3Y=�d�k��;7;\\�k�Z�s=���I�<��a=��7�-Q���;�h=4p=H�<8U��8�<k�<}�=t<Q<u��P�����_;|�<l(#=����rC=ͫR�"J=�]�Ewżc^���S<��<��!L��^�;:��<��$�D���)�e9%�J�;��=��<�HY��ƺk���n���<"����a���S�Oռ_}+�In<,;��L�Q=�6=�M�|��xU=�a����t=�3=��:2�qE��������G��;��q��u=Qr��ܘ��nW���R=��+=����)����j&=�Rh��`r���L�<D�D=��<H�L<)9=�	=Lװ< �)��u=�C;�l:���ͼ�}z;7��ms�;_�@<J�L�Ǖ�<j�F=��a�/�����<�L=��E�
2�<�SB<�)=���~<A��f\5�	`��&=�W�<wC���j�;��_=���;h/g��7�E��
I;H@"��MD=%?�<y:=�>P�ȍ;�<j�"�<���K ��"�z�Z��k���;l�ݻ�Ӽ�J��=�-���>=q�$��h=���:��ٷʢS=��<�$��&:��j=P~=�\;���4=ˑ
=E[��w�y�<���G=Z�*=�w-=�9�|�
��zk�
�üb�n�iJ=l���$-��S��=�"<n5�<�͹���w�>��2=*	�<�PC�x��S��&'��i�;0Ȗ�9��<6|Z��*=!,�Qan�Uc���=o�:~�$=��.���='"��G=Wa���9y<$J=�=+�@���ݻ�	=7�="R�rQ���:��A�֨ļL:ڼ��?�`��
_�<ц�:<�:yi��Ǔ��w����<��@=�*b<�pq<�uJ=���<}�<l��8�x�u�F<)-������+=���Ƽ(�&=��$y�<{�\�k(=eD�b=QC�<h[o< �t��k���=�zA=�� �,;���;C�=k��<��������X�I,'������#�<3�'�� H<�`v<h4h�/x=�H���y��Z%=��X���6=��E� �=�@
��d/=�%�<�4]��Ӽo������J=����������L=�\v<I��;-��<u�<2�<2=�f���oh=k��<�<����y}=����*=�3H;��v��>�6��<����=A�E���)�T�u=��e=��I�
�=أi=�����1�����l����O;�*=���<K*S���<��μ=l�=n~m=)��<Yi鼎���Y�13��{<��2�ɟ2:��`�vR��rZ=�w =�2�<���<v��=Ƽ[Uz�vAɼ?G}�i���@�;��D=�e'=��?�5�
�-U�	u8;��9=s�(�ʒo;�@f=I넽�V���=�~ȼ+@G����<��E<�޼3@=a�V=JR���H:6R	<��B�%cN�Y�3=�c>���k=���l�E��~C��d���=��4<HO�0ɻ���%Ǝ��ή<�(��=�<���8Y&�`�<�R+�"P=��}<�+=�PB�+��`���P��i���`�o�;F��R�Y<�cȼ��?=�T��6���E��#e�}���WH�,z5=zR�;9⫼�4O=��F=c'=a p;�L=1?��y:�IcX<gϪ<����<�^�/=e���-�U��l��ː]=�@���=��F<��?=ٞ��y=�M =�����)7=���<}-e=>�<�=9k��w=��7=��[����ƻ8󪻏$[����<�̼A�����N��;u�j�@�<��j�<�K��˿<��'=�y���꼯`+=�����;�d�����;�H=�g�� (��ի;f~�<d����z�z��<�]�e�<�(1� �w<�(^=^�#��J=�=,I�;ur�v�=fR�<��F�'id<�&4;�	�`w�<� ��uɺ퍝�ֻ͗g���9=�����%�ᨢ�%W��2b=�%9��wz�S�5���0d2=&��=� `�Tt#=o���U; =<�=��=yU�\WK�����.��O(�:�<5bлvq=]�+=�yN��7����˼�\=C �����}�l=��3=�aN=;;�;�`�<&;�q�7�f)���=�3�����Gqf=���<X��<��=�Ԫ�ԝ��"!������l= �L=ȗ=��t�.*T=�������AY���:�<��aWq��n$�����b����:���;Զ�<Rp�;�^�>i=O�h<>n4�LKi��aѼ-\j<��<�'<�������!�<��=�i<��!=�/f�V�=��F=6��:k�=��?=Z󻓈=�����9�;�rN= Z"�k�'=HY�vF|<�TT=˓�Y��<ļ��A��ͥ��G>=�q���e=�l8��dc���=#E���A�<�u��� r����ؒ==��.�%#�<
c���rE=�=LP�6�==�L�̸�;������컎���C��g��	=}��<T=���<6�[�-��q�<��H�y`:��{<<ʂ���<��	�<�P<R=�_I=�_Ǽ�N�V��:~(,=�釼'c�;Bm��Q�/<�켸#�<�l޼�7=��<�?N�p��<��;0-;"U=�<���;2
�<��3���#=�u="w<�w����=#��z^�����<G7=J�V9����ъ�<4�
��=�
ϼ�$i��D6<ŏ���P=,R��_P��O����/��V=NQ�<�x.;��<���09=�z>=)%=�Z���ܺ/Nt��.=F���5�==s�_=ȁZ��=/"�<H^�����j)A=��;�K��3=j[v=�0X=I�i<:a=�+=��U�Q�==&1�<��<�[��0;�i�]��;��L=˼=.Z<�d���7=�V=�]O;L�4��۲�ө�<(�Q������8��6j�[.�<ؑ;̎�L<|~�:Y< =o�ؼ�N�;2P;��켣d��8�=���;����T��<�Yy<$��<J�y8[���ϼ\W�<�=�/`��o=ze�] =�^�J�$=\����л�7����缓%i=@I�<�U�z�=;�7�Z<�u	<�\��с��%i?=1�{�P�&=�(=�N���*=X�F=� <SD���&=$_=�"���G=�ݼ����P�,W��Q����)=dPS��z�;�܊��Io��'�ex3���<�=g�=P�T=/�;�=�V�<	��?����f'=7���Z��<}`�<.�W�,�=]�V=V�=
"Y��b�<��<ξ<ع%=$}�5h4�=�j)=�߄��w�I<��/=v��kٹ��J=�I=�
꼔T�����<&$G=[9<*�(7�5I=3\�����<�^�;,�=I�7���L1=aꀽ�[�z�ϼ�z�;&�-=z�}<Z�=R/l=�Y�<4��<j��}|�B�RY
=���.l����cؾ<B��.�<�<s=���x����ؼ1�)��A��8�H�{Py<�"!�;�#=k\h��,�;��N�ĭD��(�^Z:=V��81T��Y\���1��@���C���_:����5�<��a�P��<S��<�r<N)м��?��<�C��͵<7�<���<��6��$�ѻJ��<�zK=}@$����;�#�=+	<�"��j
��8Z��q<=�'��N�;w{��=�����<���<��/=o�T���R=񹐼��̻�VټxxB�0�=�Eܼ�l��V7=X��<v�3=��;��U~�<� �X3 ��w1��PƼۆ*�s)W=������<%�;%�#���,<�W!=l�� *�<K;�;��Q��Y;��,=��B�P��.Gܼ �E���\=��g=����}Lܼ��˻8l�<k�<=�S������u���}A <��.=�p(�e�~�^�T=��|<�M�<���,}<���<G�.��D=�Pɻ�P����(�ϗz�kv�<y��<�1�|A=���,�9=$yb<Ų(��Lj=ơ��ab=��&�����R����!�27����=Xk�<��=e(I<��s���<�+��G^=t�=��O<�����E=%gͼ����]=�~��r���S��-��2���v+���A���A=_v���3��d�<����h˻/��<�p�<D�5=@�0=E�r��펼U���\���w�p���(=��<-�= >����<{�<p8ͺ��z<�ݢ�JQ��݊U<d����^*;H�<�i	��(�%�ݼS��q)�r�޼��ֻ��5��d޼�O�<N�<*��$�,=s�Ҽ�XN�O	=j�=���<�R$��p���XI���=ia�X�X:�s�<m�=�=�G��<Щ<�ǹ� S=:�P��q<X��9�mG���XE�;��<��<ڕ����Y���X�S�<{��;��=�Z��"�=��I�w�q;��B�9����t8<l'�;�Y�t�=n�=�^<�6=#_�I6=I9���TG=�K�;�pE�yO��;3O=�K�<��F=-�<0i�<�t=�'Oλ��7�'�<V�O��O�<^��<r/���<�==QؼE�*=mc-��|7=��<����Լ��<��N;���<��<���;�<��;Ɋ�<�μ��<�f�� �\���=0�F�y:�<�w\:���<�6�;�p����<!X]=_����U��i�<#���a=�4�<�����y��Pn=������<t�D�9u���z%�.!����D=@�U�WM�;e]�<z��<{9�<��ú��4�=�`��Y� {�</��;�A<���Β="�4����<{�=Pg���\�фd=9E����Se㼑67=�[�W6�<Y���:`<���;���<X�=#Y<=�$p���\=�n���.�.��<D��<�Q=�f=:i(�,��<�A�택<^KԼ7*�<wXr=�#�|�n����<�!=�s���!F�6+=tW<�T�'=�m�Z!μ�I=,�E=t@���N�<-�<�综0�; ��<�8�1=A%�<[����+<�e�<��#�%�/�Z=�˻��K��x��2>�G���s�/X̼;dͼ?-d��l���,@���<�-�C`=�x)�wMD=M�c=EG)��U=>���P�<R��;��=�
;�0^�<l,�<�E�=�-#��Z=#�� �=��<Hp<����Ą%<o���JxB=S��<�A��iM�	��<���aѼ��5=`N�<��U=Z�d��=^N=+�<����&+��x����Y�T���ad=�Oȼ��e��}�<w�7���;�u�;�I�;L�޼Ŝ)<+�f���;`7�w�	�����9�<T1a���.�ɂ�<k*�`tj=}&h��G8�P^=�#�fa.�Sn=ۼ�9�C���d��e�<��=��=��9=���<N�7=̩�;ڬo=�63�a��<9��<�Z�Y�B<'��<@z=���:��:�Y�����KE��"�<�����	�Ԩ��1==�mW+�2���܀;s�=Ѭ��=n���Ӻ�ﾡ<c�==�l�<2<�<����Cw�=� =��<Α=�
�2��<�V�{���ɿ���T=�fJ��*�<n���7�R� �<���l�˼~�U�=e5�=<p��:Y*= 	=y��<՛�:�c=������<�^�dN��=h<���<�_7��4�6� ��(_=50e����)@=��<\� ��[���XR=\=�<��B�l�&�h���"�Ѽ�uF=�H��M�-=�]<��<(+Z=��"��=3#�~�H=P: =�v\���뼮fR=�Ke�I$=L��H���2S��̯<]���ji߼=𨼱�$�P�u=�!�;0@=W�ʼ>�<I�[��<:�
�<�M<$��<wO���C��G 3<��Q�u�A<�?#=G�����<�R6�oW����W&�c�=�����<��b<!�j��b�Y=�0��K�;<G�=��̻�O�j���O=�N��g=�@7�C�B<��`;y��<B�7���M�I��KIr=�DQ�K�}=_��<7B�;�����;r�Ż�fq�8x=hh�<�<S���e=B>=}��;�y���;9\�<�u�<�,=s(=:�/=�䜼(��¬<�Յ�uҦ<�1��<��
��鼨�R�*��B&�m�=*c�;��d=^2=��;1�;ƅ�<L�:=c��C =Y-R=z?="� ��)Z��<1�<���%`b=�;.�`b>=e�};�XS: �%=�F�;��=,����<ӊ�X�=XY��N�9<�P�W:��<��S�<��+��g=m��BU��v �T�o=E��3�ü;d���<���;��=�$=`��<V���Ŵ���^�[?8=���[=Wh�<���<�'����2=xk��H���(�<U���a=?;���U���	���3��uݼ�|(=��/=�&d=Y�������<�< =�F�<�Q��9�UO<�Y=�Y���]=Qq�<�k=�7U���J�����^.=�2#�T��RĒ�b� <��`��$6��bT���z�Fa�8�>;~Fj=}�K<�1=�ԉ<�ѓ�[jF=o��j?=�t[;���B��(��{�m�~�	��9;-�I=�B^=�>=F�鼱�ż��R=\��#T�<i�E����<	��|��<��{��5]���q=C�<�=r�.�|��<�K=4 �<�WE<� =c�/��u=e+�<��I<6l	��?=!��zl�<�{��xY���*��O��#$=�4,��󼹼=�''��S=�=�%�G9= k=�]X�&��q2?<�䌼!��ڀ�Y=M�=g��<� �<�7=�K^��P�g�K��R�<0�=�6�_+8=-:��̢;|���-:=O��e�I=��'�&���+���J��j==p�TԎ���D=�7n<�^]=�	��+=~�=��l{��Z�l�6=~�Q�+�=�y�;�Ջ<R����<���<N�<�b �?�.=�;=�.@=Q�y=�E^�� �X4��劯��f=!���E�"����-�=�<=]f��p<�x�<��\��׭;�F/=��<��м�4=�ɢ���,�#�H���.�y��<_�m=d�&�~"�<����$�����<��Z=X��J��7����;EN�<7���/1�<�v�<t1=)���`ۼ}2 ���<�~=�=��P�;���<p�S=���<��!��ab=�t9�$���(^�׍�=�9=��<��6=浒�Tk@���,<@~�<�h|=�A�=�%����/�)=߀=�:j=U�I=���M���":=(Ec=�=�:�=9_%�ȱ1=�N=���H��%=��i={d�<�GQ������=*��<"�Ȼ�����һ�N��ʴ��ꚻ�D�/ż/x2�C�.=�?=6E¼�s���=.D�<���<>�:d�T��x�<W�=Jf;d�=�c<o{=ό<�O%���:�pz<;�λ�*=I�q���p�J�I���!��� <�֜�6�޼J@e=[�*<�G�Ϡ�ҧ<G�o��8ּc�<XrG=3+'�5�W���Q��,������k�<ws^�e�׼)�=O�ໂ���aټ� <��t��<�c��Z�<5 �;�/S=�.�<��A=yL� 6����:��&��˂<8�.����9��<��:�x\=r1�<�L�<�=������`<��*=�yI=�A;=���Q� =kW��nbH=��X�o<]�޼s�!C��!�I=!��m�@=�X��<��<�m��`P<7<�m��3?�<]���ռz?=�60��{8�q<j\����8=��Y=Zg<iJ�;YS�|=f�@<;M��~P=K�ռk��=	C ��Y����=��<Kb;q�5���<s��<k<Sކ<����PUU;�����-ּ��=�h=�2L�{4��J�F<h08<�~0=g�7=��5<�c�!>=����G=ʯK�zB=��!�;]���Nڇ�M}:��l�X�L=B��;���w�l=�%��7��Oe5=�V��J }��S�]�a��.���=Av�"�<�/?=�z*��_= �m��Ҁ<�Ő<�ʋ�4�<=�f�<Y�<e5<�;?=��f��>��H=v���V =�K=u���4暻P�5��qǺKvX=�b�:ι(��v#��9��4Ѫ��	�=�j/�Uy�<Y���a�H�~F�9�3�1w�&q�<D!����(����<zL�YZ==X1H����@&=^���"�Mh�<�G�����;;��<���<IK�<(��V@�<\��<G�g;O. =��#=�4�<u`�<F)$=fBL<V9,�|���[f=�[;]7��K̼�XJ�ޠ"���F=�i ���=�#ԺMm�}v�OU�ǣd�h9=���K�
g�i=M;e�\:V�x;��a�
�����K�B�<�����������;8[=�z��|>@=�p�B��<iB��=v��:p�����;�)=���<m�=���=�kY=��h=�y�;�dr<w$�:�@F�Z"=u"=G�=�6��ڼ�R�<.l+=���旁�q�Z=?�,�l�Y2Q�p�_�J�߼�R�@$1=�׼���<}*A=��A=/�o�=�7���~�m�1<rfF�6l'=�~�;�\���@�.d=\�f=�`,=x��<�<_����=!�0=��=��+���b=��i;x�<����V<;8����˻ʠ2�9�,��AH;[S�<s��`�F�6�<�!ݼz5�<x�U���;=�I=���LU=���~�B�N��<n�ļq���9�<	�%����GƼx	8=��/= 1=����5=��=��j���?���$<x)���p�!E�<vAe�C@�߸E<�=|���6D=���<o���l�C�=�n=d�n=M!=�-���nD��+;��E;�q�[~�<�W�<__<L��<Gx&�j�==�����;Gw
<���t�=����[r�<�s}=����3D}��

=��Y=s�����<$=�<�T���e��p[��G���^�>V<=e-=>9�<�[9=���<��=`���L�<�3�<�.�;J����6=�Pܼt����e�l���n==g�<���:e�ͼ�c��,:�<;���Ֆ<�:=5^L=� =�Ҽ��=�!�<��¼Jֆ<�^�x4�<?E+=f���}_W=s�S�!�D�>=!��<q�)�`��z込�T1��.E;�C=9><�'=���:�=~<�/=��'=R�<96=�KX<��x�Xv��缲����W��!M/=d��<�aj���)=Z�D=�#�ZHK��-=c	F=:�]<�/N��n�:9�H���6=�������F�Y�a=;�9��iW=Ys>=7���m!=Zo����<��-���R;�J=J��<�-�<��ǻ<c���$�<r�L�ME�;K����9���̼��=�Vg��6P��n15����B: �>�>���w�#<=��;��l<YKb��WK=�`Q�%�?�i����������\�<��V�¼���=��}��<�q=�1�=b�<T�L�E�==X��E�=v�e��#�������ޟ�<7�=U$�;��v<o������<'��<gL=`jI�M2��P�<�ɗ=�k�,�=o��7W���o�o����&�#>?��s	��$=�(v�jz$=��n�$`J=�0U�˼�<�>=�<C�#=�|߼��6��b>=�c�� �!=O�$=��ʻ�o=l�D��!/�oo0�U⬽���<}�=M��<�� ���;5"
<������}�ޞ =7�!��<�� =1���fZ|=�VG�l�<�}�s�(=0=q��<���e��:�p9�L1�<p8=z��;��$��R�]	k�&2=sƗ�����R滝]I��ۼ��<XV=>f=�����ɶ��8�I'=�y��7AJ=Y�������#Sl<��d=�n�H����<^��<�IU=�;}��<CZ�ºz�m�:?}�<?��<6h=w�E<�z��0�9�_�=��1ۼ#�	.R=~S=Z��<u�:r�<��v=u� �YwԼ�?=%+�<�׼�A�<�v�J�����;Q�)<u)%:�2���C;��:��N�\c<(�I<��(=+5�=�ü�R��)�/����M<�B2��45= Q����=�o�<�+�=�ӊ;KY�<��$��+f�3^W��$<�7=̍��c1���Q<���;����s�=t9H�A��^^�N<�<���<��7���<�S>��h=���<��O=V���e=��ͼ=/�[<�N�<�=�==�\=����H�Y��@�P��>hH�X)���Y�<}��<���<���`����*�}�м�ѼP�=��=K��>m0�����K�|j��
ƺ,t����<�{y�f{�<��`��7��m�<�1�<6�� !=�Bl=�F_�?�=���<�<�d�;��<��5='/���NK�JzI=�݄��Kh<�Ey�QC.=�����=5�7�<3�4=�ԥ����IWἜk�<������:��:=lq:=C3��\e=����~��<˚B=b�Ǽ�s�<z�uE�<�b�<��*��ⅼo>�<��H=�J�:4Y���=O�+=���7����";�x��X%���#;E�����<=�_=���d���\#���Zy��%I��dW��<�o[ü����g㋼�>=��N=B�i�]�/=��s<�r =�ka={���ǥ<E�J=xq=g��-~i��W=s�<o3�;�_���/=>�Ż�����~�ּ���v�<����><�Z[=�h�;��=T��<LS���<ӯ<��Y���;��;���ç_��v�(cv<��"���\6=��<���;��O=�Oļ��A��#�8�=�*���\=W{y��|��Ղ;?4�;���/p="&�<�-�<�@��ԑw���F<��4< J�Elv����<F<N�j=�=�����<r�ӻ^�<�E�<��)�$l�����~,W=	=�!'�H��i����d=�9�Je��P0<~m-<͟�;�CY=�� ���==���!�޼[tJ�L}P=U:H��\0�+�P���8�T ���~=}�������*t<����lV��{9D�50���[=n��<���<���ټxD��ļ�L����AQ���4G= �+��>p��O< dM�:���v+���<��]�^I<�R�<nN0�H%u<x!B<���<�2�;��V=]������<�&���<�z�2^�d�<���-����<?�<4)�<�=�w{=�V3�V�껔�h<�v�-�����=OLR�8R���W=�}<��b�&�0=���;.�<kf=$� �$(<���A�v=���<����Q�3=�Z]��-=
[��� ��G�<\�g=ҧ<��Ѽu�<�P<�m}=�B��;eF�*��<�֐��r���<M��<��ȼ�����J=DbW��6�y����}��"=�g�<�+ػxn<�1f	��q�<�@�K�K=�=L&���o�9=���<
AJ��u<��];�D:"�:=�[�u|h���/=O���Ơ<���P�*о<��g:"�:=tQ�=��<c����=R�;���<߀��	?�k=�1"=�Z�que=�����N���7�EZ�D�\���=sU=7x=^d���|<�����<�t�=�&1���g=�g�;�?j<LcY=M=��dh^��=ήI�^���@ˬ��E�@ր�+p(��L<#C}�2�&���<J����%�=�,���<�u��f��;���=tS�t����<�z��ߦ<x�/<�{=a|t;�������M��*I�ܩJ=��=%�=��A�6/,���L�� �<�X4=��	Z!=�n�<G'F�0︼W=W=���H�&���e=��=mG��q፽ZC6�U�K��x`�J%�����k�=�d\��Ŧ<�Jd���
=���D=��R�F¹��C�<C��&'<��<��<X�<	-�}�)����xX�� <
=���˝�</�1�׹;o�<�ht<x�>���U��=v<m�����<���<����_�3=% �<֋2=y�K�
�?�HU�& ��n�<H�2=�=�<��(=�JQ�hO�<:�`=���Yy��z�<v�L=GB<����<r�,=�G�C�.=�=���|�����<[���\�E=[�X=�*��f�>=���;��?��gq�'����,<=.ۼ*�.��u*��mB���g=b�|�<����w=e=H�)=ѐt=2K<�=��)�`y�;���S?��w��[N<�"}��]�<�I��3�=�)�<���<��<cl�<�g%=��)��u<̛@=Wj"=�K=��w���;���<�6k�Y�M=G�<�|ʳ�n�_�_H�D~-=��<���30�9�+��-�یL���;=� ���8��6y<Qd�<�R�;���:��;Y��	 �;�<Vc=��Ǽ�>[�!=���S=���<�/���2=w�H��!���d��(pY�M�e=m5<���<�F\��8(����7�h=A��#*=z�<��ć� Ǻ�R8=�N=�2.��''�ܳ����$�b��=P�n��^=�}�<��7=ޱ�~�T;�O<;k�;�	:��d=�x�D�=D�!�]�<}�S�B<y$f<+=7=>�4����] ={R=P�;�K��;���tB#�eh[=�k=F?������伭Θ�+HW=�E�<;�q=�W�+�p=[�$�!�=m3��뇽�p�<T����+<jH��9�=���؝(=q]��� =�
K���K<x��<�+{=6ü��o�׍���?<�ȥ�7O�:1��;4tn���=�$=/ ��gQ����<4J=�醼�=��9����<1M�<ؽ�<bO�b����T�!=�<�D4<3��z�`=.��
�C�@�<U���_��b=#�l���ͼM�C=b�;B�J=�@��AH<V�H�|��a�� 1��\=z�B=��<B;Iؼ
�<�0��`S=@R�a��=\=�>=߼Om2=O�6< ~L=iN���=Ę�;v <"��<��ʼ����a��}\=)n�<9c=!:+���C�̋<=�l;W=E�"=*����N���0� �;li=��/�WhF�|�1<�Nļ��b��� =ʯT=��;<��<���<@C�<�oj��IK:D��<�	=�*��-ռC�<|0���{5<=�	=�q߼t �"??=AM/�E�F=�t�=�4;�c�=�6=��R�(iN<��<t�,�$,�<����>,+<t+F=��p;z�"<���<��d=k8=�\�����<�{-�r@i��֨<���<}*I�|k�<�e��f��j#�<�<,8�zF;�
[=����l�<��o<׵�<�s���U�����
= ��f强RA=&���=�I�<�:��]S�<��j=L��<��~�$p~��Fd<ܞV=	�7�@<%P\=1.=��7=~���sP�$��<���b1=J_��MJ�<O�=�>~<1v/=Svk;�<�g=cIؼ��?<��"��T�<Xt��`¯=ǎ����V��-<�9=h^���������f�D=�v�wU=Q�~�����能v:���<�Y�<;o���&�ѢӼ�'��8=݋j���<^�!� +Ȼ�Y�<)\;H�=���� .=������<��<̿��ʡ!=���<��<�<���<�+3��%q����;�WM��꠻9?�<{r��Ǽ�&N�4 )���<�⇽M�<H=�B�@|*=
[><��O�gi[�N��&����k��D7��Z�r<{�==B7���=N�ɼ��<5�Kx=B����	缕�����$�_m<�r5=��O��=�A=��=	���;��<�=���8=�\�m[b���<������t0e<C���G�Q��ټz\��7�P;-k��$�L=��r;*^9��<
 ��(=|����u<nL���
P�e��"�`=7=1me�J���K�=���}_��/��ؐ�<g�r=o᛼�Q=��d�}10=�U�<�a=��Ż�����M<�g�<_=��<X�.=�u5=�:���OP=x7�9�L=^3�;����u���/=�_�<�;2�e�/�=��;c=_W��W��CV<@�y�e��q�ut�<���� �ܼ��<Wi�;�+�<n�<�LT���;}�<~�F�w<�
�<7�8�4
��s=/�<��d��>+���)���\=��:=�Y=p"I=֮���ȼu����OP=φ<	Z�<�M<2�Ǽ"%t�I�n�I�,�@���Q�b���<�\=�P��]2�<�wm��/��VF=��/W=�t�����1=X߻��;�7 G<wJY=��R;V�=��=��0=�o~���e��Q=<V<"Ys�uP�<�x�<�:=���e�7=_&���=��<�=.<��^=�ջ��8�S%�<��=e»�c�b�����4��?�;�UE�M�˼Mp?��Hh<�Y=�z�;?6=�Լ��\=�؃=��<�uo=-g2��yO=���l@���j=��<�x��7�U=DGL=��<�41������=��<ȎO�Eͪ:�/
�ׁ<1�B��+�/� ���E���S
�<7?=�w�<HA�[bJ=�c��)�m�A��?4=�OP<E�!=@��s]��Ӄ�{��0=��<�$�;�9��=��D=�|��oN=HA��
O�<�I=���;�0B�� d��ނ�wЀ=V��զ3=ɰy<�����w=Š=�v�<�?=<F@<�œ�<�<T�:�Ft��s��t�I�=��}���r<�>������<}�<�
=s�@��V<�
�d&��>#��Y����B=�����V��<�?��m3����<�A�R�<c�{<9��;r��=���<�˼�Ix<�U�9u�v�DI��(�Ԃ����<�u=PC����<*�2=���<�>c=V�<�Ir������|�<��S=�9�<��5<�E7�w�=�]>=z<��=�;P�5��=2;������k=L!���ر�Iɀ�����Z�5��i����g<P�<�A�;r'�w\:�<�<�=���Zg;t�=R�<��<=I�<T�?0�<��<�g���J=����V����˼M�=<�B�N�м��(�D�;MG�<�B=���r���.��CJ=�H#=P�*���:=�"��@=���@=
�
=�^�<�j<yX,=��Ѽ�[=���C���7��S O��2,�>l<�������<!n =���� �����b=�F�	�7��M�Ug�w�e=TA�ĕQ�}��<�H�<����e����9,��� ���	}=RS=�'�	}��8�<�l�<��q��</�=�^!�+�<�۳:d��<>�U=�E!<X/�<Lv<��\=!(�;�˼�y��{}���-=1; =�5�ϧ=��<:����8����;���<��F�t�	=#d/�7��<�/B��m �<͕�= �� �,�&=d�&��W<B4�;� ڻ1�׼����7=,�>=�w�<=� =�򵼌����*z=��i=��h���=
Qt<�y����<�c<&��<"̈́�D��<+D=�;= /L=.X��}j;#¨<���=�:=�q:=�����j@O���<<�v= jo�'���"X"<�O�����<8:���=$��<�hk=&L��;*P;\�G<c�<��m����;p��<^�)�b��;�g���A�������E���<p��<�o��7=ʢ�<W��:��"�5�2=s�C=��׼p�.��WJ�:¼��V=c�d<�?�C=.�7��i�=&�=�}�[=��*�@�elD�ǖ���r��l��u<�p�<��y��T�N�<R��AE<ժ�<;��{����
==j�$=����=&@<Z`���^7����"�ռ�Z���@;�#��n�<=d�*/�<Z����!X;\���*�;d�T<jޑ=#�B�����9�c�:���=����F��Z_�&��<;�!��O\��:m�K�<%iH�M#�wq��I@�P�=+�Q2x=�a]�2h����=@R��<�#9=��=.
b=t�=�&J�r�-�Ao,=��=���z�<H�\=��<�;(�X ��M=�.=]/=��;�G�<�sȼBTI�Z��Ѩb=#2�J��e8����)�;�kW=`�e�ƫ�<�Q��k�r<#]� ��"��^=QΧ���=�W�&F<o8�<���:B�f�I���#v�2G����<�DC=��j�ܾs�5�d����䄽�ч=�Uu�EW=�.=�&a=�7=`p�<�A=Q	��S>=��X;���<
)��Տ;̊l<��һ ���<=�+�<��(��:μG���<"����/�,��s<�����=�c<���<�r����j�*=�c6�vi=l�S=�<炞<�R)�ۄ�<���`=7J<qH�<���;�(��q��1s=/�k���=�6��������;l��M@�&�<_�H=��J�LO�;S�%<�	\����<\�%=P�!��=��<�8!<><4=/NԼaa�:Bqe��
::^	��g�<�4=M�C;����?/=�k8=�o=�l�<g�$=���9�>=�p+���I��=-T=en<=W)�<c���L����;�z¼�g<t�'�,t|=0��5��; �=��Z=���'��<ᛒ�y =����:6F��	������<<��-=�
��f=��V<my��G���,������/��<%:���S<�S=+�R<�ԕ<�8�<'�R��!;��(=w򳼺�D=;5�j!=�=�9ƣ���H��y�V�]�y�:��=�j����5<��r<})�&��+L�֯�:��⼾�N<��5<���;v�;��F��\�<vN��N��/<��;L�<C?�B��Z>q=��<:��"K�;���<�C�<m^$���$=k��;S<"�r=6X������=�V�(6X���}�T��:5���-=FϠ<�3=�,���B<v�%й�4����-=�:�<���<JN��������<�2=c��ע�<�?�=��6=S
�;��6= GH�3X�<z:
�	,���-�Į$=e��=:V�G<$�.=�b�I�+;Z&�;�
����;=�����u=�=o�R=|6�𸍼��<���<f�;�"��Q�n=Kͣ;�O�<�<g|e=�=�<d[��9��4�<V�{���-=zn��<=!_�<J�M=�;:=.�6=gH=#W3=[�]�1~`�d��<�X=��5=�7��L=*`�<��$���A��/<���	?[=�<�<��h�<j,�qt'�7	���<�ԕ;3D�;tY������^#��3:�-4�c�Y�,y��cD<T:<����4$<�0��p�C�5�{�C�k=�K���m���&h=Ƿ<\��+DɼnA=���P�)<6�<���;$��<�Z���e�<F>=#��=�����<s�=c�A�4=�}���G(=A�=�	�E�޹�l<#��<3�r�у�<b\�:��Cb�<�n���qɻ�x���ӻ\�S=ZW���U�<����Q��R�Ĝ�<g��;Xk��<i=3<�D�<G?���I��| =��c;H�=���;)Ꞽ�$�����kp��Y�=�����û�a������4��<�4�<���t�Y=��!��\]�>Y=A }�GP;���K�3�ɠ�<�@&=:�]<�{��^�<Sc.=�VF��9 <2;_����[��<ְ����E�:��{An�漥t�<1
�����<6�S<��<�m;�t�<תM���'��D$�D7�=�B= JB��������P"S�D�<�`*���<� �����#�Ѓ�<f��<8�#< �b=�ʼH�z<�-	�Զ�;+R&�3+1��+�pC7=+%X=ۗ���L=��h�E;�LA����<>ڼ���<��8=Y�*<<3�;�r����;3,:��ݾ<A�=���C=�$Q���к��Y=\f����<�=�i=r�H=��:<�~<��.�Cy�<ġ=&=N�_;.�.��M��-<eEx�o��<j@=�'�;��N�ۊ��u=d�W����<�+1��go���~<IK麀 Ӽ����|����=��[9w첼��<�n=.#3��ӎ:/2[�\�j;�P�;���<^�=̔�<��N���<��<^?
=�[[��U��,=�ɬ<=�;`�B=x�/�SjM�`J�<뙶<��z=�L����<\��I(��m�<��=�q�F-=?�9dw`=�����<Y����Ug<��o<߃!��v�����B��;/m&�n�S=��=0AW=%?<;D];��⼘�a=qZG��3`� C<�ϥW�z!�����|:='* �v�����<��*=Ar5=9,j� �g��� �Z�]=��m��o��{!=yc�|�[��t�<��'_=�
=�&<��[=�Á�_Z*����Dx\��c0:
W�<�K𼇦�<�D;�*��c��d]�	o�<��b����W��$9�<�����Q�u�v�?=��!=�Ik=�I�})�%��<N}���M�<��=�d=�"�-;.<E>�;�W<֖?<��ʻ���</FE=�,=ɜB�^7�Z$�<�>�.�t=�K��[<�&ѻP7B�a�Q�¬=5;%�]=��<v�H=x-=��Z�}i�;!�w<�=D���=�>=]D�[I��Zr}��9�<�ί<��꼹�S=FJ���J��#P��v==f"�*�a=dh��3���9��v]<8�T=%
6�6�?;�;3=�%�³3�b�B��0<�������<3�4�`!���^=�+�g{g�I�z<��������b��@G=ˉ���ļ6�?=e�9<�D���yh��]j=�o�sZ�;Rp������w�M4G�� O<�&��d�m;����S�k~�<u�8�z4=�晻��5���=�4`=h�=�D�=�ʃl;�Fq���ͺ�:�V��:�*��-�<����4��gѼ�G^=�z7<-R���0��1"�� �� �:��<1�k�$��<�������L঻�%4=���;�Z�<�
=����p��rb<�o�0��<���<��ot��f=�q�;�{d�P��;��#�Z&=|�j<$G;��ز�� �<��'�o=r�c=-E�<�=�p���fgT=c�d=�z@=5^��5Ļf�?=]Ç�VʼƉL=%4==IB��=�����V�i<ș��T7=���	T��o�<ؾ;�$<͜�;�B����N��v=��;$� <Raq�r�мZ%<��8�-=��?=>�{��m�<�&�nY�d@�<�y���,���q��!#=��|=-��ۼ�p�x���*�Y�=��ܻ��1=W4���TF=�����f���������=�',�W{��չd=��<�D����0<)�:c]���ռ�L=U]λ���<l`�<G7�}z&=A��^l���7f����k�s��=�܉;�:���O=�mW��f����;_�2=��&=���<'�Z<*�P�`;v�N��>ڼ`D���I=76��5��<\�Һ�R<#�<�*��u�)���i��1ļ�k{=F< '#�t(= r=�s2=�}�<IS{=��U<��=��m1����n.��?X�ާ�<�&q=a�D�������:���<`́�KE4��Bb��{�<ω��*�<�Y��oy��:�G�=���b�I���P��ȼ���;�;�9	=��z��'=4}����)=�/=P��=�k�l�#��!�?�����9�(G=�U����<n�O�t�'c-<��=.��<�z;��.=�t��"H�SI����@;Z� ���Z=�|�����<�$�LX=%i:��=�u;J'=��,�;����=�C�	�i��?^;�Y���\O=�k�<�O�</i����!={M�P�=��j���(����H���1�����ش��%���&�9V=o3s=*#c=�<=���<~��;�ya���<=6�����<������.==�*<[�
���U=���;����%<$�=7���|=��Ҽ�X�"=��[=��U=�ה�M��PF<�Y9��FZ<\�v=��==i�8;���<'���aR���)=�/�<��K��l-��<&T<�v==`
+;�禼D��*[�<jݦ<ɯ�=f[Z:��M�9N�;�)������0=� =%!����<��:���ݼQ+=_��I��s�W�te�C�Z��nM=��U���y��	�n\{<�,='��3Y5�3<9���av��	e�<�p�vr>=��k�s��V	{;[W�}�F=�:3�u7��>_p��O�<|�=�#�vmr�^F=M����9�<��ü��*���<�f��o<�'=�<�74���);yA漪C�<��=��M=��������K%=L��<e�<a8:<����n�ټ�D���<fN
:�8 =��:= �n=Y��q���Oļ�W��JW=P�=-��<�,���4b�^���N�<+^������	̼-��<�����;<���;�T��=g�c=�)����=ݜ�hf?�S� �6��;���������<�dq��ca=��E=rs=�*�<*ͼ
4=Մ<��̼���#=���<�pL����N�����:����n�;�;���Zo==��<!�E<���9��/=�S���07�jl=_Id<U�<��)�n�d��c�<Q���#=�?<r��=��=|G�t����<�J�
n��k�ӂ�gq&=��ռ���������C<=�:1��B<a�;<����Z<�	=�w?�?�+��Y%��+ƺ�V�<�,N���;6�Z:�*3����"���'g;��'�Q�m$M�u��<k�<[�!=����������WO�<��.�-=_RW=����;������<�ז��NW;��P<~�I��~=�� ��==����Ѽr�<�P<N��=�!����ީY��=ֱĹ�U�?W=�c���2e�<Ѥ� ߐ��^��3��<��a<v
��1z<��<xF1�t�=�)R��;�{~�ja#=F�F=�n��|Q�;@��<��<��/=T��	p�;��U���E�E,(={�^��=n=K��<��;�:=*7�<O�#�{�h:x䮼0���=f=�6�<�!���μ�|b9������Y�<@���,��[��>�d<�pF�x���3q<#`��`b:]K�ɜ���,��}@���s��q=���<b�6=J�A=��<�ٷ���k��B��J����|<�2�<f�B���B�tݻ4P�;��<��1�(�j?L�e{�;��<l�m��a�6����P���.�<
��<\�E=���wU	=�h	;(��<�:D<�94=���JwJ����{��aa.=����e><B~��s�C^O=��E�Сn����<��<��f=.��dz=�;�<[7	=?�a<u Ҽ,�<|�f��E0�~
l�](�<ȣ>=��B
ڼ��������<�ɂ=$H%<�b�;F?�<9�<�Q^=�S)<�"���<������܄<6H�����=��=6�n<��M=�4�<�~Ѽ�=��;%�3���^�%��<P3�<-���>�=='t��>4<D/=?���D�<뢢<Hs=}�
<�:b=k�a=ƚP��:;=��J;5.�;��<�$B<���&���2zD=q���Ħ�<]1���V="e���Q�K�g=/���=Qȱ;ș&=t�k=��%�)=n�N�O�<'\�;:�q=������<ta�<��Q=�����>��=a,��x=z��<
�'T@=��;x⏼�Ӏ�� ��[#ທU��qd<�s#���<J2=$\:�#�d<m:9�WN�g�@������oD�E��P�:V	<�����j=�-��������2�#=z81=�����>�2==��;��Y�u�-�^���A=`�=ZB�<��<�[d�m��;ljN<)](�ܯ�<��a=H��oJu=f%=/ $=k��<W,=J�=E�!�OΔ<]h����<Gsd��d<���D�]-���=����B��]=���<v�z��Z�ֱ"<�~��!^=x�!=��;5`�<�U�<�mӻ�=/�d;M;��<�;=����Xc�{�p=�J��'[<ᘁ���<=��������Ao=���<�ra<��C�l�Ƽ}��H(���*��l�<	H5��S]�(lX<��<5�"�5���$��;�9H4%=��q��!����<�&=�~��T�v���U
���.='�p�\Xr�J&�<䘑<Vs�<og=CRg=ߩ�<��㎽�D:��
��JTU����<Eڪ;4Z=a3���&�E�L<ڃ��c������<�S��٦���ż��<ohԻ�-���%M<	��<�2]=,)�<��2[Ƽq�!���)=�1*��"0='�,=%(˼b� \x���%��S������!,�<
lQ�K�0=pRq�;�,��ϻ;�xu<�f�8e ��x�;����~�.<�H.=��=���<��d��)���C����%<?ּ�� ;.�����b=���<N��<�;�<g1�:o!�;���p:����?�(=��ȼ���N^=�L<\��;�w�<Z�<?�;�e<m[G�(�������;�|�<G��>�<xmx8�D
�Gt"�d�;��<��<��)���W<E}*�D33<��t=��t���*�<ex6<�k ;1��;��<���;�[�;d�<�
E�-~U=ፈ�RM���"��D��x�p�kڭ��?���xO�����]>��?Q�
,���|u��F��b�q�_�=]�����<[�L=$57=8���,�(� �� X;�z,=�kM=>-x��A<@�:�=O�$��4�x�Y�6����<��/����@y�
(`��C ;�t�<+�!=�o	=���&�E=�K¼���=a�<R����z��<���QC<�"=��j<�冽�=���<J%�;=�h��9<N�
@�g�h����<�����c=��r����< �g��eO���l<��<�gj=�x_�ZH;:����A�<�r�9�`�'FU=�G��!�<&ݻ�Ǐ�v��U-\���U=d�0=xZ�<"����0��䧼���<���FZ	<�[�<v��6�*���H�&����:���<I�2��d��I"=�
'=@�F=��<���,�:ݠ =�<ؼa~<:[u�{�� 7��{x:8�<�߸�����u`=7�;�=��K����h=������	=�N�<x`�������:M�5$�u���@r���z�<��<ߦD=75�5f�<,<3=,�;�}�9C�^��"O��C�<����d�ݼ
��<��<��=Y�<n�=��艹S�R��by<��2<���<������Z:$�o=�z����?�="������B[|�r��<ȕL=�<d�.�;B	-�����S�`�L�N=f�'=<n=1�;*OI;��;����<:��<�)�˲0=*�1={Ǽ���<.��9��=��=�A�t�<mg��
�=pJ=0�<P���AG���x�N�<=&95��,j= ��<�EL�;;=��G�h�?<lU�<�<�<�����B�fd�;�� x�� �{���;�.=��=ne<'\R�J�����WK=UK2�lxx�o�=�X=�|弶w�<a��<;�<�7Z=�}�B����0��6��$�<��;=��:�ˬ1=��=h=d�r�S�R8 ���c=�3���dO=C�;� =SO2���U=�= �<f!�_���<�����	;��<��<���<,Xy����טw;q<I�����;YM;=nV�`n����<�"�����'ļ�A&=�S=߬t<��7���	=�z����L���+��wS;��=s���~�&�[Mͼ�`�<]�;o==c����P�;6��jJ<�a;=CS<�Y;=	6���a<�J�<t	����I=҅�������R�z�|7����A�B��<�M�<�<��=]Ը����=�.��w�ټ8���� ��p���=x�:=S��<(=D`*�e�e=|�0=2E��H�<\��<���<v<�D�1J�<�W <���=��?<�S�<��<�n���+�{}=�==�Tp�Bɭ��4�����;�髼�[~��$j=��%=�q�<���l��:�nJ�����Q���Cټ�W���	=9?=[7�+�-=·�<�m��v�<i���=�X�QQ߼X�m;=�[�2m�<q��s�V���F=V�j=�"?=5L�����:�����߼���2�"�v_7��	$=�7[�O=G�1=��S=��v<��Ӽa�Y�ϥ=��b���=������<��9��<N"�D�)�x�<���=+=!�`���漗I;�I=Q��;B?�;X�==(T��<��D���[��c���?�^�y�T�K=�ܡ<�l=���<6�T=�l�,$�<��(<\�$=Kr��%YJ���c<<0=�� =拷9�B ��%<+ "��n[�p�Y���/��������B=���'�c�yӕ��@=���y/2��O�t��,�-<�d�;�k79-��W�J��uż�:�<���º���<����F���4�T�"���<J6K��<�B=��^<㕈��}�<n$�T�䦹��t���(���)=%�<������=d�L��8=�I=]Lż9x-�׵Q���M=ե��r�;�j*=S7;�� =b�����=#�d��Q�<^�]E=��l=���<m~����UU¼�$T=^�8����=d�\<t%j��<8�������+6�̏�;TX��,�z]O=S�C���9�v"����s�Fx�<�Z��U!�5W=�2ɼ^6Y<�~=�2�<zD�����#��9��<f��<�^���<T�-����'�=��g:d_�)�=^*H=	�*=��@�9g�<$=�7��I�T%=�.=i�+<Ĉ';��,<B�8=�P�xD�����L��U)K�����el���^��k����=i�;�;.;��Z����k({��@�<o�<�|E=�Q:�s4��.3=��N��=}�f����7Fμ��= �K=���H�;�U������2o*��*g<�+=Uä; �<�"<���<O����#�i��;#�I�\�{�ٔ2=}�<H5V����� J������M5<��	<
�4�>�x=�B�<�y�;Z#=>��;+��tYu�Im���t�?yD�#�.=1؍��(/��g��4c��$0��� 8=���;zN�;?_r=��� �8�4�	���g_�=̌�:�Y=C���z<*J=5|k;/YG=��)=-�Z=|'N=��D<�
&��sb�/r��O?9�H+9�D�I�O#K=�v��,�u����/�CW{=$�����<Zd��/V=t�;�k��:�c���;�yN=ĭ����;�<��Y��$�@��=B�;��̼�.�;S�<�]�;s�<�_�<���w�=����,%=&�e=/yw�_�F<�S=[y.=���3Qp������i�L��<��M=�S�����YY��i�;�,A��л�FU<[���o=����T����B=z-�=�H�X�S�Sss���<��#=�^l��m=L��<Tӟ;�c����<��T��<�=�GL=kp�<��J��Ҋ�cH޼R6��F�Vˑ�ŘT��R=�;��@-=`�O��H�V������;t����=��L}弌lh:��w��~;�8ջ�k=⢔<���oj=��(=�xq;*	��$1=T��<��;��R=6*+<�R=`�<*a��'7��tU�FN�<�"=<�˼��u�;�;=�$�+&I��1/���=����[��<�c�<	Ҝ<&Tżཱུ�l"9���=��=���ߩ_�A�t�4���[=��;�=���M�FEֺ��<�q�*��<�D��M�=�6O����;�I�<Ӎ���;�W�;}�<���B�<�aR=���m����e�:f����8 -=\ r���z�-=�&E�������J��)�<-��<�f�=,���=5�!��u���s��&$=�d�N�v�<1ba��5t=򾼼�D=If2�C`h=N��g��W
;c>=�1� ��<0�J�/ ��`_;p�M�(K�2�Q��85=���;א]=)1B��Wڼ3%���b<�`�t����n=��I�'�� �=��=�_=��
=��;�#=n����X��y�.�����9=��f�`h�;�CS=�:W�==@\A=Py�i*= ,����,=y�ȼ?����(�<jU=k*<�w5=��=�iZ:�ټn��	�ܻ%o2=s�D�us=㉘�f~=�4V ��C�mcR��m�;�j�<��:=�~ӼG�=Z5=b�I��Ҟ��]�PHm<X�=yk�e$���#=�g:�i��v<OA������Ӯ<o�;͝�<�^X=��:<� ��+P��=%x��ͪ��VC��W���J=$����<?�<:�=;�)�;��<��<�_׼��=I4��=�Iu=��=Y�׼ %`�=D[�;��<�Y5=�M��:=��\�M��᡼��q��奼�>S��]i�v��< .=�N=������<�w�:Z��˳�<I�'��<C�T���;o�<�M�<��i�Qc���으yb,=����du,=��<{N�=��+�c��<;N?�m��;1�X��g��<M=��=4����!��&#=�K:�W�R=�#ݼ�Ǽ��=�Y���$=6�<�/�A��<4ю<�#-=N&��FOf=�L;-&={6�<�B�|��S64<��C=�������u\�<��=r��5��Q&�<旹<{1<��.���߼�Zi<$�&�!�$=���i=�/E=�MM=A�M=C9�����\
=V�5Oe�Tɦ�IQ6<@�����*=�z1=���u�M�p���=;�l3��W:=��%<��;^!=T=E?M�ҽg=8�<ǔ�<TGp<��<R�#�[��G0��G�<��<0l��60� N<`U0����9�;�0�>d��Rμn�5�lh%=��; B5=T�*=��(��r��|=G=<�J=t�<'��<�K��~����:�$�Ǽ%T;>o�H+l=��F=�H���C<����xF�(]�;�y�r��v���g���<Z�=��=߇O<�˼l+<@f�I�2�l]<���]D=�u�<wK:��:��<�mj���N���=�U��ڒ�<[�e<QS=qk-�Q˼zbd�h�<��Z=��3��qJ=��Y=�P��`<��3X��^���Z��<8��~SԼ�I=�q%�� =1���B�<��Q���]=��<��
=)���')�&s>��V1:�tW��+�;���<=2��!A�<R6p��x�~%=�⻼�j4�gan<��;��U��I��/�g-�f=�c����<6�+=Dt�<娉�&�a�I�ܼ>i�<�BƼ��^���<�^=&@$�����Y��[M=VJM=��v=���<Y�|�����@� ;_��<qs���[=�SR�h=C�ۻVw���5#�[�l���<�G+<a$����e��<�=�8<.N=v��v��<V�%������2=M�6=����Lټ��μ�-=N���::�<½�s���.9�+��<����~���ۼ{_�9�ؼ!�(=���<�^�;�B$=��<@�(������K=�D	=��<تL=^{��μ�X~���F=�xT�o����<U��;)d=��	�d�<t��a=<�Ȓ:/Z�x�¼K=Y����=��,0��=:`�X<�<3��<�K����<������4�%����<-�����r�=�۲�TY���<}Z�<�^"=P�c=�c=����=X����<e��QL=��2��Yl=_�G�=E=��=����j�h<��a�9X��B=Ky���S	��\�7���.�=��=i!��
�4=���?�jP<�V�<Ĕ<�7׼�sj�
�g=�.߼��.<H� ��g��j�o�d�.=a���s��==�����P&=�t�<%��8��4=Cc���K��<=�v��ſ;ϕ�m}��D��!ּ�-z=���02Y��X=9&5��U=��_=c�7��u'��i���G=|��<��O=��>�}���<�;��Z���`�  =|���O=(p0�R��;�|��´~���J��W�oi�</��<S��<���ԨX<g:;y�>��<:;t&$�� =QJ9��Q�g	=~y=F�8��(!�l�]�&�<Ÿ?<?�uIܻT�0=��b�T��#ؼ��R=f��<��Ҽ��Ȼ�W<��T���<<�H�Db���+�?��v�=�1=����G��!�7=�,t���=�0�w�:=h"��u�+�=]��[�f�Y0��l=�q=5��<ٟ�=�0O=��Լo���C=�;=��W<ZNH�9Y^;ȋ�&�<��>=0�g<3̝�b��<��<��5�^��g�<�Q=��W�b ,��	�<�L�cIp;��o<�_\<Fڼ�8���X=6In=5�=���<f��jCK=/�^��t.�0�ż77�<=�H<
��=�Zּ��j��˼�Q/<�+m<bg�����<�(��wB������ =#�S;�q�;o�h=XL=�sE;?�4�y�=�ZJ<$����80=�v0�x=ft/=/�=�=��{����<$�Y=��{����<:r[�n�<Z��;���;��n�ua>�48�������<��p@3=���;��"��&��_��p=gI�<�[V�W�o��[���=�|!��	=܊B�����MȻ����/ڻ5:�<��7���<�t�J�vuZ�+l�<�����3=�=�]�����<Cp	�E]\�˶�<r��<� <є����c����_��9�0�ݶ�[u=s��;3�=*�v��h_�=�\�W���n�;�'���y��,��@� 4O=���9�@=n�ټ��e=�r�\e.;�o��YU>��=�!�f~�<��j=�+<�����E^�����n<ct%=�
�O�ѻϽ�<�Į;�'0=>�����<�<�I;�=�"�'l��&�ŋ[=��5=4�A=�	˼�� ����<~=�6?���O��sY��5��˺;��]=���;ս�<��׼7橼���;�R?��2j����CK�*X��z�<^��n*I�Co�;��<�O��<��=}�n��c�<�ڮ��=WH��s�x��=�^�<`	`���9�q�)=C��떖;/�`<@ �)5H=_�=��D<�&�;��&���c3=#��<�A�<ch�< ѻ�\!�rz��V�<F�N���=~7=��Q��Z==O�a=�_=�=�b
=�=j�>�G���&�|`ͻ�w��|S=u�h=jT=�kL<�4�Z������<�ʵ<�ê�����B=�<.=¼�(,<Jg/���A���=�U=�0=�f�Gl'�Y�X��]ҸΈE=�~ټ�1$����1��<�,�<  �<����<>����L=Fǁ�b	���_T��<+Y*=�t�����Y�o&=H}#�Z�o��q<��+�ݯ��V�3=qS���K�<��+=���<^
=�<=�/�SЍ=�"�<��g�!�==B=q=[�<DW3=1���e����g=�������H�='8w���\�0A���<^G�&=<���<�[�;�j޼x,C�3�%��Y=�F%����8�S�<!BF�yD�s=K�;�<=���<��<�f	�aU==);��FY<��Y=I8���ة�X�	��'�X�׼�q��2��7�<Ő%�O���-�S���,�Ł<�&�����<�Ma=]�2��e�<�?9=-�|<ż�������<���<$]&�0?�;s}9�ׅ=��m<J���)Z��	�йS�ۼ�r =�;RO=�=.�=m^=��:�ˍ<Or���=C��<zۼ�&=���$���:����<����a7=a���qC=QČ�!�]=--=#^0=)(�<��f�eYK�;�Y��e"���4�n (=.E.=���=)�<N(��x)�<!�<Gż��=�����ȼ�|:��:E=-�z��ݓ��_��\.=�Z=���O��;`A2��#8���̼�MF�+r�t���o�G�Ǻ�-D;��i=�_��h2�<8�A=9M���_�:a�&���¼���<��
</o��0�<i<�<k>+=�>L=�L�<�=Aκܒt<$��<��<����]��Q={����%��.T=R=HҪ;�CG=���<xH���=ȏ��D�1�={`;j��<z��P���R={[��V��<�[=|5�OJN=�f=yK�+�n<�?e<�A��dX��-Q�1a�_=��;_׼<4�;R�<�C�<���fq<~�)�5D�V˥�_��<§ۼ��P<���<T�=>��<�����,=��ټ2��V[[=���<�[J�F��*=G=
m�;�݇�Ù���1�Z=�T$=�Į;K/��8��;�T�;��ʼ80��e[<=��:=�o=��I� =�W�T5=��<�o1=k,�F��<�4�<�����傺�f=k=%<-%k=�i*=P���i��JN���̼9�g=?�=]�r�7"=��c=�����bm=��0=K���!V%�O�߼D�����Y>H=��<�����Q=�,J=���<#�H��S=�V= I=`R�:��I�aH�;!J=ݶ��'w���><���<=��:��jI=A��<��;=ЀQ��%!�V�Y<��N�����B=�Q�<{����¼d*�<A=�-˼����oX�kKH=I
�*;����<�<)�=<L�<r��L�J=}�2�b�I*�r�.���J<�O<~ز�M�5�S���;�<�H=q����HJ=��N=gx��	�0�?E����<��G����=p��<����c���C=��v;�f߼�.�&�X=GW� R=<�(=Ã�<�X��Cf��R<2ip�+\��'1���=;��<����)?����<C7|���gR��� �<���X�f� W=��s��0�,��<�o�t�<m�u<_��*�A��;@���M=@~�<���<l���S;���{�{� <}(�;�i
<�X�<:X�;K�U=�E���2<�Bh*=R�=Է��G�뮁=�N>�a�j��rR�x���V�7X�<0�=��`��g�;[�+<�?=%%�_�5=��@=V}�����T����P��1o<I�6=؏E���������-���đ~<0�A�lz��qa���;�b]T=�s��	��0��v�1 Q=��U<Zq��Η������E*l���A=u����;�^g=!h�:g#�"��;��b<vW(�:�<ܜ��P(_<��;�L�>��;$a��h=��<��w=��j���2fk<g(�<��;1�9;�H =߅��w�<��)=����U�U=������<d�=/GA=CR����Y��<i�=X��<)C=X��j��~!�<�1��t4�=�>��XjS�:h�<=�[=��C�_ܵ<��4�4'�;N���ˍ<�&O<����}!����<n��ڈ�;)j�=�[g<���tP����Z�y�T���x���<?{\�������O�-�~=����Z<�[=:��<2@]�X=�{+��K�c<�<E�=���<���Sz�<�G¼������9P�<�֡<S��<�ث��	=g14�ֺI=k��;̸=i�#=��E���;T:�<�<Ů�|����O=��߼KG���=ơ<e%A���F��BP=4eC�(B��{P��Ib�Q��<̛\���g�#�R=�o�;�}Z:�X#=m�;�eϼ��=R�d=DD��{D=C��;��=h^ �YLc���=�[P=�<�ݦ���(=��M=P�$=x��=e�;<T;�+I���<�*�<���౑<�W���I=��=V}�k� ��_\=u`=�ػ�z>���<V�;�Z=�:Ƽ^ʧ�oc��%<�����I=��g����;d����*�;Y���.<=���ٷ�Y=��w�=�,�<��Y�6y�j�'=�e ��vP<Eb伻 :�sLp;$]�<�J��d�����a6P=!�<�9�7���5� ��r�W=�j�����<�;=J��<h"<���;�	;-����=�·<�Ǩ�D���N�h��;Y	��.���C)1�̣G��c,=������<f�#<2|(�d=�;=�P=q���I����FY=�wA��9=P2���ͼw�o=���;�ı<�-_��%�;
$_<{���3=�F=��a��K�<��<��m����	��a<�q=t�'=�>S�XF[<.�=�I;<<�Ҽ�a�<K�x�+��8�)=��o��i6��=%�=��b�0� �K+�<��<ڌ�=�,�::�]��!G�`�\�0�޼�>��\�������=B,
<}U$:'��<�}���<@3�<B����:�3���C�Z_c=deo�r@������	x;G��<�p(�.�@��=D(Q�n������<��9��@@��K>���=����r'R�!0�<�k9=�d�I6=O�a=�Q�t�j< X�<��p=d �;�a�<�oB�Y�)������N�<�$<#��s1���$,:,�"=$�<��X����=�.V=mBh;�-���P=�#;=�䦼�X�<ź�<�95��r)�w�=;��N=�������,<�=�<�#(;�a=Y�A=`�<��N��c<�"^<�#�<��W<�a��S��R��]=h�K�����u�=I�!=��C��X?��,�翤�6����:� =؄3=#F
�����}<<�"=��
= �<jC��z�������<��=�*�4��<�<��
��a<��=�"�;��j��Ý<�b�<L	�=��k�� �<�KG=B�<�c���\��rK�<�*e<���ۯ�<�y=�c��Ƃ<=��;�H/�7^j��v!<�X�L�;.����ü�<9;e;n=��<������A�����[�Fe"<��b=�x漈�s=1�A=HȂ=�Y�<�<��C��B�.z����<��Y���V�����<�?���(4�_n)���~��;����L�<Uq�:�<j+D�f�Q;�V���0��2z�%|m��x<�e��<WX�<�rS=��E<��	=��^=���i=�/O=��8�c=\N=��K����+`�<���;����ټ�@w��O��֘<�J�<җ5�!�J�Ϫ����^�/v�:�@e��!��Q��'=�<<O��$�R�:���K=][��/=�8i�U\=�`<��+=?$=9A	�[}j����<Q� ��U���=0��փ�<�d�J=�8-=�����-<C��<c�a=���;��0=+:漤<U�u�����Eмd�)�0.���<�)\��3F=��<��B�Yo�<xm��+7=�i��ݼ^��^=�<#�.=������<*��;\� ��,<=���V=]�����C�ge���b��(L=�d`<���*o;��]	 �%��0t�;=ƛ��GD�놻<�s=�±�<�M=!?^�+s=�"�l�E=��<��<����+��7t���"�_�0=��%�fAx=�c��ҏ���<������twy�v,��6�;$�:="����l�4"e������!<"s�<G��'�ݺ��F;�f]=�z��H>�:h`���<	u,��!:;��<��<�
��h3��1޼���:X�K��K=!�,��_һ"�K�"�1=����=��y��hڼ�z����<;5_=�Eӹas��2O�%��;FE���=�r�<'F���$<�t�<O���>�]��p=.�ۼ��J=1�3=s[S��C#=Ho�<�<̻=p̼�
�;)��<9�<Vg���w�i��(�.7=��O=�=̄�:e=R1=[�<XkS;���kCb=��<������|=�<�i#��P�z	4����<�/':�|�hw<\p��e���+'=[i�;pR=�߷�%�0�ڤ��񼠃�<�|=���ښ���au<�:D��&
�-4�<e}�:.%������� ��>�< �r_��Z����;����XT;��`�<j a:��8=�L����2��F�:2�ݼ��&=���]=�[|�QzD���!�fw�<IN=/Z=��P=�U��Tt����u��^w<��e��kb����<E.4��d%<��e�@�=R=�L���T�W�F��1����:*	f�%�W��<hJ=��ż������ʼ��<f<'�����3_��y�;R:�\g�p�n=A��wJ<ܟZ=�쎼�_=��<© =rlP���#�F�H�����<]��u�� =WZ:�}�<�	=��p=n�<�'(��O=�~�B=�.S=Y�F���g���L#v�֤B=�!=隌=��=fC���ZԼ%u <�Rۼ	��<ؔ=����\��<8���3l=N8<0�����.�6.O�$�"=*�I�=������?��k�;�!=�hK��bY��<�$=o0����G=
�=�f�;$�������蔺XO4=x$J=��<pѼ�\A�x'9<��D<��<C�X���>�+F�<_f)=I�R�O� <��y=tE���U= b=�W�<)�Y�Ѐ0�X+���=Ҷl���(�0�<��<tP_=�
�Qx�<�Bi=���8��D=�vE=�]�<~a�:��O�=�ڼx��C;�<�;��c�4{�<�ZN����_�����=	Q+��q<�c�4�8-=�_�X�P�T���p��;��	��Ȋ���<4Z���	�ʫ�<�|�|ܼ4	��H=;;�'=�:�$$�Y�컨3`=ܨ�<�]=�z�;D.�u�=���>�@=��������;<q��<ڕ�;��;%K�,�p=�k�=E!=�ZT=�I���Tv���Y�{�W�Q
=��h<`��7�<��=hE�	R
����;��<���<&<V���<k�<
�=��Ӽ�� ��z�<��+��W(�@T�|K=�0���}����;=�%:�%�k=.�d��d�<���<�H��Yoź�7���3���,y<�Jx��ɰ���=؃=Q[D:��C=��߼H,�<s*���P;�d�������<�<4��P\=�f=��M�0j��y2��~�Ͼ�e$�rp���sj=~�G=��һs8=�:E�7=:���d�@����]��̰<4"n���<K�$�E�q��(ֻ5������dxb=�n���5���;l�߻���f��%�����<��t=ް/�a�/<�OV=f�L=E�q�ٺ�<8Rp�k�=�D<�W���`w<�'�Ԫ~=�a�&���&�<i��I���L���X6���U�"���9_V=�l� =�;_Eq=�	Q=�t=x�0���ȻU�����ռ�;�<�R�O��QJn<���ZG=�B"�I�G�9=����a�j=T�^���O���]=��p=2.�Z�I�:ֻ�V=9�`���{<a#��S3�:�6�<��������=< =�gϻ?*���]H=��<��<��G�O�1=G��!���Q���͑g�� ۼ�m=F��u�<)~`�W�����ڼ�X���5L<��=
=gGq���3�<Ӄ9�n���d
=_`9�Ȣ`��x	�����$<&����<Z�M=��<�E=燺��<����Y�t:м���������E=Ӈl<}*��+<���-��TE�_@>���#=p�<�F=s�����5�=���<N�y�� {;��<�m�V�G=b+��;�t�7#=Z=�n<ݳ�<G�<��h�<�ZG��U��V2<��L��.;yc_�/=p�{�K�<�7l;;a��y3=�R�;�<��<7�y<��E�ē`��`H�����
�L1=Y|:��F�9�(=U0|=���/A	=���;��5=4�c����<�6Q=�ot�н.=� z:zj=[s �B=�w=��g=��k=�E{<�W����;���<��b� �p=C=��
= ��;l�4=M��<>�?;"�D��;�:�N�<�Φ;�.=�����5�<��/=�oX=ٲ��=◌=�'f����<�=����4���<���akY�@}�� *&��X�<"����V�u!�G�h<��ɼ�=&�G=�̬��ie�g�@<��*=p��j.�'���a=���<lN��m��S�⼫��:k=�S�;˼hC�D�<oF=.;�4o:�� =;<P���̼rR=<�dS=�.��8�<�N���I���%��XE=�*a=��S���=5�9;q�=�O2<��/�<Hs2<���=p�*���P�r'�<c��<�&���=pp<�
=�8�=�s=̻=h��<�?f���#=�2<�����t+��HdG��:1=�w�;��=l.=V�V<�B�;��<���b0���'�gl��6�<��!�=8����w.=>�����b94��V2=�Q�<��<=�G<�/=7jּ,�<�v"=	�g<L�]�=e�<޺>�|�`=�l�R�O�	ͼ�5=�(�<4<�,�9:�d�׼)�`��#�<K-�_�R=-�<�_�ؼ�hL=��
<���$���4�<��(=Ĩb=ɒ4�ـ�����Yy��=���?)���S�5n�<��&=�޻��� ���SF� a�bc��72=Y�t=fBJ=�$,�b(*��#��XH:�|�<�1�<�  �c�>��27�y�Q��=/hw��9����5�e����:��=��=B9���<�?�<��O���)�ۦ�<B�U��u�<��1=��]�ڼ
==:n�<+.�;ڀϼC2=<��v=(5r��<�hKü�	�L
W�wC=>Z��:��{����3;=��\1�<~�H�J]C:�6=sH�<r��B2�>\=� ;��}�<�˼E훼L)"=�K���<��d=]�n� M=]I$=�
��ƭ<�������<MsZ��'�;�[`�s�6;��@�:=�<g;$=���<$�*�d�2=�o �>�=���<�х<������.�<����rԼ͠����e� #<{�v�!	��;���u;q=����X�<$�h���v<�����=Sb��Jy[<��<�����׺��?a<�W7=�3=������]���\<& =9=��2Q�k�e<f�{��p�<ZV@��!|;
�<FsT��̟<�q��>г<�9<ӲԻ�Հ=[st=}�<=�q�����W~=�w�<Ւ`:�;:D��<�>�;��p<�%�}��<��}=/,��o*8=�)$=t��;8�K=�2^=
&�y�P=��C<��/�����=��;z�h�{�7<�9=��<�0�<WW�;E��XG��������=�hG���l�hR�Q�����Q��	�ė����;�[��{�2�`�+�|�=hD6=ni���6�<�����%1�Ȟ=�����3�<�?� 8.==D;�8Q=�R'�Ģ=��.����<���<�kN=�?<W�4=����=�& =�g�<�+�<@�T�G�=��|�����)��B_F�5T�<4�9��|�+����D;S;=�0�i�<��!������ �F诼I��<ԫ�Oi��)V=�PI<b�J=�<���<�R�<a
��6��Ȅ�7[#��]�)=�<=�W�s](�4]���V��
�<d�<)�i<|2�=˼�_Y�f�u���6�~����;��0��O3��ػ/�<c�<eVM�\��������;�\���Q���"=��^=#=z{$=W�u=#6=I���� �p�/=:�@���<�mb<��d��r ���.�A�%=<�#�s;�b�)=[it<�S	=6>5=r��7��=ѿ=d{=0=-ň���̼7��;�䑻n@=s�=�B�[=A�ŕ�Ř�<��-���c���<<t�;L�3s=?�ɼ��� d�u����c�u<��<�<�?ʼ�F=�$`=!�D<�i< r}=���<��^= ��֫Ӽ��g=���� =&����<�=n~���_�<D�^=�K<��Q=�p�1��ዼ��P�c�+S=��׼��b<�^=e	�;t7��>=hzq=PL�;�z=<'���.F=.�>�)>I��kp��1<=�Q=��<��o=Z�G�?���.�d�I7�<���<��A�����;V=�b��S���R=�XK=�<�� �v4���I_=4�P=,W�;�*=���;����3�*�fk��y
;��<<�)]��cc�� �<�.��s=3s����1=R�<@�P�����3�<&�1���<h�s<kd<��<�n�<�C6��<T(�;�&�~˼<�4�<��v< �[��냻��;)��<R�L���1��%n�F�F;4Xܼp�A=�BZ=��L�Q�9=U\�<
��<�+0�'82=o)�;��,=�=���@=��8�zF�<�q8�	F��6q�êW:H�S<T<�a)��_=�����'q=-��W�<���}�`��;'`�<��#�T=g��I:O[�����G��<�Se<7�A�n>t<�r�<���<����;C���\=�h�<컹_��?�<��5��A����T�5�;@�;D�~���|=3e0��IB=;C= 94=��I���)=rW=:H�1=�a��h�<�~'={=�6�[�a=%��*	���<	Ͱ��"='��[��<��i�8�<6�!=$O1=8�<��/�2]ռ��ü,�;�v����<�!��^μf��^J��@�9��=)!V=���=�uy�HI|=l��;�� =��}���c<�s=�O)=��M=#�7��2=�n;��B�'�ϻ� ����{��`y�efo��]<	�=jj_�5梼>�<>�<A R<��̼
�y=�
9=eT���D�]Yʼ����iZ� 	��G�<��<�}=M�T=Ħ@=A��;�30�_����8��:ؼw��;I�'=Q��=�=�����t9Ǽ�Է<W��y��>�ǻ^�;��Ǽ���<�6�<��C���<2�A���<� @=�[�;��!<�y=�<��-؁=&'�X��<���O=r�Ốd=�n���ݻ�r-����B��H��9�*��};�`�=�vj�?����<7����;���+=�7x�┼nI�<���;��e� �==.�	��<��;�ch��#I�����<)�6=ߪU��� �(��<����8��mp<F~m;��;�����5��)�--!=��I�q8<�1�;eJC=��ֻM!��c�Y�J��<8��#��6:��:`��2N=\.�;�c��֡�^o0�#vf����<��5s=�[��=�0	��]�<Ѭ
<{!���;S���B��<Ķ<�M�<1���!v<�l<����W��;|�<]�-=ӭ�<���<ә<b맼=�Nd=�E+=	K7��&ϻ;Lٻ+$<��<�l�=��j�W�-=��=!6���/�<�,���so=��<{,����'"=��7�8Kc<
�7=c)=H4������k=����ʌ��ql=��k��;-��׼�ܳ��ف��L��� ��p=Cn�<|h=c��<��;�V�<B�J=b4��C *=cqx�ؿ=��<�
��ؑ��,6<
�<���<`><ps�<�߹<�u�<5����=�����oH<�4�<���#V=�	;�3ں�ߺ�}<��	����<E�#��]���+=US�<@	�<$�{��Tͼ\�;��<���W&�*GL=4[�<m�H���s<E�ϼ�>#�} �:���9|��q� =�C���L��۷��iU��ڇ�8[q��7�e��<U�
�=0�;���Q2<�-q��4 =b�r=$�����<6�=�f�<S�Ƽ�d)��a=��O�<�N=�����W�;�0�^^4��8=1h!�%^`�&g�<�$���C;�}���(�ݖ�<#�<k��==��<�Fi=�M���<��<�мX��<��¼�,��𿷼��.�3E�;(�<�+Y����?��<\�]=s
�<��8^˧����Jü�:�M�d�S=�R	=��)<��x�S��;c��}T����T�<:Zż�
=kR����ļ�C=��1�1	=�[=�f"��E��vk=�ѧ��?<oŊ�g�x�!=�\�<|+��t���@�3+=0�᪟<[,:��ً�ЭV�52<dB�t���u���I=�[�;��<uJ�C��tI���<=�Ɵ<��=�#<|�K<Q[<�Q��w�<�})�&�G�^=�����~��<ֈ뻠`#�;��=�ut=����'n��5=�=��1���F,��4@�p����U�E=�V��;���<a,*���S=�1�=�s@=)r�<��<�8@=
�y�
�<�BP��H:= �@�'M���b�����;�u��8E���<���$��<3�;��N�kl&�T�=N��=�yR=�h<shi�@8��-L���<��3=�4�^Q�<s��=Iv5;=l��;oR=�n[;d��<Ce%�;�D=�^��}s=@��<u�
<��F=&�<ī3�![��u=�mx���g� �\<[>�I�;�	�n-�����Y�?�@03=��A=�b�;��<�aּ�[]=�V<���<��<;F<W=^�N<J�=	ȼ��(�3=�;K�B=)#;�§<~�Ӽ� <W"#=��T=������<{aq;`���M���[~�z�k�L�J=ݪ�<��^n��	�v=橤<�B|<y�=���<�a���2=f? <�.<3�W=��4=սm=-�<[��<k�<�Yz�����:��	{<�J=�L=��~;�I=�3��
6�@�&��5�<��}=��!=+��NT�<�FN��`<%R=.
=��w<�^;�2�<�����|�s�<���v�9�U�>_;!��<r�<b���!.�>�=%���Q�ܼmL��M��l��i�<O�M�=�5=qN�:��9���;dϣ<
=K�<��J=q�;j��������%� ��[�<��F�/�;�����,���޻|�;~��:+E<e�*��*���)׺�!=�>�<�ep<F��:�p@=gk<��<Փ;�l[������D�;����i�x�\��](�-��<n��^�*�c�,�28=tꟼ�YD=�c�:���>�<����ڙ9�܅���b"�#D�<}��b�YdX=��
=[�����<,�<��Z��:`=M�P���"���!�`�x��:�<�`!�O�I�m�<=��^��),<�=�&?=2�^���%=aZ=�Dú�6�<3l<l@�<%t<���7�
=T=�/ ��K=�31=� 2�"@l��H8=a~V��i��i�p<C�r�/Z�<0g޼�4y��?��zu=������0���ɻ�
�<��_=�F1������=ɸ���<N=�UL�^~z=�V��:`�P�ּ��%�{;<�l<o�m�
2S��ɨ�h�0�-=0B;�/#�<�g(�#����A�<�C��s��<��=�ڔ��=�}��n��(Bk=�<$L��U���.]=���͖ļ�eo=���d8=��<4��e��<�3��tJ=awj=��n�h�8<بD��3���P<ɛ*;���  A=/ߏ<�0>;�҆<{�C�0=@'Y<y
=��<2����]Ἓ��<د:��[=��8�nE��<��;Բ<�@����/�X��h���S0=��<=,�<�1,=8�L=��l<���;R�Mʼ2>� �%�=OK�؀5=^ ���N����<��*���f��3=cr=ȓw�L�o<���<`}r���2<��s<�:k�KgR<yY�<�F6�.Tk��⺻��:�t��ɩO��V��?����7��i�=9��6O������3=<�闼gC���ci���5<�n6����<4*=���n3=��M=�O���zj=�U�;�<	�M<��!�����K
=h�L�d�7=����?V���Ҵ<��=�xe<.�)�I��
vq�a�2<� P�@=��Z�ޯi=��={}P���1��c<t,<�t�Y����;*�:�A<=��B�=Y;���J�q�Z<��鼕uT=5�@�u�+=�|���e<�i =μ���s��<s��X���Y}<6�M��3�9vb��?=�ɑ<��};����O=�d=]7�7�Ƽ$�ι4�Y=�N%=f�H�~�=��,<�a(=[]��ٍ3�����!��A��L[����Rm=�f�<y�2=Y�C=D+��n�����H=?�`���D=��8��V���"=�����=�u<Tc=���/�H��3��m]��^\���H��)�>���(�1=E�|X-='!��o�<*1?=6QW=�3;�%�<`�8S�#�a�tD�<撅��u"�#.c=R@=��(=G�4�Q�=�
x=�]%�1�?=Cq����W=H�#���;�Y)໓H���d� ���^�/<�����kM�=��=�B�<�߈8���?#=j��;��Z��z��j���f"=(��7�1�ڼ�T=�
 <y��<�<p���Ҏ<�!p����<�*}=��=�s(<��Į�;�ኻ���<T}F�
�a=�=�e>=��<��=t"T�>:�;/c��,z����2=�����p*�;l�:���h��;6g-���9�ɱ\<1�<xD;�� �<�C���d�SF����ڼ��h����<K���S�s��kL=\6���S�\[k���<Ou��{8f=0�J=�XI=����B��<�W��Vm=#�*�ǈ�P�5��K1=Y.&�� :=�i�8F4=#��-4-<��l��]�C��;��V=��<S�-�-�:�~;g<Y�T=N����Ζ<�(=���<���;���<��=���<Z�U=�9�#���<���<q~I<h+=�F�aiY��4=J�'�XX*��s<��h=D�T�ڠ�<��;M*B�W�������g=T�-��VO=�e�<�9�q��=}��<<�&=�==O=��L�g�lǧ<LZ;�P��;<`�%�qt9=ԙ�;�|Y�_���cb<�c4��Yo��?����<Ȓ�AA�=Pv#��}�d�=��x�
�>�,y0����;�%M=*��;�J=5"��z�<z�+��7D�@�2<D��<J,e:k�����;)�Ƽ2-�Z?�!6<��r;�Ye=�'2�P0���٣�YQ&��ؼ݅� =�*��Ju��F5��ڼ�-<��:�M#:�cJ������W=^%<�,̼s�$=\S�:�y=�D��{2�<��:C��ӮO<������KT����<|B=����=���=�\+����<��;M7�<^	�<ˈ<��,=�)�;��� �{���;�ֹ3=
��_�|���M�<�X	���K����,���:;�ƍ��� �<д4=��l�<�M�<��}��ͼq�{<����[3���=���#\:=��ں��6��1�<�d[��E=��=5�=�=�<c�={���<�)޻�m����=���<c���IQ�<:;�Ur�<Z�P=8�=i���u�<�,�y�<=��<thN���;�休c��m�G�x�s���<(�X���6=A�,=3p��2�j<4ϼ��8<e�Q�����}�=����Ɂ=�M�Ĝ)�1Y==���� < US��
=�>=����yL=��)=gp�<���<��=Uq\<��׼� ��e"=��H=�=N7q��jC�#�<� ����-�=Z��:	vV;j ���ݻ�?X����;�*�����U�:�&�<�eV��k���Y�U�B=(�𼐅�<����ت	�6��ϕ�<,�d��;��<=!h���<=��S�|�y�5��q=;�'�F�)j��|;I�/=��<������ͼ��R���h=�<U1=N����E=�}�;�7=T���M�<�i=�2��J=��B��I�;�WR=���;��8�����3Ƽ(�<eq&���<�n��h1<�ԉ:��=�;g I���?=9o�����,o��h=6�����4=
zN��#=c�7��I=#�~<&W�<͌G�گ�8�5=�ᗻ��t:�=g�<rW=�G�9�<	�5�h|��9\�<�'=S7��P� <s�-��	G=-U�<}@P<Z��<�>+= ���W=4Du=�Zȼ��#<��¼���<n��<�k=�F�:FG2��oK=��:=Ia;3K=��K=[�Y��-����V;ͫ=�D�:U<=i�k=�<�<Mw���21��%�}�;���<c�>�m��<#�=��<F�{<W�C=��a;Q�T���O< �Y<<`�C<�Ê���T=9��</��UzP=-Y�<�8r:J7�<{A>�A��O��<	=6<=�]��8X<�u=����C�����d���Y���G��.(�x_t�Iƽ;{>�tg���}{�k]������a6�}w`�3���g�<�%�;��w<y�����;�Ȑ�T�=bxJ=�˄�zI�<��<L]��U�}xV� $#�̉p�c�9=�)ۻiL���Ǡ<�8c����;��= ����X=q��=��
=��p=ӏ���D����H�,�=��$=&�1<�&�<���<��̼��<���<:�D�ڢ<zC=��J�<
(�Y�;=�9�̂�8�j<��?<�s���<텀=Ϩ��Jm4<5z�:��E�w�< 7i<}C;�CV��
��fH�=c�1���ƻ���;�F4�|"<gp�<�(�x��<m��u�^;�n-=,�1='��g�<��<E�<�B&���(��b$�f⳼0�1=���Bh���c[=\�<�d�;��=�l�S앻J+=�3�����
�;P��<ȟ��<Gぽ(`��w;��p��<�V=1��;��[=e�S<��.�4uH�=)+=�aD=�{=h��:B�&��f<��-����=y=@S=YX�SG�<G.N=��:9�5=�:'<���e���j��<���<B� =�=�;+���"���=�e���tM=���<�};E�<Zq��Ćռ��JD���6=g|��+N���J=��5=Ќ*�vv�<"�J=򑖼�S�<rS�<�O��ݼ���<h�|�<�O�<-�n=�#<t�L��`3=L�	=,/$�ح�<�g���=�ü��<�1=�7=%��<�	�g��<w���:2�<�f�Jj��h������� W=��F���^��y=��>Q�+���^���;)A�W���Q&8=e�W��=A��<X��O{��4(=�녽*/ּ���<��"�e��<�B?�bK�<V��<#��<���R�=�&=u�E��DW��j=Dϼ�xa������
�������=���<�*H��'��=�4~�~�=���"ɽ<�.:<�c����[��!=^%{���<W	=K^c���(�I��<{��m7}�/L�<n���k.��_�!���,=������U=;�==+qt��0��<ȷn�P�"��/=J���1<d+�<./�<>�3�*����qK<�.D=(�}<.]S�!�ϼ�WP<5�Ӽ�@=ŁB����x�ۼ"�
�}I�r�l�ge�3@����P<�`=���<j��t���/�5�%7�����=�� t8;��=��E;J�Z���0=�\9�=��=�/�<��<��ʼ�<\=1�(���ܼͥ5<%�=�����i=��P<\򼌪�<��f�=�)�/�v:��?��r=zR=i������Z�;����<�6N��Ɂ=3=|o�1(,���:�(=�q!����5���zG==`��=.�Xռ�ݼ��	��\ =h��<�l�;��<�&���S<��i�W�C<Qy���=sނ�Lຍo��f�;l(=JP=��޻�@=zf��Q�<�;�=8����;!.�;c!ɼZ�/=+�<�_���{��TO=�bp=]�0=ÿ�<}c�<}�h=Qd	��h=��(=���L`��eټ�޼��=�i,��j�=c��&�d��$+���!=cL.=���;o#r=N���FO�76=E�K=���~��<���Z�,=�|=�#�;++
�`<��]=�V����;n>����'�<��f�Y=S��;�K�`�;}����漝�"�g�s=ͪɼޥ�<��k��r"=Ss�"CW������8;:��Ϯ�9���;F'��,�U~�<�= OۼPW�:CKJ��$����<�\�ھ���<����|=
��;V�K=�=K�L�y�Z=R����\�\5�m7�=��T<F�Y=� ỳ6U�]^�;gK��a���<JJ�<�=�#;��L��9"�ԠJ=(�`�f��D�v�"=�x�G�%<z��OVp=����3 =v�C=*�!���H�P�k<��+��i=�5����;3�<Q���hU�<nUa��}I=l�&���/=íz=2���+���T�D\�<u=!�P��;�Ej��J<��*�$��;��<����0=��A���:=��<e�ڼu<ۆ����j��4N=�A>:G����;=\�kh=q%L�N���'=|xl=�G/��v��t9�U��)�w?�;�<{R��C=J9=�輤�V=�+A=��%��<2�,���ȼ�Z8<7Cb�^&=�S��i�GZ��m���`=��A=�w&=.�;��<�́��O�<+�0�q�ʼGo���d6;y|�H=��=�h�U�=<��G=-oB��,���<�,�@�z=5�&=V��;��b=91=��=Q��+g=~`=e�3/�< �<�;=f5}�RRM<�pZ��i�V���	�ü����I�j]��D=$�5�wZ~��O\=�U,��I9�܆���D�;�)l=$I<��<h�F=��;����ͼ���	� \�+]�q��<'���Ac�^�8���T���F=�M+=y<=��-=f[�F<agW<x1����:fqʼ�5��@�]�Ǭ:Au�?G�����U�&=�2ļkPU�P
�;�����P=�f=/�;���g��{��<� �<ц)�ȳ_�e���z=C<R=n�<��U<�V�<4���(q6;�zk=(#R�Կ�;o����>w<(�%��U<
�W<&U`<��H=
�>�����G�d=�������<	R{=Ɇ�<�e==���;&�x=�=<��r�ϔ��F��M��ڪ�K2=�.�<��^��|�<fOm���<#�T�u�?���=곺i#�9B��<NH�-/<�T�����9����e�<��<_[;=�1T�<���zg�;EG0<�hM�	j�;;2��<c�7�.@=q!<d$�a��<��%��ɻ�.�D����@m�=�	��O=�P�.�A=����B<�p�<��<Q�#=��=��=����O��h�<(4s��<:�<r�<���������cJ�}=�V#�`1�;n�+=�̔<N_�[ȼ�k2=\�ۼA�����F~I� '=	꼈�c=32�<mt`<'w*�Z�
�4tP9G4J=֥<Q�\=�"��1��<���<�:��~D=����y���-;Vך��zмD�[=,�=J�r��<[��hmS�n�<ߛ�<H=��B��-��G׃=�R�<?�]�.�;�u=��߼1� �}��<�`D��M=�~==ꇼ�'�<Mro����lQ=�x=��7�u�<<�;l<�0 ���D���(=�����)���0<j�f��(���Ȓ����<�?7����<6�<�th=��<bz=i�� �G�����-=�<�,<��g�@E����(��#���"=�2;P���JO�Ú �,��Q=�O=S�:=�UB���7��-����_=>=҃Y�&�=�v��	�T %;�?���9<F�ݼ�l�;�������<G)�<Jel< \o�c���jr�4�c�ل�<@�F�sQJ�(��662�m�2=�1��I9��F=
�)���=��ݼm��<f�<ss�9��.R<��H=Yv=(�<�/��>=�L��49�<�d��]jF�u����]z�{�=T�=���
��gȼfxC=O3=Z��<<?���L=�<�A�W���=K����=GhV������L=�w�<����˫<тj�a�o<��p� F6=fI3�lP��ia��ɕ<B�	����<�<�p��<Z���+=c�[=T�׻T��<���;e�B����q��<�J��☼��<h�=X�3=t���Fl���7<FV\=��)���w=)��Cb���0�p�,�4�U=�<�;�s�6� �<E4i=s����<��k<h�z<�X�<�G^<l������I=?�f=as��<������<�g3=��R�O_<<�E6���S��%�`�ϼ�#<U{���xD=��{=J�<F����9���G7�<8�6���r=���7_Y�%*�<�M��EL��=���<=��<�<���(ƻ��/=B�Y�G?���<���]O<��(=��h�<聻O�p��ڼQ�;=�=�&D�{}�<F�x=�}Q���O�M��:��7�x=�Ҽ�2��0��;M? �=犼^�~���s�F��<�P����=� �����<	2&���{�T'h�f�~��_=8Q=��7=ʉ��/*�of����=�E7=��Q��d�2�/(U��=<#=�BQ=�����Z�[�n���\=�^0<O���S�^�O����;�ҩ��7^����Um���;-�D4;=<]<��h�6=}>Ƽ+g�;�m!;$����L=R���FӼg�<*��<Gl���I��Lm��F�х<���,=�=>�d=7P�<g�4o�<a����W��KQ��l�	q��G��c�oW��g&=�9=��軀��U�=��=��L=f��G��;��<�:i="�;<".���#�mX�<�9�9i�D=�+Ѽ�%��*��<%�����<�.��Jf��;�<�'>;6՗<��
�]���n$�<�;�&�k�X�C<�����6�A=I�w��{J�g`���t�y��:�_�	=�[/��{ ���+=�^=��G���<���P�~[<�0�<��=�p<�i���s=D����H�;�1�$Rμ��E�S={�ڼu�D=S�7<�4,��qS<�����K�ݫ��m�=��Լ��׼��h=ʬ�/��<���9���;\������<]:�����Q=�?K=��-���k�3���QG�;ę7��b?=C��ݭ�<!�>�p1�f�ͼ��!=�R�<����FHϼ��Z=΢�<Q�4<e��j�޼�`G���V���|<�㦼M��:.�#=�{���b=#S����N=�s=���.(�<f�8<�q�<����
���<�S��P��������ŶF=��=,�;�2�$�~Sy<z�U��t<�{X=i/��Z=z,��^�=@�<�X\<��E=$
=�X<j���<)�-��n< >�c=���<�v�"Z�<f�Լ���<�d�V�y�q�޲�0�*�tv�{��<��+=ꏴ�ҹ`=�y�<n=�;�J#=;nʻ1�G�L��;�#.�$G=bW����Y�<�9����:�*\=j��;
YA=p�t��k=^=1=oy<6$�<���< =��#�ʬ[�G˻;t=���<�!�<1��D]��X��a�K=6��<}λ���<+:�<��J=N�:�J<�h�;��<��<�j���w��ˀ<��7�D�_�==�����&=	�a����<��=����2S=��{=?�8���L�3	��=w����|_�r�=�=]����}�L���;�l����^ ��/ba<U0�g؀��+=�?<Ŕ�<�5j<Xgh����=hl�Q��:a�!��,(��9<��K��<�O<�2�V��=7֯����;qI����'�W?κ�U=[P�(WH���-=nW<�ƅ=B�	���7׼{�T����<h�l=��=쏣���;v��-<�N�9�C�<Qi=��=8RS�Yܥ��}Z='�<���)(�p�<d���{=6u<aoe=u߼�;�<I���U�hEM<נ��S��2�O=9����pi�r���)˺c
���=,Hi�J�P=ʁm���=H+=�`$=���<,�I��z��];o<�O3�C%W=�P��<5��ؗ��8
��;+�k_üɑ<�<�/Ӽ�>N={ȼ"=��I�i�B�c��<jD=����̶=$t+=�a�=�=������=eR=�`1=6����;ńo�z2��J��&��h�"�<	��=�һ�����gU�ƌ=jCU�;�(<�{S�# J��XT�A�V���<��5����;�5<>��<�a=Qa=��9�˽��䎺���N�O�%L�#�'��^p=1�<�VT<��S�b߼����`�e=T�3=�EC����;��6�w�j��c<��:fbO=ᆼᐺ<�A=%�p=a�=�(=�L)���<H{�</��6�_��[��B��7S�<��/=��*<j=�&�<B~��띺Ge���b[=��p���L=�]5=}پ<�q�;�(�<? Q=�F�=��=���<��Q�v?=��n=DMU=�%��N3<�a���	=�B;Y0���<�#F<�2a=��9�_ޫ;��i�/���L2h=�	�o�����˼h{z��J=K��&#Y�F�b�w4��>��<��.=�g =��k�1�k�)�	�y�B=x9=�`�I�@��=��8<#�7�����½Q=�
�<.�3��n��K̼�mټ�9�\�<��<��<�\=�V8;
�6��'E�π���ͺ�߽<׵$��W+=�=#�=$�ݻ�K�b<��-�e�z,�/	;�)-=�ⷼ�䷻�PA=?�<�5�r� =�y=~A����-=>񯼗+=�&=5�_=����9LO�g���N=��H<k��<�L=���=!0.�R%Y������+D��<��<���||&��84<�
,=�>���Y=eK��Y?�^�o��9�R2=���L��<�_q<��<l0=FW���an<�ü��w=aμ���<�S5�{k)=<���<Ǭ=���<��-�ل��V�S�6�#�-��<9�?=��=P㹻��&�8��x�l��<��G��R�����<��l�QO3=�g����<�'��NE=��D����<�</�*��K=N�/���*���$�:c�G��P_�5�V��-����<8�<�կ;yv��~����<��<2[�:L���cv������<1R�<jL�<�8��;����;��=�m=��ۍ���D=����D=="��s�ɻD	[�0|;+SZ<BU�<&:=W�=<>J=�U4��Җ�vQ
=C1�<��#�yS$=�t��eĵ��|\��>0��˺<4D=�Gy=;�=to>�e��[^9=ZB����<�h)=V�[�qb��?޼��}[�I�C=�e���v�<ƽ�<,�<���j��<P�j��Q��򂻰�Uh�<��
�a#�'4j=a�c��<<EQ��e@�':\�ű7�����qc=�<:3=� E�A�=��;�1=;�7��R4v<���40���n�a�S;c	�����)漇��<[��<8=���3���];��^=������<�Kc�(�};�׼�e�;��=� m<��2_�q_w��u�����mM6;7�=��<�N:���<<v9�w�#=��a<ME�;�0=v�<j�i=�B�0�(<���;}S�/&��»��<��o;B��r��0��;���t�]��'M=�G���@��3
�nF���t\�~%=�0~����0-��3��<R��q_=+x1=����G��������o=�]=��ͼ�:@��!��T�w��G��<��;�a��H�2�КK<C,����;R�J=���<�-��B1�+�N=�\=y&d����8V���p=��=�G:�+޼��Ƽ���:Q7�<fm�;��7�5iH�t��<�J�:YG=��<���<F)D=B��q+�<h�N����<�t��#��;�*+���׼�\*��ϼ�s��Ik�z<=B�C�ڼ�sV��X��9�CF����/=��;(�=�m<���<Zu�<p�L=�fP=gۼ��=
=�GV=F9�L�L�f�=�4<��U=�/���0.<���������8�P9���h�<P[V=D�Z���+��w�92�6=_]м�'��ݼd�=�n�;䵘�pu��c�<sPG���v4*���0=]��o� �^�
���� 1=��O��=i�;=g�9<C��s�����;;�fG��8==F?�(�\<�͹;�=�=��<g�=�z:=D�E��5���l��È�<���<�~T��b�|}=h<+=Q�;���S<���<���t�:<�[����<�Ɇ��8�<|�I=S�6���P����<�z#���"=�?�f����2f=\Vm<}U(=)��<��V=ߍ=<[������(��9��<� <�.<;�B������<[�T=|�=�}��Zh7�=DV=��I<����~�	����J�=�j�I3k���S���o=aO���<x��<Jw|=``3��,S=R�ͼ�
<�<GC=_�m=k���@�;UN���<*��<݇�:�c=T�����B=����K���8=:�a<ۏJ<�y =�{���ɳ<�Y���$=ڷ =�?[=��1=Q�w='��<�I�;���<%�	�~�<6��1_/���"��^��`h�����������7:S$=uջ}s�<�B��(�A=�#m���7=%�R�?�=d�0<7yE=>��;��ͻu����f�YW�<�=-�S=�QK;�w�<�V���s�m!��9z����o=< �f�r��C�<�=�z���Q�<�=�/����U=�$�Y��;���<&�a=���8�=�=ꔼ��M=3����
<�Fϼ�;�삼�{B={�<���<�z�xp
=�+�<da�q��<�6t;�_9=q!��@g��(�zX�<�+������Q=���<����w=D�B=^Q����<�ӽ;T;N��=Y(=�<?�`=T�=k0D����<o(��yb�'�Y���G���=+F�8��~�m�zQ<��V<��j=���; 
��c�$B�yQļ=�(�L8!=�jl:e���~�����<��:=I���
�<�w���<+���=�<SM%��=��;=���;JF/�ӵ�-�0=7Y��S�B<y�\=��I��<�:=]{3<[.Q�݇��R;Z<Zy:U� �7jh�,M�uW��(�=���<��>=���<w8!=l_g=���<�5�<��#��C�<��*�!=�H��̼~'��ñ<Ò���;�&�!<o��;����*���L�;R$�x��<W<�^���k̼���<L�<��M=�<�;�P=WB ="���QZ��#,={jȼ|=������t4=x�G�&�=�=#==��Wa=�<��N~�_=����;�<ZC~��-n�'��~��;��<�Z����3=�ǖ��H�T�1:�z9<$v���7m:���N��<9���w�<��J��X7��D�=I�׻�/���^=�H����v:����Y�5=UYƼa�(=,��:Ô�<�*��6=X�1��5��؝�K���)=�|�6V���[^���<�~�;ϳ�$Η< q=Bx�E����:)=k4k=��c=�Z.=��d=�@=�.&���=�~�
�^��N!<�"���<e�N�[(�<܊��o�hs,��˘<4�Ǽ�=d~ټNd�<Rm��a��]6L=�I�<� ���u&=ĖG��L�<�b>K=���*I"=Ȁ2<�6B<�y)�?=B;c:��Q�M�8��� l�u�R��<�z¼�o:�=.b�k�a=�<�Ȯ��4=Ҽ;�Ӽ,E��q��7��Rr=��<���<ˎ��p�<o�W��O�)�+��/=�&�<�^���>=���<��G�;ʪ)=б��j���²<�<'�<�2��=|��K)u<��w�t�˼d�ҽ;<��=��<�]ɻ�H�<���o�Y�jE^=<�u=��<�JϼS���6<�]@���<�߬��H�<���i�~{�rDm=���5��<�A�4*����;a[=wC�<�+��x|;6�<xz�;rK=<T��CdQ���Ƽ0^��P
<�	=���=#�(��"�)@���+=_�<B躒Y=a��F�<��ʼ�W=�����]�n��3D��2L��F�<��9�d��uM<v�:=��=Q�X�'3<��<C�`=��<-�(��!�,���D~�<֓�<�dL���V���!��|\�z3�?�~�������ʼ��=���=�+d<���7	��Ȉ{<��<��=��l=3;=ފa<�o�:}�ι�bT��t=��y�NX�<�;h=\��<'�<G�T��(Q<U#)=�/=g�>=��3�hg-=�U �y>=��4��K��+	=�m:=�;���._o�7��*ۻ��^��)V=�=��zd�<E�ԼL\��O�k=�_=�/�����8W������s��뼌T�D�8=�"�<e<��<�Y|���=�f�������~=fH=O�*=��<P�O���=7�;� c��6����jΠ����D��h�=[GW<�s�����/�'�
�
m�`�]=W�ظ�]=���<������_�W-=L�Z��*���s��#C<��;�*Ҽ��<��&�28I���Ͳ�T=W��Q�<�ռǖI�߭�<��]=|�d=����8z���Pm�W:��F�<���<v��<�!=��D��`�<;Y�1�I=� ŻwPQ���;>JH�(�3���=H&=�Q�<×��s_=	�Y�<"AA���=d����M �^�=�0n��O�<m���B=���ؼ���;����׺<��<s0=��;��ƻ�)=&6A��Z=�<κ5���(=�ռ��%<��<Wj��/D�;5�ʼi�8=����A����ؼp�;wN�v�=���<��뼷���Dod���������<�#�;k���q���=�RI=�*a=��D<{�i=�)='�U=;M�<U,K:6�k=���Yu=���;<���.��Y����V=W6�<��<?H���Xݺ��<rO(<���H���:���6="����=m�.��`(=]�&��R��,��VSK�N� =9�<��#<]C����<�-<b_�<�\�:7��щr�Щ�<�u_�m!O���N#p��<�wq��H6��YV����2�<�BA�2���|���DvQ=�u�;(���1d�%�;��Lw�� �<�>E��*�<-=�e;4���-?�����pT��j����������^����<~`�<?t2<L��<o&$��xS=c9�<?b=9�<~���<�7k=�Eͼ �7=k�g��q��O���=<�X=V�Y��{�.5������x#��7��VἳP<$��<v�f���5�GN?���+=z)�9�Q�E�(��)?�v�U�]��<�.=�J�3_Ƽ��P=��=#7�<�,=V��;,��=�p�<0��#���G6����=��;O��<M�H<JB�<øa�l'T���G=�a��pn�����x��<;�@����$=s|$=U=i�M��Q$��k=r3��f���.e�<�<��ټ��<��z;��"M�:4��B����m=}�<·ڼ�N�;�2H�^��r��O�]=�<�<y�ӻ`#=��=9\=V;%� =�p��Sa=��B=�кı�<$�g����Tu�;�����8E=���<��»��;�"��#��S)�^�#�e�4��$t��K"=��c���,=��<��i=UQ����<9L��Ռ+<����o�;�	�<6t6=ͬ`�m\�:3b��*0���2<��O��@ր<|,�j���V=�v5=��Z��`��8��4�m=?�8����;�q���׼?!���7!����̮<n�H=& =��<�2��>�-<�@�;�,��.��/�(5e=�8�Dz$<;ͼ��I��x�%!�|!S���<�b^���L;:��<���|[>=.�^��/L�,�m���¼6�<0�B�0��Y�ټ�m�$�A=��T=ASQ=����]<0��<;=r��R�<f�<�Ě��T�-7¼s���c@���ͼ2'M=+	v��NC=�����v9��9��~V��-�c㴻�R�;�bK�컣<�oü�f<\��<���0������_��5=0��<���<ޢ���bf�mge=_P��iO<}OB<��ż7Z;�H
����<~�9=�/I=`��<�\M�������W����d$=��<P&��8F<K�<���<҆B;��1=���;'0=�ge<�=�����<�k(������?="�<V��:\7ٻ1Ѥ;ʡ&�����c����<� �<�G���\�V�W=P�K�����(=1�=Y��:�hɼ�ݻk�C<m��<Z���x�<Dne=�#4=��6�6z����=�4
i��Q�y�û���<�N=��^=8��<tV\�ސ��c�м�*h<[��<�SR=,R¼[�*=�/'��}�<Szp��"%=�|!����;��[=K�����;N�6=�Z=���{Q;=o"ּ�u�<��<Y=�����si�����3,���<=�P �{2�(6Լ�ؼ��;}��%"=(0e�Q�=6����Tϼ��<Eo���<���;j�F�0��=+�Z���N����;);3$�����^ܼ~�5<��-���M<���
'�;��`��h�;���<>�ϼM	��M��<e|V�c�ռ���֚3<	��<��I=��O�t�w�nd+����xC'��MN=�t��_(=��D=a�6=T\g�R=ǥ��qO�Pk��{=�x;�;��?�b鄼:Z�U+7=��"�v�]=����(�<:�������^����:2w�'1˼o�_=󑩼8����P�7�<�R�<��B��0���=t�ɻ�;����o;��j;��N=�m<6p�&�Ep=�|�����<�1w�[@�#!G=�����uo=�Em9����>ǔ<N�H��2���l1����)=��<5wd���ͼ�����M_=�`=a�	���<�R�;S�W=�����vm<�ļR1�<����A�a� f��T=�d����;��= ^��mv=��=5���%=��=��;.h=NJ�<�0	<9Ln=��<}���S=;(��Z	�Ue�<؎�XC<����OD�(B�Æ[=@5�����-�\�(]�����J�=�t6=��<��=�+=���A<������#�;bDg��C_��(�<���;
7!�j�� �'���<��]�&6N=s�=�T6��ӻqu<)h@���e��w�<��<j�;��=�P�<' �<VS,�Ʃ\�jA�9�b�<�V�;l���k������9Ц�՝7��l���=�6���:_=P��0k����Lւ<�W =`�<��׼�ڼ�۷-�PU6�,�w<j="��<\�<!���<	�Y=V5@��� �6=�`=����_����f�]�O��vV�R���+�i<ܦa�'P�;�'=g=�=�
<P9 �Nü�{$��dl���#��LR=�";b)A�ex�<�.<���� ��¢�<@Z����=��ڻ� =��
<�{'=5��<�}</M����(= �;0_����)�T��:����C<�Ķ<w����v!��i.=N�:����c`�~ּN�v�y�.� =w
[�+�X�Y��<�A='^�:E�*<�=����>�Ǘ`=�IE<�p��溚�x�*�\=�lX=r�a=�(�+�6�Ua=�#=�M$=��s���
��C���<O��4=]�k��yR��2-���	���-=��(���Z��B���M�k�;N��:BA(��(p�R��Q	���=�\E��b����=��I�nx:<8�+=�X5=��"���:=��^=�X���:�;�&=n��<r~��q��<��<?<_=.d<�?�r=Х[:v)r�t��<��d=�=j3m��8;�b�=D�4�0M=��<篼N+a=��m�E�*=�կ<PZ �V��3 �A�)<�I���TW=��=^�<����q��L-�;?��������Y��]�Ox�<�黺�.�y�7G�<w�t���(�u�B�F�F�~� =O5μ���<\pA�w�<�S��;���<y����b�<��;	#�M�*����<���m+�&�"=�»=yؼ�;o=�t�<�4
=�*<�2]�"��<�8�<��(=�B6=�͉=��X�~� -'<����m*F�7��,�ld>�'�z9[�м����D.<��i=_���v�7=�?=��E�Գ]��V�,U*��}L�MjV=+y<]�W���=c-ػQ�<z��<�"���m=�K��6���B�}]��H�=<&պ���$�rb���.=f.�<~؞<R�������1z9����<l�;��H=����><���<X��<�>T=�=o���
��?�=��(=��,�8��<��E��@$=0�Neͼ�v<0t�<�+*=�O=��5<=��!�LT�=C����Fl�q���6��F�_�Z�K�eWV=��5��g=��d��y�<�<��:�� �T�(��Έ�1$��73��}��<����G	�<q`��ȼ`g=e�v��s���^�;�b�'�x<&��O�;dM>=�kj=�խ<��<ϟ��Ҁ�<8q�;�	��ݼgȽ�� W�K�4=�)W��υ���E�7H<J긺cGi<8ws<q���:{�<��;ذ<U��<�@=/&���!��l�r�<�*�<p׼�w���b�;{.���6!<c��ױ����üQ�<�-<t]$�D���?�U"ɼ�<�gE=���?=�-��:�< u��H=�J =s�/=�|M=:w5=T%=�G<�R���$�X��]+��-=ML�<�N=���_��3��<T�]<�捼�8=�;�j�����<9x��mqO=�h����w-�D;����<��<4Y�;�$�8Y=�m��g�4�1z<T�<�7��<(~��<:��=��Z���2=l��<�<_�����)Ἒ�u<',<àU<JV=�|_<�W�<T1��@�薪��1$�R����_�;sƶ�]Y"�Z�r���ʼ����c�e2S<9O$�b&+�<��%;`���u$�'<$��7ݼii=y�d=O�=��-=�V��6���<t$�9d<jhͼ�=�bX��E2<��G=��;��:��NY�u�o=�;��[=��C����<� ���;<x=3%w�����u3<
��<�������;��+<�4��>�@�4�|�a={]=�9E�e���=����=A7��p^<�u==��=��(�P�������l=M�\�0.������y�6��<e��<�����겼�>=��?=V�-=��<6N�;��i=~h<u�n<�ѫ�<ݙ<������<�9C=#o#=�"=�k��s���=�=RC�;�6�<��[�M�W=*ZP�==U��<���<� �:��r��/������T/=P�ͺh�<s��;�N.=�a/=ٿ <$_��𦻁��<N3=��o��n�<d��� ��R|��<�!���Î�"�� ��<c'�<8�S=*4Y��쏼	
$;�i=�ȟ���缷�=��K�� `<z�K��OQ;� $�7=&:�} 8���;PX�˂R=r.4�{讼-�N�n�9��Lx��/=h#�<���<�
+=V��<tüэ< ]�a.��U�e=&��<�Y�� ��<�3=n��$�Q<M�;gj<��)�y++=�p��=$�t<��6<�KH��k���:���<���/=�#f=#�q�s�o�9�=$V"=m�`=�1<�y9=qI��;ƍU='a<��<�T�����:����X8=��L�ik�bU$���;`YE=C9=#'<�-�ɺ<_�u��'>����<�x=1�[<�)��%��*��n� ��.g�5�E�xj6�fMټ~M<��|=������a=��;di7�[��Y	���;��9�q�^����<ꞈ���ݺ��}�M<�<�B鼳�l�;>*==Y=�w;;X7*=�=��<�^Y�n�ļ4��}�E<�k#=�*�bm< L�:���[= �r<Z݌<�k=_z=<V�
�7=�ͻh3��{d<�`U=��u<��A="5G=�l�<��ȼ�S=z��<������<Eɻ�=�j=�G=����C?3=e#=eC=�� �%��9�R$=���<�2���I޼�Rs<�|Q<���<�.�wе�p�;���)�=|��<��Ҽ-��:�f	=�#[�̘�-\��?=Pg�<�ѓ��"���|{��@=�ų���=�T�ꆾ��-�<�[x���v=œ:�#e=�ȼf)�:��B��d��2�2z��zM=��F�H_�;�c�yU��1�P<�r�<�k	=�u�q��!y�m���p�?�ɑ�L=!�G=o2`���<�n>=8`��Z�<ՙK��Z��u �<���r������<f�"=�%4���'4=&n�<�J�;d^=j��<�>�B�h<����t���O=`1�ҋ=T��<��C�	�����S��#��_�<���<�%���ϼE�<~�����};��<V�<��ol0�����#���q��ݼR�={0�CA=��<�<��븄q�:�z=�=�( ������:��v�>A=T*;��V�B���d=� ��6��Xa����<����w�ƺ:�<���Qu=���lq�$��=Cx��?�
���d����M�=3>��r=卑<�Zj=Y6%;v�<�'�e�fZ=�5���ۼ��V��,c;��<�B=e
7���C��|��GH�<Ջ4�["='��<EW��i��=/i(��t =��V��ۖ�Ҿ��C-��ϻ�t�]%E=3�L=;XU=W�c<�+=(X�;���<�{<1����P=�K=T�=�ӓ��YF<�/<�o;�e!��_:<7I�<�,�<r�N����0}��� >k�ƥ�<b붻��i<��!=�86<=J��k�r;%�u=:.�4>���V=�mJ�c�/<�ϣ�+GN=�kH=؆��� �|���\2.��*��[<еM�	�=�����$�U"<�J��4��øU=���<���<s2%=�[f<uD��=5Fv��,A�۞��G[�y��<�p�z�<���:`�0��fw��NL��%�<�$=�&���NA=n����U�<-���}RD=�Uɼ�q�9%x�Q���fB=]f}���#<n���c�J=�����2���i=�J���n=���<߆��
����;�"`=}m=ys���0U=�7=}H#=9�l��<=M,7���<'�T<~���A<�b@�\wüG�T�;��;���<�:��X=Ua��O~= �'=��K=��=!c:<3��`�<��<>�0�d�[�ѼИ\=�f=�5���(�.=�R��(���B=������<2@=�=���͈$<^�o�k�<��>�W��d5<�����fB=;#;�3�^=�wW=$�����<b@���Hj=���:_�.��l��y`n�=�$=�G�K^?�!�<Q�<�ħ�]b༲�0<�K���#�H
p;Wj'�H��<"�0�D����%=qFy=�"OW=�����m�<� ����1�N;�<��߼m�E=��"�
�>�H�#���f��B5;`�;�2\��)A=<X��$���.�?��툽�t��[��(���W<��E=~#�w`���E�ϧp=��X=��I�\���_�<�[=-л��B=8�=��K=/+
�/�=�0b=n]`�@�Y�w�X=����}���c<,��C�S=�$�;�@� M=O������<�Y=m �����a���1��6=��%�|�0=ͻ�2ü�Q==x�k=�9I�d<��=�@�d���%=��<gz�<bIT<(� �	��;w�<H�����<ܪ@��N&=]4<{L2=�м�f��R�<�l=���I=�8��=��}��z�;��t���̼U3��n\��*����:��<��<�X;�y# ;��ǻ\�d<͔3<_��<KΕ�E��<��!���1?�Hm���
��=G9e��e�<�w���� 9��O=gw=?W3�w,=�)��_F���/���	=����<=�Y���=�΍<��<����5�<�P�<x�<x�=�g<��D=�J��g	,=��k�^.���pO=N�;�{~��@	�:;z�[=�����0������y;Gx:=[l�<�%z�e�6=I:��ۼ�;63H=x�L��
=�=���!w#�`���}����<GMC=9p1��D=Wn�<d}�~D@=���[��<�b���?��'%��'<sdܻr!�j�9%���bT����Ft�<z�#=�f <��=������N�g=���Մ=;o��Hz<���m�=�qk�M�ɼ��<0�G���]��T�p������	= �6�
*��5�C�0��;kQ�<��ͼ8�<�{�<��<(m=T	<�w�kSE��"��	(=�q�<F�%��W�:Le���z�<0�(=����I=R)���;*�<W��<��Y���@��Vݹ��;Ѱ�ib����ú���<�f����ݼn�<�;2�Γ�����<��N���;T�%��xv����V���=��p�B<A`�;����sFq��yc�Z�y��k�<�2B���a<�R =ʹ<�����Ǽ�f�<������/�+��8�<EFG<\u"=}0��c�㼺<j�����.�<Xޅ=��o�iݾ;�H�<u,�,�L=�ً��f ��3�!��<��0=ީ-=Go��IV=�������<8�����=p��[
���ɂ�x^^�^�N=��8=�=H�q��w�ĭ�<3�˹�g=��(=f�9_�<��4:OG=N���Q���`�W�=\�0���X<F�'='����K =���C��ǭ�zʸ�x���[O�䡺*�>;_=t|�<;��=���:����5=�^��c�;(��p-�����0p5��h����;�.<�>0=��I=�	<ĵV=t�=\Ư<��B=W�=��<!,<�J2=��:�BX���q��Щ�[�<�VT=�/[�{
�<v<4=���i�<�Ç=����A��;+��=�3=�?+<��s�|�<=���=z�_�J�߼�><cJ���6�<��:=�����a��jY=<*�����e?�3,��(=}�z�h<�,p��Ն� �2���-�
�=� Z<}78���<�o@��k�������ļ]P'<$�R<��3ĻmD��z=0yM���0<#$y���B=:t��?1<���܃W=:��Q'���^�<{� <y"�J���� ��+���iռV};@$�;��	��D��6��;U����5��X�Bӻ(��Tj=�9�<a�/=�)v������Ի�:=~�g�4�=�!c=Gqj��%���<"IV����;�.f=0��* <���;,s��>�1���bW�:#X�6�&��g��wy�
3�mͼH��<f�?�x6D��>�<��1<e	�<S<�"Ƽ�]��\`�:>z��U�<��A�˵m��w�:%��]4�K< ���f������'&<M�D=Ŭb���`�{�A=��C��9�<F<�Jh7=��{<���<Z~@��.=Ŋ��-� ���<��H�?��p=���<4Ɏ�!'?=�G =��=��f=1aE=ޙ�CE��Tr=<6<���<y�=�����=.��=^K�S�$��@��;�T+���i=�f����G+3����f�a�NW�<�_<�	���=O�R=ml�<�-&�E�S�!�<ݹA=���<?�=Je�L���w��}��3<� ���Q=������<�[�y�B�El��.��������~�|=D�@=a
=�l�� �<8%=p�N�=�;=Q:�=&�-=~�M={TU=6��4��<�@�<��"i=p��A��;�%�<�1<��<�`�&��Tu2��n<�T�;bܼ��n<˓t=H~��~��e#E=��E<Bl꼐e�;�=o���,�=�ڻ=�h��N�<|�<�n<fZ���!�c�Z�1=��<j�}=���<zZ=zJH��(=�d�<%�=����n,=��<�j=Ѽ={a����X���3���B��u�<ɟ���:�<}S�j��<[��>C:o2�<Q��<cj�o�ƻ����Z�Zu�	9�<ټh��;}�Z=��!��J�e/S<}^=o�<>D�T=﹦<"�r���������f=��<4=��;=�\M���+�7�e�qV=f���=�&=��H��}�<�����G=�b*��ኽ,�@��=1\<�S�=C����X�H��<���0�꼒A�<��=��꼙����;�r-����:��=�P�<�J��ߵ)=�u���*=*�>:j�r�e��<V����q��,=�켎sR=
J=d(<=�3�:���<Ѱ!=�,���ŀ�
\=�o�=h����h��A��<��j=�w=;�<$G=�������<5�o;������ĺl����<ӓ\���%�ZT�=�O<ā=�?����Y���Q=�O��<=��L<M�`=ޜ8<�D���=x⼟!�;-!����<'��<@ͥ��5p�VE!�ڹ �+2Ｉ�=
��<yQH<Q����;�+)�l�3����;�Ċ���x=�PٺQ=�!=���<ŭ�;�ڼ�3��l����	=�(�;��p���u=����W�м��<F�A=0)=�X=�g<͍T=\E =;H��Ў3���7�=a�<!�E�6v�<U�S=�к:������r�ZV=R	=��	��Gm�y�ռok����=dJ$�\�Լv��<�'ӻj��t
Q���X����<�cm<������;CĞ<Z�"���мBw�<����'\�z��8?i�<U��<I�q�� ��t[�_�/���;��;g�<�<� �9���)��#�<��K � �=,����Y=��ܼ��<w2μX!C=�]M="����-0�W����:��W6<���+�����Ϲ�\ =^5��E�=��R=?�»���R��=�Rs��C	=��;�%D�g�m=]�=��,=��<qRK=�M��w�ҼaO�V��<ȁ'=��0:��=���<�b��߼S=Uv��:x�7>�<#G=��B;��`�I�N=��;l�j�wd���T�<�2G=+�L���%���I;8)��O4��fYG=Em�;�[��/^����<�'Q<qμ�{��()�"���@���ӼLA�\g'=��;=�=���ټ��"�F2=�Ɯ�:���L;f��W2�;J�Ǽ��b�K��=8���&�=)�'�~�ͼI�>��k=8��<܁���H��j�e�i��<��s<��;��N;C�[=�j=M	=ɣ�:�Z����=>~>=g�<��<u`#�Y[L;���;���=�]=�zB=B9��-�p.��2�;S5 �n\��&�˼�ݮ��=�����i�9��"��� `��}=��@�P���m�U=ˇ�<��<SB=]'[=�ա;���Hx=�.C�� �m�<P�C��&=w�����A��	J;Jt �A�>=������3��]?=O���yhC����R|�<�3= =��;*�l=�R=Y�?=ك=C�#=�1Ѽ���<���0�A���c;����;%���S�<�;���]�v�{����<���;ܵ@�?S�����z1�����"�"�������V�SF�<��<o$��u�<,�k�\�1��G�="�%<��=]*=��a�~����E��n@=)��<-�!��Й�y[�H�:k��Ոi��+���=�|�<o48=��6������ռFj:=Aև�b=?�����|<��6�/ V=JBn��n꼜����ӟ���)�}��;�Q=L@=��<76����g���<1����	���=�:��T�<J4)=��%�<;7�=:[��ξ6<���{:<������|����C�0<]ԃ<�=�?�<�ym�O-==vq�<�40=�E�MA3���6=�x/�V�Q;��(;�J=��= =�ߨ<��ӻ����J%��V����S;��W�hK�g�=�s.=���<�vX���,������a5�_�$��a�=��'=�3I���=���:��<��9�fH��N�h�L=��=��M��lh=��;F�R`)�D���=`�J=�҄���?=2g �%/*�e�A��N��s�����<*n��W�7��`5�<U��s=d4��G[�;�����a[<�2�P$`��=EoD�gI
���<���<�n���=Q�&�)�~vB���d��\-=Xr=Bw�;�VF=�Fq�E��=xL�
h_�j�}p�;@a�<�x�<�a�<Yv�e}�(������<"�*=Nԉ<C�I��W�<���<T$�H�U��;�4�o��,Y=��=A���uw��2�<h[�=|�t=@!I�H��"A=f�D���+�4�c���W=&��E�b��� �R��f���LD�<�c=�N���N �m̼�Ӽz���7D.=J��=Z =Ͷ��2[�D��6Q����Լ}d�#�`=q�ͼ���Qe0=���;7�;	�8��a��,�@�=Fݼ�'E�a������ꭼ'CB=��<��Ѽ^�;=FL<��2��=5=���<8�I=��L<$�	=Ϳ;=��<����ؼ�<�;��<�2Y=lّ<��M��=��YT�� <\=�;^�V<�[�Icz��Lg=Y�J�0^v<>��;[�N=��4=�7��U*=/�;>^a����=:d�D���aC=tV�|��:e�<ة@<��b��DN��1F�Er�<��=Q�ݼ�R��Jƻ�<�~�=O�=Q3M=h7缵�⼚ J:IC�<b�=iP��.��<o_9�к���K�.�E�:�p03=a*=��f�JW;���>��1X�L�-�N�<��=Pt�<zr=��<�g=%��H����%�NG0�ʰ�<[�:�ӻ<���@<{�R�OE���$i;#��'�����	�e8=@�8=S�y��Si<X�'��;��+u=b��@<���<#��<���<�:k)<���<h�w=�?�<9�=�;W�=F�w�t[T�*�3�����0=�ۼ"�Z=/����&�t�-�*Pb=���<��-��M�^4	=���<�=W`2�U�&=�-����Z=�N��V=Ri����<;�;�+�R�=e9������"=��?3�Q_=zsQ�����μ�HH=U=.�"��6�E{��=�Z�:yp_<L8�����g'*��pd<$��<t�<�"ϼ�<uy�<W�����9<j=��l�<��+��]�<8���Ś�;'T=#+R���M�W=��==�=~�)=�	�<[�]�8rb�G�=r$*�d (���;,��<hj�<kT=b��<�\�<� <ݕ0��	�<ے==��-�B ü�q�<w�>����|�<w�W��n�<�A��;�<�3�=����{l����¼]J="��<$�M�mS=�n�vO<�	���e��:\�ˤ߼���<��<2�=���<9�B��;2��=����꽻1Vk�
�C���B=�t}<��>���w)=z��@�Ӗ��aD<~�;��%�"��<�o���; �=������͹A����<�fE���=a��P~�<ƛ���H<bb�<��S=˅6��/,=�p#�ɥ��rI==� I�KX
��+�fSc=e����Z#=���C_���:z���;8�C��3<��;�KI���ӼW��;9�Y�^��<�: \=��<K4�<d=m���A<]�����<��=ǳ=H�Z=Q�<��+:�=�5��]<��Z��	v<��ȼ�'=q�X<[�����漩��$�)g=�f�<q��:)���U<#6=һ�	��<�b�<)*���?�Lv�<�1��\��ksW�8.��-a��w��*��(v=�U�<A8��''�L�=1t|<�%_=���<x���Ŧ�8��;��=�Q�<�>M=$>�;p��<��h��HW=2N������>�;�*�h�;b�=��<(:\=���� ���<�Yݼ�~��S���;'���.=�=]<fϮ��Υ<��K<�)=���<Z�<odƼ<��<Ś�;ǅ�<E�@��`���F=����8K���9�Z<��j����<�c(=�6�.��X=,�<`m<����p⼩Q�<	���W��b�&;z���G=6U:=��\�B�9<iO=�bK�ِ�<"��=�Dp=�7N�q=��k<���"w���߼U�0�! ����<%@W=8qi�9��<MwP����I��:������<>�=���<�)?�曼�>%���������γ�<��=mBE�E�E��A���%&=�<I=U�g��sѼ�E<��=�ٿ��H�<b�<�$D=c�����Ż��i�����~z��e=�d��2�<�ׂ�a��355= y�Y�=�0�l@=W�μ�B=Z[J<`���$`<l&���k�<C=֓C=��"<|k@=Y�<�(=G�\=�40;��1�
����!�<�=��<g�W�Wq�<�+;�@!��<v�U��[=�E=*�ػ�'�c��P�"=C�� 6E=�u<��#�g�b���k��^':���;����o�z��!R���9=��b��i�u���ļH���%N���ѻ$xY=���;R�$=q�кSr<j�<k=�c�<�,�hp4�I���Ea��h � 6I=����f�=��8�#�b����<�7<�̳<�=��˻��`<����u�=D!<�]={��:�s�<�a=x*���< �Q�	��<�j.=�(P��f�SN=�����߼{ ��ċ��ۍ�<�O��md=sν;~�e<!'=��=:�ֻ��=�$����(=i$���]=�N�<<�ȼ�>L�1�@��Ǽpv1�M{�<�U�v�Ǽ2@=g�=̷�Ҩ==1$�<P�g=+*V=��:\d�<<����`�<�x8��<[P���00<��D<�?>�v븼��*<�;�:7��A���<��Ӽ�*=���;/c_���<�*�H=�I~=�,ǻ��:LK�����~74=Xr=:�<4`o���q=P�;j6���<bF%;+�Ѽ�(����<=I�U�B�-="H��6!<���Ԟ�<�S��oJ=x�y��J��n�s =�-x�^�%=U5�?��;aK�<NF =��;K�=�\=��P��!=���<��</=pFK=R�S=Z�D<����z�L==W�����%�޼3,��^=�p�<�<�ɺ�F=��=��;���<�(=�RB=�U���r=dFE�M�<V"=�wU��z[��e�!�P��}�<6O2<�86=ƪG��Rڼ0}�}P�b�޺�D_=8��;�*���]=��<��a�ꌈ<_)Լ�$E=F =o�~<�.��:<�eѻ�e�:��:;bu6=���<�I��_=3ve=�Ⲽ{��x�<�����n�f�=Y�<N/��8=��J��`L���<E�==Hxĺ�:=>�K=T�?���p<�P�<�mD=�����׼Tf�U<=}X���Ľ�Q0�퐼�3=Dݍ<j\D=<�5=#9<J[y=1*��d�<��<���
<��8�j<W� =s{���<d=}����<䵒;��=�<�%	;��'�v�D�c/~��� �~N��.�'����[�mIC�9 E�f���T��ڸC=o�<�,�=Z���v��� =]#?=i��	�R<�<Mժ;13�<��i�K�=L�<�h񻔒�C	=j�Ge+<W�*=Xj��M/��9���e�=�G��V�T��;��<
S_�܅�;��'�[��<�i�<��y�fP=����� :��R<�^ɼ��'=u�<, �</
G=�򍼮�<qgI=���C9'<W �<��_���2=ͳ_=�|.���\<��5�?=���e	�Χ����'=�*ԺU=��dg<I��=O��=`�<�V��6;YU!=J+��=�=o��[�d0=@�<�u0=K)�<.]�_�]=�\���1�4����NV:��:U���;�;Zth��\׼� -=���
@�9�X=O�X=��E=A�l=�Fh�DP�:�/��:1;����
S�N֩<���<4n"=pG���ē�a�S<
�=оH=�6N<�=��.�11=F�=�z�;�"G=Q
c�4V����=ڼo�X"��z�;�.1��H7��S=~6Z<��ݻ����{<�;:��<�c���<k1%=E��Bo[=�.q�H��<���<ژ}�mJ;��I��Ue���b�\�Z=�J�:igV=>M�yCW�em<O4<��<ed%��#�<&�lh+���K<��%=u.��{=�$�<�2�<�/�g��<��<��=� �5�t�
��^�)��K�BL弯��;7?<�F���4�<P��<di��M�C<Y�;ѷH�#�9X�����+=��^=��h<Te(=�P?;�G �|������<q�<�ˡ�,�������>�<�?h<ᢺܱ�<չ=��|=���;C|�<�����=*�<�b�;�9=c�;���L��՜�Ǵ1=<��-u=�o�<L~r�|�L%��
y���� ��H���l=��w���Z�^��	��T�ܻ�|=���:.=�������ݘ��;0��j���e��fU���w�̢�=���Y1���<�*W=9n�<��9�u�{=)X>=��f=����z=%�$=R�<w���o��u�< 	=�<�눼FJ�</(�w�D��M�<2$+=z<��'=�uo���?=�f|�r��e?P=�R�=�]��<��)&ƺ�\=�#��9Dp��J<���<��b���=jp0=�az���|<9�3=�BA�E��Qd<k�����ѻ�<�F�W�<z�,=
H�L����7<�B��rT<*����{3=�/)=ȡ�<�ǫ<���"�Ș=F��:�	=G�^<Ղ��<��I=$�F�g=�6x=-a=ɟ=V>X���U<ܿ�y��<Bߤ���)�G�
��W=2�E<B���Y[��F�<�DY��}�)hּԿ�h"c�7�<�<�����10?���.��LF�i>����<vr�$��;��|=�`<��l���=R�==fl��%�o1=&h���=��*��h1�<�`='آ<�9ļ� ��V�5�,�p=��O;M�L=�<|&ۼ5���,=�T
��p<���  �;@�e<�#��X�<g�
��{=��7;"�G�m8&=�2G=�F=愼��!�N]%����<�|<4A�89���4J=����FO=/%<I=5�*=s�A���%�=��_�s�<�$=�y�<,�����<�w�<�#J�6.^=(G2��p)�d�M���6��|)<�p'=(�;%���x`'=1��v%@�R�9=��H=���I�����9;lk�2�c=z;8= M���V���+J���?==b���SH�:E��N�<̶<��]=��9D.����b��/Y���W�{3<��K��!�9SѰ<�O)��]��/�R��<y-ռf!=��~�%s=S��<m�=��Չ�����+�KI�<g�<"��<�Yu�&�D=Wc<�����;�c=�6���+����N��U�<N.2=��M�Q��<J\�<wz=�{�;~l�~�.���<E��<{Ǥ<��<>
c����<��M�O�[�u|���Q���'=ҠH�D�=��B�zs����;!�=/�Ӽ�4H<^{�<::��˰��� ��?�}t"=>�U=@:E���T=��=I�e;b#�(����2=�^�XSv=�p�q�<�/=��=�i�R=7��v�n<v�:0d+<��#�*�A<�b}=\V����c;E��;���<���
\�;Ψ�<κ�� YP=����	�/�h�c�m=CH"�	(`��ü�@m�E��;ʼ�=S����ޢ��XGy<(��ޣ=\A��M���C=Q�j< E�<cJ=�w7���!=?�<I2�=P&�o�
=���M];�/<M��<��i� ė��3 ��󅽙�e�>r��H	�<��=`�|�޴=�<ߺk=�A>=�1�mH=�iV��7=}bz<I�]��2����Ƽ-�V�L�<\X=���0IV<W8�<8%+=c^�A��b��<3�j<�r��}�����-�D-=M̱�ղ�<*B��	����}=��
<:%�<3�O:�����=A@��/=���V3O�q��;>}������R�=<fz�<�u��/:<c¦��Y뼥ܵ<s4=�U��~�G=XTQ=2�z�.�6<�R���>%=��5=��;s>�;�g�̀�<=ث@��4u�e\1=��;_����W��3A=��0=�R�<�hX�A�˻u=����ir`����:*m,<#�񼞵e<�"=��=,R��ɀ��;�:�<���<�ڣ=9G��9��=6���b:�3��,�%=t;H�B����&��
�QZ= ;����e�;:6=��#=I3=k��t��=�`i�Q�h=�V�<4*'<%�<8Hʼ���;S�0�����'[=
����9=�����=	���=t� <�IY=�5��\�;��뼴�=0���oL�<l�-��n=���U)<�5O��%�	�Z<~^�<�Zp��_�<�W=�Q��t�v;��!=Uͻ)O=e�-���<� ��Dr=2g��Rּ�̜<9E���;۝g��B=� =��L�1μ�r0��%�>I=�3='a�ȅ�<߼��V=��<{F�<17W=sA�<_�;�=���h/�� @�)�A=�U=&��듇��R�t�7��s<P��<�㏼'PX�F��F<�0q�q���ͼq�<�����W=L�߼4C�<��F����!���=���:X�=pz���^C=��Ż!⇼�5+=i}O;�3O�Su��Gm=Z%=�z=^Z�eh�=�qV<:F����1=�m켳�B=@�"�+��C��<0����>���;�W���@�s��= ���d�և�<^��;&o=�%X=V[�<{<�B�n'��\���p=S/w�D��;�\=��"=���<�И�
=.rn�}�<�=��/:<r"��3ƙ��A���=C�ϼ+u=4�9ю���R�`��+$�
]���K=��Ѽ2���K�<��8=�a@=G�&�r&=E丼\7�{�2���<���=CԚ�z�=�żH�J���A����@�1�'=��һ��(�<1d�f�=��>Ry<�6��+��<r:=����	c/�Ij;��D	=j��Bv����[='X�h� ���`�+;L�C{X��+Q�_m��gv!=D�=c]j�+��4�0�]Mr�c�=Yt�4v�:�a,=$=�Hg�w�<�<"*1=��!��H<����#��q�<�%@=�r��ƈo=Z�<#(��Q.��~R�X�H�;I��!x�������<Ci7=t�ڼw�<��"���Q������׼7X�^����k����j�m�r����4�:��=���;SF���<!jc=d�X'<��^<ӄ��l�=��=��7=<�=�ep<�ԩ;�)����e=�� =��%<l��<#o�;���=Y�c��+=勢�9�o<|\=���< �=��A=k����UJ�f�.�+$�&ܯ<G�-=ZL ��MD=$ /�O�)=N�;p-O=��w�����p#=�E�8_<��1�8������?�<�$=}t��8`_=z���L�<�z��H�]M�<Na�;1�>��E=�H�;W�-�5=�m�;��;dj=�=x2=1�=�~��tz��I���@�/�R=m|��Y}�W$;JD
=�b@����]�����(�z�K=�9,=ˡ=ߩ_��-��^A�<�g=��_=*|�f�<Z���O�;'��<U�S�Ov�<��~=Yd�u��<�<�B��Jp<@Z
��#м�`ü`�=Q�<�g�<�0��9�A<����Y켥%z=�>< �><��O����;����n�}/Ƽ�z��F�=�,�=�����= IZ;�{e��Ԉ:V�h=�ɯ<����h�޼�\&=A��<.�6�b�3����<1k:����J��V(���?<��=�=vU�=W���<������;=n?�.d�;�n6;�56=��4�n�k=���:	7=f�мbH�� �B=�rH��`3�L�r=7�x��Am�j!t<�Y=m��<�U� =xhż��E=���;������;�"�;H<���<�wݼ���7�c�Z� Ȟ�fx<C�R=�A=v���@����<�FN�R�;��0�>D=�!�<p��E���_��=��<�켼�z�<Y�<S�1�G�!�[A@=
n_���P�rj��� =�=[R:�C����P�{�_�	= ښ<	j?=��f=���<��9��=���%�:�^�c"=��?��7}=�?�=�D�6Յ<����g�<e�S��ԋ<�{0=�쇼R:�z�,�\jH<5	|=�)���,�(=r�Z�i~��ik�:GH�$==3�<1��<�!=X-&�:�<]:6=�0�<9���+�=���;���<�; ��9Q�ܓI=/�����<P!���?<�]=e�<�����ͦ;��\=G<��F��<NI@��0=������;��d�d�m����:��\���ؼ'��&W5���<��ȼ=.p�]���Ր�8�5�=������B=�P��%��?�<��8<��6=�8=KC=�j�;��H=����r�<��<<�48�$�[<&
?��w��c9�=�Mr�n�a��Q�<�,��4�:v�I=+��:!	7=���<(�̼�#����H���=���V����@<�z(=sT�<���<�mH�Y�=�ּ�`�<���j6ؼ� �� ��L=^0b=��'�P�'wk<�_p�kЭ<��9\���&,�<���Ps�<K��K[��TC� 85�q�=� ;{��<�cq�tIC��9#���9Z�����=��*��8C�5�2��,=F̆<XI��c�k�q?��N�����:�y[=XP=�%��MD=Q�ļT��<��X�g'���(A=�?���ŻU#���Z=��򅏻�򋼟�"��aw<��ܼI. ��@<Z�;3M�S�<	��:��=梹;d|ۼ@���c=nw6=�`:8�ȼɗ��GN����<��I=��f=��=oqT=��;Nq�����c0=�� =�󭼬W�<���_�)<o��<_��T5�<�X����0�g��<�J5����<�!��¥-=X,�塄�K
�<%nP=�eI<1o�<�J2�!��<��=�p�<�<��4�,�c��'
i��c==%�L=o=�a�<����E׼���<k��a��� ļ�o�]=�$u��s)n�(�]=e���	ʼ$?� ���E=Iu;�2Ҽ�N=c<.�C=F��;�j=��H�+=О;�h�<L4�n����!=��O=VC<�ʟ�<��k���"�W���}g�?���`u=�t ;��?=�/��k�d�3���	h��z��&A��4׼s/�<�_�5+G�r��<)i'<i�;������=9���`�2�<=��}����"�<N�<���;�u��ZtA�${/=��n�*&=��0�|���ט������?�<~�g�E<�<�al��̯�P�9=�V(������ng� #d���;��7=$�K���V��%=��=&ee=F��<�<�<�X���]=�fY��	\<*���10L=��]<���<����<�r.=�8�/"�<�W@<��C����=�[g�FX=V�G<;9=a5=���<B����U=-!�;�^\<C�V���=w _��aɼ�)j�)A]��T���/]<¤�<��9=��C<���<��Y=8k�<�W3����<��#��7���;����6��<dr<�t=�6�;��l=��`=:D3=�\�AH=���üM1�
ƍ�lR�";��s6E�U<H�_�A=ڠ�����:��<���>N��H��v޻�FU��e�<�"���=�H�^g��=��F�/�<�`��n��.��~y�;m,߼�� ]-�M<W�G�߼$�)=��/�Ӽ�(���|Ҽ�@5�'�,��=�%H<x"�:c���f����<�%=Z1`<[*�U���N��=諸��*<�O�f=B>�<[��;�;w<�1
<���'�U��u�h�M�<�s����_�M=R���PeH�dg���fM�>�<b�`=���;R7��<T=�=��7=�����$��W�:�#=�|<�	+=	,=��0�����'=�J<#Lg��f��h'<�`��ch`�9�
��Ok=v=��T<� =G�F���;� F������`<�<NPb<�>=�'K�����d׺�C*= L=YE=�Y��*�t]3�w�����;
 <�B3�y�E=*�X=�� ���L�[���K���ƠW�q�6����
=t��<��j=s-;�kʼɁ�VLr<��X=:v
=K'�滷;3U@��M�$<99=�~�����<|~=�Z>�<h$�<�E=�!���R�_�;5�����~�;�=���<uc��=l�4�C={�X�N7�<�=&@C="=�ゼ�v�(��<��:� �<�q��P[]=TCs=��1;�=��=�]��v�h��<)8+=X�="���T#�+1�:m5G=Y�<��1H=`G��%�=&<��5�����Lͺ��8`����+�Ӿ��d<���
<N0�;��;=���;� ����+�N��wn���N <�=
=�I<�US���A=���<=-�<=NCX��G=#e�����<�	,=�,\<�{�;��7<ꔥ�Ԍ��W|�<���PtY=��˼�K=_�8�ز�|�=�x���=���*�j?g=�h =��<���;a�I�鼫�����<���9����7���˪��W���߼�h�i��e"�<�Ղ�����<�x�>�m40��
�<�@�=)�d=��3=4�Ƽ���<A��h��<�3�<P(�<����/=��Z��"�<U�%�h^=��ü�m��S��I/=;bs�<R=���b��qC�KI�;϶��4�<���=06�<ig*="���_��9��<7[����;p,U=4򨻉Y�<�{=P�=6}:`*3�y�Լ�+H=s.���v=�~=tu<���9�X=�Cg��#�%�����T�T=��<�@���A�Sҋ�x����N�_�=�����R��d#=9�p��xB<z���r�941= ��<��=�)%=-Q<�ͦ<�D =�t<d�X����·�{�{���=D�=df���^�8�=;:��<z��<h=)=W��6��<��J<��==��P��-��+���!�0Dr=��u��c�<d�i�k�o�^t���&��Y'=~L=Ԙ8;Sd�X�b�y��]/���`=e�<n[<�'�C��<�K�����OUj�~�{<��#�*�=L�ؼ�4�9&�C�hh�<dߝ<�<�V���(�����`�Fl��;��(��f�-h
���A��J����=	-=�~�:���_A9�~�;V�D��+H��K=<�e����<����S��<�=��R����:�a��]S=$�/=�,~=�;�����S=��u��A�<��<D�8�T��<�df��)'�I8O��&=_��Z��<�	��������pq<7ͼ���<�
==�;=��&���g�<,x�sn<�<�o��>=�_5=r�=;�M<[>�N�<�"=x;b<R{��������<�)=��E���(=TOj=�N�<�~V=����$=���<��0=bJ�<����ּ&Me;��=���;>"�Ȍy=�r�<��r< \��n���ze=��1=?���A�"��;�㜼�QI�E�켹�j���b=q�y=@'���ͼKPs�x��;�&$=L���O#=w�<��>��I�ut�+H�;�<܀���S<h=��=��b=u?=�����y��`��y(����,<E� �G�<;��N� ns��Y=j����˼C�Q��_���ǘ�iv��	.=nu�:%ڼ%������s,��Y�<���<�����<�D����%������U�<��3��"��?������D�g��<�ȼqֻ�s���k���ᖻ:]��s��El<$V<��0=B�{<m�3���`=8�d� �B�r~<�Ύ�M��<4�6��)ؼ�T)�(A�Ll�<`�M�]�s���=��B���작�K��<�/`=U?�����]�<'��<Æ0=�li�1�`<�J�� ��<��?���U�[�W�=�Ⱥ�8M����<X'<�.�K߲���\�
{I=����=t���<Xiw�f�<�VT�u7=�Е<�$�-Eμ@ß<�7b����pL�̙���<��¼���;|���9=��=W������������9�M�|�!� �Pr�aBk=6���'=�u5�_������<�m��G�=F�O=t.9�	�&�֩��H������;j�/�T,<@�ܼ4��<�,�<��g<S��<��˼��J<�<�� ��k=�_\;�WY�N�N���*��a�;ܪ7=��<e�=���<�	�C��<�^�<�S���S�ޢ<>��g�<��4�s�g��2<�Җ���E�$b���� �p�R=K�)��{�xV=�=����?��/=���Z�P�'�XH =>�1��tI<C�<N ��<�;,�ڹ8�_=n�O��U�9�[<[<~=4�=�0=b�v=	�=�Fm=�fl����"��<t<�<[Y���b�<K��˕<�O7���~�bN=-�	��d,=�1�#d:�j$�V]-=�CR��&~=�����Ϻ<nO=X�A=jo�<2!�e���{�)�@�� ;��y���v湮�W=�z��2'��c+����;v���<�<r;��_=��w�m�<��5;X�����n<�2O=~�O<��	»:�V�<�J��H�<�/k;
�ٻ9kB=*�2=�QD� Ƌ����<��:hu=W��/��%�=�ݹ<-�<P�(���<j�&�R�=\R=e"�P���M�
��@��<�m���-�Dm7="�N=
�g�+�mS���=��;D?L�>P��6=��=k��ycg�0�x=�:4=�$��ʯ��w��!'i�;����*6����(�s�<_#�<�k<�����7���~(��zC���ڻ���<��<jά��d<?T=d����S=�
�Y�;<lU�N=���!=��f~���<K��	����6�z<d=pI��x�<�R�@�@���7�$=���OK@<��_���0�]�n<� ��<�h<JQ%�!�(=�h���=���9�W��=�Y���s<��M�'�u�A=YQ�;O���sA��q�;�Z�loüq��	�;�'ۼ<���!�F��ſ��n�|����K������<�H ���`=�P�<xق=l��O�	=�_Z=e2�<Ԋ�;��L��/պ��X92��o�<L�=�@�<6�;���<ь<I�<O��<M�=a�<<Ì<Q�/�v�[=K�N=W̎�sQ��`h�T0��Ή<3Sf�A.=�c�x���I}W���=%�r<6�=��<zA4=c/=:#�>�<j�=^H�<p��;͌�'h�;��<6���]m�:�f�\s���(J�o��''C=Z=<�	�Z�+=�0��ђ�;� ��n6"=�[�<G�5�h-<麼;[���;�
��ʹ<'U���<�[��}T��xO�e��:4?��@��<{1��/�;+gP=]:=�Ҽ�y�<�p=uς��R =����ju���6=�D�<5F=�����<Ϳ����c�Ih=�=���;��"��&���D��OӼ�z;���h��je<�ę�.�����mB�;��z��ֿ�pt�ťk<���;D#���;�'7;�Z=��&=��b���<a��<��D=O���;�`ݼ�����@����!�`=N=Cnd��O$�� �;�E<=(�<i�=А�;=���q�<���<w�4<���<�%�<j*J��<=��<+�.�5x=WU��]�<S�+=f�=�,=ۻ=�c<=tXW�_���M'==%Z�U���/�<�u�<��=[^��Q�����N<CX�;�=�u�<ī�������'=�b=WuA=��Z��'�<�&ǼU���e>-�-�������h�O=Bz<�vTz�pAY����<Q�>���=n�}=Ʈ�;�,=����3_E=�0"�d}m��,j=%���E�4%�<��:�h���C@�+_�@�P=��+;"u�<��#��0=3�(=R]�;�E�<B��r>�<F֛;�PF�����/�l�<��3�ѽt=3W�g��<z��c��<�s:=��<DrZ=�ұ�OӅ<_<���� ���B-r=�����PH�;�K= A�<[b��lE='=U����y<i��;@�)���*�=v�z>���=/�j�	=�=h4d�,��hiu���x�\^=�*�<,==E��<�R2����<@����|<�ש�
����I=��/=��b���;4��}��<TL<b��<z���',�@�|�I)j�d|�<_��߱�<m�M<�e��3)�<z/]����<�����<�N�:������=�u�<(�g=V=@��:8l������jw=28r=���kK��2t=r)���=#U˼\�+<o�{��hh<}&�<�2l=�,=���,��6{�<�:N=�{���B��^<	��j{P���<���r!1=��U�S�<�iN���Z�$�w�Pq=k!*���< =��ػ�J�jGb=]���K=�jD=x���a�%i:�����g���'����T��x�<�`�{1��K�/�2v<^X�<�9�<��̼��!������<I�M=LE,=��	=$�;l��<2�Ѽ��%=:��<��G��<��<��9�z���@sp=J����K��}�<���B�<�v��č=�*S=�$_�ќ�<�2ټ�����u;��<j�Ҽ~��<?v<��^����b0���x���H�<�W��ۻ�l�ī�<E���qp����<mˋ<�=�-���8�<?^H�n%'=�G�.ϔ<�%=\>C��~����v=@�M����)��#9#=fR=_t;./m=������Q=R�[=�ȃ;]��-Z�i�<Bڊ<-t<�O�WQ*=��)��d�;N=c�;F!#=R�<\Y�<�J���B=�J(��d���ѹ5���q��o��;�1=p�=��L��Hg�n�,:�r鼑�U��:?�t,ʼU���=�[��R#��W[�<��f��U��gp�#>=�$�<�-	=��F��.�<��t����ҷ�<u�=���<��4=�_=���;u���?�<�]��ս�<��<�d<������=����4�;"+ɼ=�<��<���<[�L=�p��c`1���=.8�?��C��:��;2Y�<tĨ��s��ʧ+��? =��W=��Y��.��D=���<@Fu�Dｻ�*Z=�k�;��d�=���(0�<L��d<^,W��3;}���vջ'9�R,ͼYD���-=�y<	��<�5��g=.��<�F
<�k��툻D�$�D�=�;��<j��ݼF��<뺘<�Z�=��ع]r=�c�;{��m��;�<�����<;�=XU&=:������:�j<�w�<=;����K\=��;*8���<�(�;M<�cּ��@=�a;��	�=�C�<r�J<�J�ѡ<����鹼��<��<~}ѻq9ۼ�6J�q�����L��$�*=@ߖ��׻�s9=i��<7h'<X���G�e��s/=atr�`#j=Ou���;=uռ��;��>��� j=鶍�������>=[���#<=��5=�=KD�<40<�g<o���z��;��<o�"��W#<��f<��=l�l=,������G�9=��!��pӼ�j3:S/��j��ۗ;�xq=�=�x�<Fg��=o�(�nv$=6o��J�<i
�<�N㼑�0�2�D��=p=�ʱ��sa����c������<��<�ҿ�hMżil^=�/W<�b$��L=g�	�9*b��.�����<$ڹ;z����<���;�z�Q�<�5=φ����a��;=�&�Z:�=�~����=r-7���>�Gsp���<MC��$� ~�<�O=�o��0W=�D�� d׼�E�<,�0<ǆ�:��d=��6���D=�f�	6c=�3e���=�d=ut<�]=o�J=����+N<r+=��;8	]<@lg=`m�'R=f|�<X$���3=/Yv��+j:�=�U<������<���=96Z��?<=xbT�㓕=9yx=Rc���R=�8<��@�Ԃ��3<�<���<�]�~U�I�޺��M�ˊ=8���"�<sat���C=$��;̽<0ܸ��M=�@��k=E	=}|໗�@�eII=h5漞ɬ<jV �P)�<ŀ=��=�(�&�<�#�<*���k���,�<�?j�*r������)���ȼ��
��ᬻ�8�<G>�6)]��o����߼�?=ݩ2�~��<z���5������be	�]LT</�D�
�C��ʞ<�%=����OU�<kp�=�W�=yC��S���H�����|�B�;B���W�D=���%џ<OFN�AE��ja6=7�J�i~�<av2�����"��<l%=�� =S�<7Q�<3壼.�?<�z��i'8=e�W=��-=��ü���:�(=Oj>����:˃���=&&K��^Q<�p= �<]�<�G=.\u=�	��I<=Κֺ�)���x�<�m7���=�q:�X2=�d���1*=�,�����|��<����' �ݶ�<�S<z���֢<�za<��q�{�Y�x<�R=5f�9C����ڼ���<��-� 4'=4��<c� �!g뼕yǼ��_<w�M=�Z=�h��׀��f�j���;�=�9=�9�<���<�1κ�B3=���<M[�<m����ɼ�\�Itj;�=��<t�b��y����ؼq����2�<��=]H̼��=�<A�2<9�p����<�耼� p=h~c=�Od;]�i�w> ��b=߃\;6�)���I<���<f�.���<�z=Ju��|ds��`a����ƍ�<_��<>��;��>��l=���;F�;�S�<�C��Q<�#*=q��<Σ=<���Ӄ<�n2=�w�l�F<���<-0����P��,=�u�B�p=�ۈ<��{]=U�K=��<���;�.=�=�����<��{<���<\�+=��=s#h<@�+<ӻ3<T�X�%�U���<�K�b�|;�����뼬~�n����^���(=��:�C��[;�������;[�ͼO���A���k=�'��u�Z2/<��<��:���<��q���=���<)�f<�򗼃�#=#��:T^��ɋ�4O=$)��|���<��`�Ȇ<N�<lJV�\V=��<���<A'	�.$��� f���=�4�6��:%�(�N�˼0t=��V<���<��<��ػHf�N�üCi�yJ�=�3���L�4P3=���<h7=��x=\}��,EK=I�%�X�=&�=�ʑ�M@�����;�@=:���{.=cT��SZ��M#=�4�����r�ۼ	$���=|�!<�e{�0BN<�Y.=D����0:��cv��"<��=�"�f=D7�x�D=$�Z��2ӻ�ɼ;�N�2�Y���v��;=��<y�d<��O����=_�<j�@=�&��xO<AS�W�<�K4�6� =�

="�:ª<M�<�qƼ�7��߉�������a/�<'1=r���P�<�J"<�(�rF���)�n5����h;��9��-�;�S�<�u���F\=SS*<F�=��μ�y@���n=�R=TJ���j��J�<� =�x�<��ż88=���|�r!U�S��
ֿ��AV=s����1�R�=>=[�ɼߝ¼��]�H	���<^���s�<��/G�<��<@���G�G�>=��Ӽ!�P���=k�.��;֭*� �u��r����\�p�;���<��=��Q,x��1%�Մ��Z��.`6=OA8�"�F�i��W-�<qn�<!�<�m=���WL,���i��u=��<�H{���[=��9��,2=u/�5�;4p0=�h�<R���J�=�0o;q���j�ǰ
=�2��xP�5�P�4�=t�o�d5żCg=��1&��#�<]D?=�	�˙��R�S��;�l!�3�=!S=�W<ԅ�<��<���<΢�]QM<��=�<]f��R�<�����<A�=r�j=� �<�Z*=g�ĺ���<�2��=�U�7"�����}��dz����K��;����ywA<�N����G=w��:ŐK�o����<�Q�t���CK�����>[9=�ƞ<bk�9��;��,�v��LT}�����Z�黪d��#�>�'�0��j<��"=��'=G7=�*�+=i�\ z�Iʼ_W�< l=T�����ڼ �g��|?=BY[����<�\�<x@x�ه���b�6��u�=j�G;��=ݍ�<m4n��[�;i5=�!=�v��$
=5�=���<�)��ҳ��0�<��B�ނ�<V'w�{j<[�==%R�<q<�;���<@s@�ļV=�݊�rU=�$�<Ve=���:��]�_<��q��{=uh<�x�<q�={����C�3=��!=�C	<cI��8�T0�<��=�y@��K����jH;���<΍����7;��B=O�:<#�e��z�<�lF=!�<C�������ꝴ<����F�(k"<Ux=�=_��<d�N=!Ҽ,c�H��+�=���V.=��ü^ű;K"=l!�B�-��/�<k�E;�Z����P=~��<YMü���R8;���?e�<���<��<�j�<�p<AW�;?kb=+�=@�!�,?�<��<��ü�����'�<�p==x��a-<=�ŋ=䛘=�<��K=�F��E�i�\=��ֺH&���<��<���;�I�<����ԣ�yp�:ex�;�W#=US��n=�q�<���<{��<�%F�NP=�D=U8��_�P;]��;5�O�~Ɂ�F�漍�
���켾/�< �C=��C���^����,(��I�<0w&=��<!��=�ke��b�<Λ�:Ef=���j5�<9��ï=f�<$?
�F4=�=���<G�I�9[9<�<�<-m�:�2=��[��亿?����5�������<f�?�T\�<��<;�I<��=C����HӼ�"@=���<����Rv� �v=D=��<X��<����_t=�0���\��D����<�<�;2��s-�)w<�C�<���<$��=;=��V��i#��M��
��;�5�<*�=<>��g&6<&�<0$��&=0����߼[��H=8 ;��
�]�0=v�+�t݁��+1�*��<��
=�m#=��ۼ�U�<�>]=k+=k��=��s=����C�<�+.=]��< M�<�]�<T�<�B�0U �ϸ<wT�y�`=,^0<.=��=�0=���{=)�=�9<������x=�(<A�^��=��V{��GQϼgp���p��Ǘ�.�5<ݸ%=�D�%v;�cz��w���H�c�!��Qs��B�<`:@��żO�P<1<�(<�;���Lm5=&��ǀ<�)̼%p��*�"����[=|޼��޼\"�QТ��o����6��c=)P���\�E�e���X={ <=�=d�˼����o $���{�ZV1�O�n��^���a=��0�]f@<l�\=��q���<^�!<��;r*M����D_X�1�Ҽ��=m\�&�<�7�<[8�<$,<0 ���C�<lfȼ��)�U�X���J=:19=������<�l<��༴=4=������;9��~9�<^9�<��A�ֆ@::�^;�)<�1�cC���HE:d��<L?^=;=x��5ܻ`1���P��2�$��c����#��X=��:�⍗=�>���#���b�H���A��1��u�*=��/��,�=)���	����<ʪ�s�l<�������<0�S=���e���T��%(7��(=iP��O��>=n$=U_��#.��;�gO���= �<��<�^<��Q�;�B������#�E��; 1�<����n:���C�U�<��(���=L-4�M"��;��<�U=Yb�ѝ��m�w�<;q��f�9 �s�<�<��\��~<E��:s*=��2=��c=�z=�=D|����<�AZ��j=�]Z='2�<óu=w���C�+<7�<�؃��j���f�sn<w�=��O=��N=�3�*�T=�'^=�=���<����rx�n�M<�?(=��<bZ�<b-�;_1�Cf��y����w�����;���<z�H��s�<��<�3���-Ӽ�=x�뷡<8�n�hPd=6J���N�;�& ;���<�\=~|�h�<ܮ3���1�;�Ǣ��0==�#����)�n+="��=�b�=N�8���P=l���3�z�wdS=�7:���U�Q��:a<�<�z8;����m�<6�j<��ּ�7＿κ=���S��Λ�	��<З@�H�6=��+�q�i�����&�(Q�<G�:�r@;˱¼O���l=7�=���_�#=��d��n׼T�/o=��g��T=F�6�#==�@V���{��� � 7������4I���NӼ�OG�|W�t�,��}5�4�Z=�ѓ<'<v���=�y���<Dx!��Y��\��>�6=l9׼=0>����:%у=߿�<���v%�;b�<��y�wr�<��'=�!�?�v=h�A���G� ;�/��n�4�En\=<�r�������3=�I)=���<E䶼*�<F$�maW���<�)"�ǉ���Oͼ�˺п\=W�<g��<M�<�a*���t8�#6[=q�U=�»}J�=�^�fI�Bdp�8���V�<�<��=���x��=[�)=	җ<�Y� ��;�{��E�E=�4<�	<:C�;��<����<t7=�Lh<)�b�;�����<��}���1=T{<�*F=[hA��y�H�=z2M�;Q=<��:<	���z��<\)��d���Ǽ$���2!J=����>�>=��:��ʼ�6��[G���=�+�����'}=����k�������X=F�N�`�!:�.=CMk=��<!ZO���=h�P�f�g=Q���t���&�]=��#=�A��m�l��`��7;�<܏6=�7=l�l�Xj������v����<�r$;� 
= Nļ�2��E=lIK��x/=kP= k���=1=�3=C"�Q��;W˽�y�����~�~<)�!�m��=�1\<5[a=� A<Z�M=S�e=�Q�K.�:�x̼�q��gԼ�:����;��;�T�<f�&=�����J=�?n<��*=N�t� b���<q�0;
wͻ�;N=�,�������]=бm�vȬ�Lx��=L�I����<w�?=���<Z~@=s�<:<����H����E;FB����<�t<�kɼ��c=jmK���_<��;N��|r׼N=\�k=�cX����0f����_0=� L=��˼&"=	��%YG����?>=��,=PO7���=Qq,<��0<�����c=d��������<AQ�<*ۍ�~��TB������뿹#�_��᯻�U;�N��+�Z��g��;/�"��v5=S���:��<;͐����aog<�-�h�``<C=v{�H=F�:��Yf<c�V;�}7=Z�=z-S�����+	<¼�<4>��0��:��� =��X=w6:�s�<g܂=��di#;z¼�`/�fLǻS*�������`�^$�=;�5�"�o=�����7�T�8�-@�@u!=U�<8����A��US�	��;�S�4>ͼ�.�����We�爂8+(��GA_��==�h.��-;=�D=�fԼ�?�<������<QoL��6=�k�<Ո$��N�R�;r�>����<�]�<^�=k����U'q�h&==i��ތ<&�Լ%%;=��$=|�<.0�y�o��&c;��(���%�'=��x��K�9�
�<�C=}�;�F�����<!!=�c�Yk����<^��<%�":D�n<!��;���$��<.�X�~�<c1����<��<�=��D<�W�<�l��UFg=�7�<pU�<�x=�f�:¯h����<K=�jj<;x�<:W*=��<"~M���=i���G޼P���a=O?E<�&=�n<C�L=�ߐ�[�l<	������Ļb�W�(��DR=��g���G���;�c�~,���K=#�,=�إ<:3�<��Ի��z��qx�@�޼k���0��^��:�����;�k�ut=�j>� zQ=��<B�F��0b=���<��)��=����m�kW��@�$}?�}�׺1>＃ŉ�v��<#e��V��/7�<��=mE=�%�e��<��=�����N���������@��<�&��=~ݼ�0;�4�;"a=�� =qTO=[%O�$M���>A=F��U�<n�%=����0�S<[	=9��;�=�P�㗌��sj�Ii1=3Z^�A<�D�.�+=�=�,<�d�4c�<,�.�f5�φ9=�9
=�=�g~<���<Vs"=���;��<�!F<2N��(PT=,�=��Ǽq�D��2`���;�ќ<q�=�?���һ�\ʼ���s�=��D=��f�A/�<Q�`���p�8<*�J�2=k��;�?=�

�8`�p�h���f<sX�=�[�<u�s���u<�}�����zB�;��k=�g��$�0�4�c<=hj�<��ژӻ�(t�3�=�	<��C=�0�5�_�*�=;��+6�	v=��t<�
���>:=��Z;����`=3FƼzA�"<:ZC���<�i�a���2�� K���A�A�&���>=>=8ɼ�B��tW��PPļ�)v=؋.<O����=����pO�8(��] ���4��~����<�Jj=
��<��"=T&�B�J��*�2V=�ʼp�<�=z��?p
�8V=�ݿ<�T<������6����<��<:nA�ДK=�-/=�39<�R���Q��H\=��=ݧd<�ꗼ3!��Գ�<][ �#,=8�<�z%�&��<�}���� �;Ѽ��(ʝ<Jϭ:��F=yt!=�i�:{{����e�5��=�!=^S�]�`���;��(='�Z=7��J�2��p=ۣ��7<�ü���<Z�R�\��-�E=aJ�om&=��<$��<b��L!=\M<=�\e��O	��,�<!ԣ����W�w��;�B=^X���|=�n;z�<�^����?=�S=c!~=v|X=p�O;Kd(��[�=JCo=W�.��Q��_S��9�v���������<�#=�3=��!���h-L<��ؼܚ[�¦���%�������<[j�<���;�4꼦��j�ͼO��<�Y=�yu�E����e=�]�"�m��c���-��u��+���ԡ<��@�����P�<cqH=޳�<�?��YK�g��p�ܺB�:����-�G�c:��<��q<K�h+Y=����b�_��x�:;�3��B^�<Ɠw�i	'� �[�J %�o�`<nh�</���<w�t���W��}1�`-9���4��h�=��l<;d��ƀ=Zk�h��k��J<Z��;'Z�<4��.w��R䖼%����޻�U��pe<�5=��������<ڷ�:8(�"	x;����;�
�x�E���<Ą=�:.=ݫ�;8aO�MWV����<7>���K��셊��=D�<�w�<��<��=�`= ]X=�����3��7�[�Y�5<�`���}6;��'=�<� =8��<���XVJ�o~�B��/��[��"����֜�A�#=�;����.�\�*=,����S>=.�D=�-�<6ހ=W54=�?3��xa= cf��=�c����r�b���t<`��l�U�_ӡ<��_���2������d=2�`<"N)�K��<F��� �A���~�<���<8�����<��<��-���<9a;]�	�����<�	f2�b�X�S�+��j���&=�'�<��=/o.=�E�<0�=_�4���>:k���=��j�o	_����jR=��_��uU=��`�l�z�t�ɼ�(K�J�F<�#�<��:j?k��eS=둮�A'7��y<�S�5Yl�c|�<���s�м�ϼc�=.���'�<�1��zԻ`��<�ru��V<bAD�	�<�?��P<��U���G=Qb =��8�<�=B�<i	�(Η<�	o=ݔf<�:��\���ډ�j/U=�0=ߍ3��JC��#�nH"�!��<�>��̷<
%�<U��n���:=0�:O9�L~�=��������<ş.�}�<��X=�}"=���:��];�?ƅ=}̼�e=9��<i:����(=�f��{G��D=��:������8=������<�x_�
=�h	�����@���Q�?�t:����mC�nBm��Gv=M�<=f�<#�����м�.���&�<��2=�����\=`X��(<�F�F����<�:�Լ�H	=g�:�P-<s0:�&��c��b�8=.���m!�lwy=!
����Z=H,�I���V�=+���tz<��漸�4<�8�;�.��"=:�n��<"==��
�e��9����2�X=�i�;X7�<9���4==0+=�"G=+�S�̐C=�<��L<'1 �F�;/[�T�A���H<I�+=���W��<h&�������<�/=�pz=�Bϼ��F�>=gQQ�u54���)��l���'=�DK=q[j��=O<��.������$��6��2P��`��,*=MI3�b���~.�+冽mK<�t�#����/N=(l=r�~=`P\�w�=X9��e�<��]�<h߼�6"=f޼�1=H�%;SԸ����e1�K��c�%T�Q����1=�o��Y=<{O�VT�x�2� �{�B�l<y��<º;˯<= 4�(��<��-<�N=�K=�}=-i�<|�<��9�"��;<�<xnH�m�"�"h��á���u��M8=U��<җ<B��<2��<��[�a��<���<HWg�G����_���8;�(�2=���<y.=1+B�=�B<l�Z=�<<�o��O[�0'V���T�A�1��d������$A�AN��C0��Օ�;Y6���∼/O�=����4= �
=[v</�=z�h�=�k��_�<�<~6=(��� ��<�'R���D=uE�<��&�A���aH�!e=����<�F;ݪټȭH��=�Dv��&�<�C=~T�����<��;�8���=7夻�B�<H�����;@���u9q�y@=�廼K��<�"�;ȌN=|jN=~�j�x�=�@����;d�<�D��<
��+�#VZ��.=A�O��r�z�7�55�<�Ò����<L87=��+=ź�:J��a<`�@����<�l1�F�?�l�ͺ���
��;�[T�ԩ��$�<"�D��<��I;[(=��h�%=�1�׍���;����U=i�=�=������-�
P�����<��<�xf���9���O���
�Ml==Xo= �<_V<�J���2�~ )�Z���;$�<������^=6��:}�P=2P<L�׻2��E@���������QR=e�5�<k���<=g�	��X��d.�y]#�V����-ļjnB=��L�<��=���ńq=}�=�P�<#���K>=���:UT��p_=+��9=ji�jE=c�(��qY�� ���I���y<����a=�Nм`�<>�Q=3_z��93<�Rȼ`K�<�Vb��bJ=yF=�BE���	�ӐR�w?6=��G��n�<㾘��8p��oE=�8���k=�QR=$/���屺&�=$><a�w�v�߼��Q�0,P=l=�����'�X�L=BA��ɕ<=4M�{7ڼ8ϼ�ݻ.�;\���d>B� {����p���=s�h=�Is<����5-=�)n�C�$=�� =l�;���>;�%�oA�ا�=Gjt=��=k˻n*I=��G=ӡ =�/<5=�7�<Uz<=t>
=��߻|�&=�
;�f���#����D�����y=,�@<++<o�*�"���`(=��A=�;��=ћ���	�<���<plM=?l�<�#�;z���@��<
�)�|nT�<�<�4�<����s������8%���$=�a=�<M���5���T=^A�;���n�!�$�<��=�>������O�Jl=c��;���[8�h����-$=��l=�(.��O<v���O
��F.=���/�y<�,]=SB/=�
D�%�<; �X=��<�<}�'���<��:.�<~�%;�����<��A<?7q=�&Q��+<w����S=Y�;�9y��\I0<	�=l��α�0�)�2"���3=S)����2�N���޼�[c;y�����3=�w�<)wI=�&�=��A�4c>�������<'(#<� �o9=�w)=<ʂ<�-���<L��;�=��<�0��?�`=_��<�k.=�s�B�\�� �v����1�<ե�<�D�LF���;J�@=��;�	�_=5)���"�9W^�;�7�<3�<A'��'�(=(�K=����<h�A��])=�f�;X۾����xE;<߼?l����%����<�#7�v"<�9'�O"���7<��\�|���I�<=�<��V�e1�<���<}���z*=�`%�2٘�3t;��O=�e�x��<����3�<�h���W=m��,7'=�z%=������$<E�>=J��<y�F��� ��-=�_K=�j=rK2=�e��{=�����P<�!�<�v=ۂU=�1�<���V�?=��\��S;d��ʴ<����P�<�<�=�� a5=^������]�k��<�D�=�F<�)<*Ψ����<*�3�di��:�)�)఼+��� ޼;=<յм�s�<F�^=
�;=ҡۻ�SC<*6<�O>��-6���g�%Wμ���=1�<!=�8=��=o:=P<��k=UO̻-;¼�:̒F=5����2=�U�;�p=B^=:�q��(��=��<rj�(�;�$���<:�\�z���3Tc=��==��B�/D�<�b=?��;�U�<>J��p0�����/=�̻���)p<!�"����>�2=v9a=��=T�=����eټ�Z���;=G��;�3,�.NI=<�c��0=�J�<b��;�@8�ݜm���Z���T<S J=(�c<gy���z�<��B���Y�=���H �>='��;�B3=b�m��=�:��<���<��)=e�8�3 3=����,g|��/�<�5<�Nj�)�Y���X<M� =��8=�)={1%�����Pe���'���=��3=9�?=w_=V���8�<�-=k�=�՚��;��A=�ټsJ=�k���`#=�.<�f2��%�<r"���om�$Y=��9� j<vZ��{y�3a��v�Q���(=v�;�l����7=r�m=����h�
�+=�=���:��~�<�o"���)=�c<�q����[�4F ��%�<�=K����<�$�<�~<bC.<k1�;u�ռ�'<�溼<Kv�:V7��\ =�jQ�J3<5D��c^��r���P=���<�gQ=m���k�<W�d��<n��C�z-�����#�����3=�U+=�0ݼ�c4�@Zj<Ө=�r����� =q�����N��fW����<���H7�<{弎�Y�kã�ƻ
]��D�z/������<Y@1=�~<��*=�bB���D��O���
=�X=�H���Ѽ�M=�o=�g�<p	,=l���Y�E�Ú�<��U�u�R�r��<�
\��3�ᚻ/|�<���=21P�C\=c�.�=��<O�<����s+=��?��<;���b=5�P=N2a=���<9�����9=!�w=�v�s�=A�0��Q���p��F�;=:	�<[�A=~�;f�t��.�\<,�=ƙ�8\��<�<.=2�<����OU��޵*��#|�?o=��=}[��-X�<:5=Q�*=s��]_e����y=n-�y�m<p.S��4��r��j��:=w�s�i��wnz�'h��~H���W�	�*��V<=p�;���=��(��{�;3đ;��%<O��<�&4�a��;�-��x.U��n�I����8g=u.����e�Fw�<x>=0�c<�a�;��M=�
F=���<�R�s�<��Ҽ��C�$l�?aj��l=piC��I)=\�5���<��q<�[=�!+;!'&�b��<�u$��i<;���\�h=�fY:w�K<�<���wU�re<w+�?����B��~�9�k=G���=�<��=B(R���L��̜<׼����<׮@�Y�S�#w�>�E���c<��<J�h�����&���1;cżd�6=:]y=Z�����:�(=�i7�}E�<__���%=n0��S<HG7=|�X�6�=�K��d��)��<�-c���8�`�c�í,=��<�1-��)��ZYS�� ��vb�A�U���� ���w=&�<D���?��m���f��S���?�2��<]o���1	<s�?�)0=��:��1�x�����@�����=7x"��ͻ�c=#��kO�N��j�/��*=u�@�+:<�2�廄0�<��^P�;�#����<���9J)H���C��v�<tp�<!S��̪=��o��bB��c=�I��
�<�@�<�S�<e���~=d����4=�}�<�j=ƃ=\���Ě���c�G��:=�t���;LY=������A:5�E=v;LY��Z<v �;���<���<��Q��k=�(\�E��<~�d�d�
��r6��sW�$̼H�_��@���<wK�<�V.��-�:�vF�� G���s��<89-=�B�����:� =�g?N=;@=��;�
B=jhy<Y�ۼ�_�VἚ��� �<��#����<c��<A�����<􉳼���;��<���<��<6��n4��k@��b%�F|A={����c'=��+�b.<�k�:=ƿ �fw��WY=�Z< "�}H�;c<�z=B�ż�ۣ;���Мd�V8[=��+�Ö�<S�}<Js=�]�t맻÷j�ݶ=��=��@=�"=u�����)�|h=|�t�U<M�)=]$"�ڠ=�c\=���L=g�"�\-¼݀I��p4=D"Y=f[�E�\�Z�<=�v=���</��;|��=�	N�D�@�@�߻����<Qz=@��G?n=&�*=�y^<���������<D�=;9Fμ�p�={���It<��=�=Vɱ<�\�1r���<��=����Pe=��G���<�G�|H���='��`�A���=�����0��X�	={���'N�v���A�<�8�<N�F=��A�D�f���o�;ʳ=��</�O=�Xc=虂�E�<,��:��/�{��<��μt�<B_ؼ:y=�HG��bK<-�7=�|��o�;>�o�(w�<B> ���=H>=���<�<�<��;��`Z��C��\�<`{�:[���ܺH�͚��aI9�U[v�>D�<�
;�C#�XI�S�W=��&���=am�:�}8�U@�_	�֢3=�([=��ҼR�N=��i=əs<
�:��=��<+�<|�U�]��E�<}����,��ݡ<���<ɀ��^<���-f�<K����1<=&�5=,<�;��O�Q�38����!��z�3+=��/=�ǻ�0˼�f4�?���J��F��|�=���1=��J��=�x=b�;��V�Mz�<��%��I-�g�Ҽ%=��H<m��<f&���=��}<�<<v<�F�=�*$�����j�X���ڼ�5N��-�︰�
<<h�9���>;[�м�L==�i�2=fvF�~<����Y�-Ӑ�8�ټxQB�hn�<��=��=��=5,/=�����̍�<klW���
�����ݡ�<є��7,������� ;d���g	��@�;��9;��<�'�<'����ٺ�tP�<�-�;C@D=��#={.��1�<��e�#(����='jT��׼v�<D=���2k=i>@��r?�w�#=Ta��ɺ�z�N���-=Xoмq`c<���<�%!�E�j��zD<K������<G�%�~�Լc�;�f���^<�Pi<T�2=J�*<���8>6�j'�h�U�o�n�;�7�<��L=鲫�O=7���q=�<�ŝ<��9=���T=��k��%��np=��M�""�;
^@<؊<�Q�<>�}=p�+=M���?o�;]U����z���.KK�\M��3=��u<��<�^u�b4b��\<�ּT7=�g��xD���,=b�_=o��<�n'<�=pջ�3<�zg:�g,��к�=J��f�F�*$
=;�i��6�`#D=��a<��<��N��3;��[������#=���=`+=w/�:wn=iVw�sYż%�=j����$=��l=�h$=���=��=�t<���0�̼�w
����k�j=d�ɼ�=��/���9�<�<�=��E����;���:(E=C��<��<wǎ�D�< ���=��̐��|/��SH��2C��=5=����?Hr=Y7k�t��W=SD�<S:q�J�<�g=���<�X�����pX�x�=��=&q�;}�2�f10��x1="�ɼ�P�<*�Ｙ�X=J>���[=*"�<��E�	s'�RBV=��<�dC���@=ۃG���<+�̼C1�<G�k=���=f�<�`h=���;������_���+=��2�*^B<?$�L==X�)<��p�xN��V�<�����м�p�<y<=ݖ��L,�<���v�������Z����<��Q�ҘM�܈���x=�0�<���vk�Q��o!=ݏ�<��< -Y=b~ <ϋ���޼��%=�;N�e=����|�;�n2=~�R�]�O����������G�`�(<��=`@=�"���)��oX�Qb=�A���8<o� =����E�����<�>��>»�x�RnY����<�2���):�=Ƨ[<������.=(�ټ��<���-�D<HA<�_�=��ȼ���:gS;L�(<�:=����i�=�����7<�֢�4J=��ͼ��<�<���暫<L�U���<r%=U"ǼyH=ҝ����r<IZ�9B;�<^ZW=�qP���<b=����("�B�!�h��ɐ�<4м�<���:�h5����@q��X��%�6���q�7O`=e����O�== �B�{5=��<m�<�VZ<S';<��[���\��x=���������I=%vS�$�Z=-m��>�H<2Q��=<6�4=�|_������p��6��HeG=�<���#=��n���$=�o3��{h�:��<�u2�<��N<�Kg�q�8=��<n߆��|>�Ƭ���<B�׼�� <u?Q<��K<dc�<�|�B��;|_]=dI�<��r=��9�#�N=N.=�f8<���E��q	�<1�=�3=�:�;�o�eQ<���_J�<6	��Ԗ�	'��[	=Ы�;���F���df�<Q(h�u펽��d���\=O�@=���<K=�=Ѽ�N)=EC�<ʑ��VА�dY��A�<��}=�E���p<�	�>�S����=�&$<�B�����]���L���<=�_�<�o<g�)����<=��<,=@�
=�K��#=�#=�f!������úPO=�-,=Ύ�1-i���9=�9=��%!�<J��<e<b�e��<v�=;Z��� =q��?=�DG=pG��4*��+=���<�zU��)w��>����VR]�#�=���<;u[���:=:����
=��V<+m�#I=�_=(l����<ό]�_�����;���\g��1�J=�F=�=�[���</��<�=�)G=�?=V��Hx<<z�W���Z1:To=�fH��-\=E��[6?��,�bR!�RJ���6�4q�<�B=<��*;t�@��To=�;�<��ü���;��H<�⼬�8�=-�<m<�}<u]���mӝ��M����2����<j�=��[�|����D�d:=���<�Y�<�#O�	�/�zb�4%��	.��Wb�W�j�n�5Һ�{T�N�s�EpC���`�=H�#�m��<�+�a�p<l�Z<#JL�#�,�{Sἦ�����	=dvмG/C9�d�<׬ּB�=�j���e����<�|=��s��@�<�^r=RQ�<av�<��<���<7�=ʇJ=Q�< �5�ʩ#=�
�_���H�\����E��Ӽ�<���<l����|�c�<dӱ<��P�;�b=�5;����=\	C�i?%=��x=�m=�G�<2CF��9�:��<���;{�<�Z=��=���B�;�-��%=��u:\�M;/�;��=�)�XÓ<Q4�����@��k9�F<�v<�!ż2��)V=٪�<SSʼ��u=�!<�Y�=�3P<9a���d����%�C=�2A�����1ݼ��=w�O=Ռ=��!=u�<�T[=��m<��=�b;="~^�������(�].
�^'�B�vUu�{���f��;�E��<"-�<��=p�;�F���p�!�	��,���� <-A�;7|��f�<�1<+�}�L�;&V�<-��<|��<7��i�:�_3��μ���<�-I��-=�_�;oB0�g`�<� ۼ"[�5F�<�FG��Ѣ��qs� F=��;�	�<a]ü�b	=�ׇ<{e�<�_��2�	=򸩻<�;�-����=0Ib��C�;�Z�y6p=�=("�<�m�;�n�������=q��1|#=A�&;-w0��=���<_��p'd=\�%�)ܼ͐9=li<R ^=	3=S]=�<U�f4Y={�<���uS=Eyp�/�<�}��UY<���kq>���q�<�x<xQU=`,d=��мh�=k�;p�U�R١�ݷ=��<[+�<�9�=:�w�d���c��V��
7�5IԻ��9<��5��p(=���=��<�%�;e��<�k�<a�]�x_�;[��Zak�kv�W,=���n3�%�⼄������%=+�Ӽ^��̅=�q�<�T&=��]=���;ܹ=?�;�}��M����8=˚�	^d��5=83o�X%A=�%�<�\L=Ca�=W#J�P=��(�ֳ=z߼��=׉%��:=a,Ѽv�<%��<IC���(=MG=<y�w�5;�Ҝ��	��<�W�<��b=P�[<�=�Au�<�K����V<��F<8��:�.'=1�q��7"��~������ӑ�<��?;��<װ��i�<��C�N42=��;�K=~�X=}�D�ҥͼ�U,�(R�<���k�����==�N���A=]�5��k=�U��@_= ���y����=�7��*=�hO= ��<?�	=KA)=<��m�<�{�:�%K��1��.�<^�:�J�<*=��\<ݕ�<��^W�;�¼���<ݾ��hl=�o����.��=;Nrh��L�|$<V�������>�j}<�\�<��޼�Ql��2=q|�;�=�׻�/��0�W��cE=G�ռ(��<p?�<m���֑.=�{U<P������oK��v��<6M=w/6=���<\�;��f=�S�<�#<}�O�?k=焕�,L=u4��z�7=��.=��=�o��=W�Q�Z@�<]ֽ��E�<濔����]�<${2=��*=��.<�%�<��8��R6=O�<�m��� =M�޼&;��;<�E�9I��9��A�F�;��Լ�֓<�R#�#�Juy=q�n��7��Ov=-�9���0<2p4����x��ފ��O�ER:_�,�3��<�m��t��[ކ;�@������:X=τ�<�Մ<G1��"�$qW��I�:,������+�#�;��:�:F<@F=�� ��<U=+�i�����[�ּ\�p�ŵC����x�<6�L��`�<K~�<��t�C=;=lX �gE�Db����v�y=�*�K�#�<"(ļ�=�B�蓘����<kQ=,;�[l�<���<�p=����Ҏ�<��L��*P��0F��p�<A�u=5�$=�<��=�߼��c=[�<�z;j�<�:=���=��:=��-=�ł;�33=$ּ�H��s�:-�8�$ɰ<V��<$���(:Uu��؛��Ӡv=��o=�]q<��:�d��r��<�脽N�Y=��.�`bμ�3=��:�Ĉ���M;��P;���<�<��r=O��<j�k��=�����p�Hg�<WI:}��:&���!�=c2����_���<Dn==*c�oм2(=�
�<Qu���i#=%��Ⓛ�ju�=r�<�7������;<R'����<�*�C{�r=���!:�?��<@��v�<��=j��	=�����X=��9=��<6��<�x=���;B��WS*�e�S�;U5=��=���_�H]=��9�aZ<A5�=F(����<Ӵ]�9��<`�Z��UC;^1��c �=ws'<Pi=bK�:g=����Z%�D�p<78��Y��;��4���*;��<�x�<j��<瘛;AY�<�tI=���	��<夨<[��;;d���P-=EA={~����<��N<��D����=�a=�;�e"���=5�E�E���=B�P�N�W͎;S��4�<⪩��=����x�<�
�;zV߼�Tt�w���%��m�<o=�4V<�����|���/@ �*�w=�=M�=J�4��u=�V��;��{<�%�9׳���r=��D=&
A=�l������WE<~1�_�+�2[��į���CP=_j*=̍!<�==
�(���<����+�5=��ռ0;)=�[-��8^��ﺼ�����y�<�=�)��,�<F�����ݿ��m��+'�D�˻�Z��UZ�C<��ۻ����u��,K�ga�<��Q=�=�n)=6N������%�-=�?'���<yS=k��>��<�~<�p;�����g���R}���]�sμ[l�#�X�+�I=��:=i���J���<b�B=��2��Nl<�,��c�YGq���`=] =]W1���B�?iM�I�8<�x�z��=x��o�;��<��<p�=-5=.�1�eM=<�0 �-�+=$<n+��r9<�d"=��m��Ņ=|��<'k���P����<9C/=�v ���6�b=Ou^�ʮ<�<�9)O�P�<�#��=��e�%	�*S(=���;���=P퍼#�=�t���_�Y����}M�y�⼏R��%�3dN=�zm�L1p�2"0�(3����V���D�^��=,�!��ͼ@��o�����Fy;�T��ܗ�[zG�S�;���<� ����2.4=<	t>;S-}���=�H<�������d(��t =���<�+�<�O �5j:��2	�'�=��ɼ�Wû�9z<qt=4J=hw��P�68=V���uB=5�<J�=�oh=}[Y=��g=3Rݻ��t=(}_�u1�</ ��P���s�M�(=]�=3��x<��A[һ�zo���T=����׃Q��@����<�T�M}���k=/�����<��h�Y�B��������< �,�Y�g�t�.�4=�R2��^��a+<�<���;ܑ�<��U�9��
�=0�缙�<�DK=>*�A��<��������N<^�2�M;o�<q=%�<�����;4=u.ļ�B�=�3@���:��+�;o_����=�򄻶-l=�-K=��`��>g��7�
�a��RѼ/$=�����2=���x,=;�w<Q[���=���<{A�����:��=�P�_:N��,/k�X�<�v�<�y)�@= 
=�\=��<�ow=Z����0=\���� \q��i	��� =��H=�&�<^n�=l���C�<��K�Er���=*/@�����ZE=t��<TL߻o�Q��Պ= /�Hx�9\�B��?�>==m��=�I)=x�;/�<{�|���<�J=���tQK��+Y���U=��ؼ��<Ξ� ��_���*a��"�<g=�<:�^��=�<K),��˼r*%��Ѕ<mvb�1E`��lݼ���>$=M�D=r�;K�<�>��H�<��9<��X=ހ=/�j=ж����<~Z��5<i�=5�e�u�.<��<�A���&���=�^�	_�}U�{F��8(���4=pw�����'=���=)d@���D�3TW��M��k�<#���^�<�'i==�?=$�N��"R=K�K=9T;������^=��Ի�vL=�O�o��<j���:"���=�CW��L�<Nv��~��8�����3<�i�k�|���T���<@����Cq=��=}o�<��������X<�ᔼ
wQ�{�ͻH�=���<�Kw��/R�=�S=�􄽈O�<�?3=�5�����%�Ω����:)5	����/p<uR�<9�]��@=*�=����y�;�W���`�7^�<	 C���7=m}�<�μ⵴�#�#=8J7���<�`h=@����<���*��ku.���!<�4=��L=�:�	�Q=�|F��E<��-<?���7=)NX��,_=��[;���<��|b�3��3�<=��<} �C7��W�hl��*o<�*�R`�p��C:h;�<_����.����:��1��E��g<��F[�q鼱Ǫ�HTw=hy�<?c�<Vt&=���=�I<�c=��=~����*;�2o=�,E�)겼�L$<����/<�l(�e��;Ӏ=d��<H�0�!=P�,�[�F��f�أ��(��$��2��G��
���G=���<���.�b���=2y�<��=
qۻ���;=0�X=�%g���Z=�Fڼ�=m�=_��<I�R=PB��= ��<@X<��<��)�y�=w&=�)=&�Z����c�X��=m [���O��
�9�zD=M���:�,��A'�Joe=1��<Kv�*��<.�$s?�Ǡ<�u�<-�������1��*�;]o-���o�'�C=�O�����l�<�dd��zY=t2���<s�=�	��T<(�9<�W����<�3�<ή<�����<[O=�&��tE��y<OS��(���@��(T!=|$%=��Ѽ{�8�݇P<��B���!��QD=k�J=Kx<��<�ʊ<��;�"��5�5�``>�*�<t�_=�l���	=��<�s(�_ �b�i��d%����5<�?ּm4N��eE=�=�;S�뼲V��($�$8=4�G=AZ��&���&�=�@=�/��=5�����Y=���';S�|��7E��?4�:���;��<?��<�80�֍�;��A�����b�h^S:޽�<a逽ڊB;�!;�<��^=�x���{��<n�c=8c�<�L�;�3���J=>�=*?�<�?#=�@���r<�T�<Z_�=}��<{v=��ἃ��<'�̼�b^��b�<��\=p��8�G=|�;���<������=��g��:9�X=��v;���%U�CP@=B;=�]_<
?=`����<��=wP�<��»��=𑿼A ����x�ؖ�<�-P�r^ݼMP�;j<=��2=�A)���4�+́;>S";	��<i��b�[=0RS��<��r<vB=T�9�iMA���?=�-���<.�4=��J=d`2=�^�<��<3K�;!�8<���r�=`	�:���<�)C�o@1=�0�%�(=�S%=,㙻Y��l8�c8J=�ԫ�Ʉ��r�H�<���<j���"�<�;�T�Ҟ����6�0/+��+=NW=fWl<�dr���%<�f��ߜ��-�=�S<v(�7�Y�E&|=��<1��<)�=Z��<_!�<��μW,>=��*=0�=rMѼ͍��:a=�v8��O�ٸb=?��<�Ph����;^�F�a�C��!=h��8���:��<�.�S��;��[<lr==�<ğ)�� �_ّ<���<�,2��^�<�����4�α��#��$%�����<A��<ݍ3=_�<6�<*=�</F)=Ԩ]=��&=�=�x�����2w�<��;�����@X����NK<8&�q���.���\=,ؼN���v�^ �<;%�T�I=<
���JG=T�N�R�<�3� �s<��0�<��ҁ=�C�<O;<����i�;ė^;g�Y���b<����H�:<�k�<�@&�z�μ%�<{�ݼ�W=�o�H��)�<�=f�Լ�6�����=�ȓ����9�Y7<���'$ǻP�*<��<�� =�O����� �;�Y �S�3��r=,q^�ӕ�)��R�2̼�~Z�� /���`�']��S�<�
=7��<�lb�S8�<���<D[Ƽ>/O=���)$�<��/�xYb�=�; ���������A�:�Ƃ<l+=i��zt`��L<�SQ�W	�`; H��o%�>9=�h4���8�+N��CJ�y�;XV=�};<�=j�x<��,�t�q;��m���޼��D=qt=|_��aO�<Ptz���t<UL=m�<��x��=�O�<;����;�C�	��<c��<]+��f��ݸ�<�n<	���b����ZE�Hn���J<����� =� =��==�?���ڵ<�/��j=I�C��-<��\�9�ɼ��u���t��2G=�l�<'�zM��5�e=b�������<V�NE&=����	f�ɲ!<�(�!eb=���<L=)b�꒡:Q=V"��.���w%<�%H=%��;a*=7�S���H=�Lμ�m�;�S[�֋��ȼ�R={�;�$$=zM���e3�Mg<1�M�E�=�A=��G���R<.�h�dr@=�*�;�����<�q��A� ��;�����p����<9:"�t�^�vv�x����R���D#=�t�;�:2v�<�J;u4�qF=Ƙ<�X�9ج8�q<� =�s=��q<ܒk<e�3�O�l=�qP�Iw�<��n�hEn�DH6��$ջ�kc�!��<�;=���<�(����Ƽ����
������2��3����b=-GT����;��|�����J��m��:\�a��u=ޡ;�A:����<��p=C��������=�;٘�<�r�;�=4O�<��1��_=O�<4�K=GW!���"���^���l�r��;��6=�6<E�����d=�p�d!
<�b�<�i=��G<�j�<�a�YX�����<yc��^<|M�Cg:���`�����:�8r�9BD�\�c<q���0=|KA=�\�<k<M�:��<�=L�S�a<7�'<��<��<�%=�-�]� =�R��?�7<�c�?d=%��<�����UV���<�̎:x�U=�L�j }��
=-h;��=�=;����j�<uZ�%=���<�VX�)�ݼ�u;��9���̼���ql%<�M��$=iF=�P�F�Y�� �<�0=k��a�E�_<�I=-�=J�o��޼��o���`�N�Լ^�<��R��̍=�iڼY�;Br��	�<@�Z:�}��n�<��D=[�4=�倽���^G���<���֥�y��<D�ܼ�L.=�a�����{�=��<؂1=5M5��]��_/���n,e�4Ǧ<J>���"=S��<@
�<�i=�	2��k��vj�/�R�'���K=���<�$u<�S=�P� ao�?���;ꭼ�Rż�帼����O༬p?;�h��%=�/!<8��;��;=]�<��<��x<�?<a�;�'W=`?�;��t;�B<�?�<�7���vn�λ-< �[��4�~��9}�D���=�L�<�n��8Q�$I=~�-=nc��̈�	^s<׍=s�<;�t<1�<W�J�S*�eӻ�U=ޝ��Z�=�~��bf<�z_�<� .����x?'��/C=zL>=�_�;w�L=&�=������#�;<"�=p���Ef�� eV=�ü�\	=d�_=�/����D��C��lp��xj�F�X�*�t=�~n<��!��/=Ɉ�9w�U=j;��(=���z���-��\*����<E�3�T��<�M=|հ<H��<6��=L��<��<ʰ�O�=@�˼��߼�AY���
��rI=<ͼn��F�<˂�<�ȼ�»*t�=>��ק�<҉��w�0�Xy� ��=�aE=0��w}<w���3����#��<ȆU��=���A�E=�`�<�|#=1�=k������L��;��:��u�<&�Z���Z���ڼc!=/�<D�=='��,=%���� ����L�T�<��=��=�!<��N<ѝj���g��5�<~�=^y/=w�S=r��� 6�J�<:��</D=�H+�a�V<U5I�9,P=�'=�_<<�=Q;�<�<N��<�O�<M�~=�g�<�R�Va6<�-�NY>�jFA<x���pf��U'=� �(�P=�܋����
Q�<����:�r�B=�X9;��t:�AX�\2�8?8���B�ro���`Ƽ�����Ҽ��D��Yq�U�<L��	;�<t��<}�&����<�lļ��἞M����<1�
=!�K�}�c=y��b5�6�2�0=�X%:��.�ڜ==:#�_ņ��P�=~����c=\e����	�<�����_��$Ic���?���F�1���CJ(��_=��,�n=$켏�	� �Z��X�#�=��a�?[�<�*�<`g0�,%;͊�=ϖ��n)=���=�tI;,G�<r֦�#��<�����q�]=�Z%���<�o�<�q�h'�<vbz�*��<D����.�</�T<{2$�g:�;~��<�g���;�P5=X�ݻ����8�j-ܼb��<x�]<�OL=�<�<�������<8�A�pl�q\ =�cE=�ư<�-�<�ļ�=���<�\4=����$=��8=ep<HWW<v���/=M��;S$	=m�	�7�=ɽ'<s�#�b�
=#NQ�d=�;`�ϼ��2����<�3�<^�=�Kڻ��<�Ⓖ���Ŀ8��'L��<vp;v��<�R����=Lm�=�Ep���_���\=r����;R�=�
=i�="�=�Gq=;�<�3P��2?���:���< p<
<��t�=���9��;���<�Zg�^Y3=����o-=�]��္�<[<F�2����^8�<��;X��<���t2�Zv$=I����=\?m���	=Z��;��� 9�X��:�ּ?�]=G܅�a˿��VN=�~��2$*=l1c=��<�Ïż�9=~���cH�1Q��խ��婼�
���<�*L���a�Ҡ<��=����,=l����D������V�<?��;��<��I=��_���Y���]���h;���;����H��r=�$�=�<q�ɺe�<L�G=k��<���U<�bZ��r�����:��3��%�;2�<J��<�0(�e��<K#
=���<�t�<�k����=�=/=2ud�]΄�S�1=ߴ=���<�6o�[FC���0��YH��;���<�d��'�<�P�X�h��a�<�!=��=!����;���</�=��=Bn=;�Xy=�����:�t^=�?`< V=�$F��A�;k�$<�ɼ�if����-�<���4<�z�2=>�7�@�B��Ŏ<M^^���A=� v� $�*mb<p�=S��<��;$�R=�Z=��8��ѝ��	ȼ��=��==�Q��Ud_��2'=�J�e=�O���	=��{�J�ϻ-���%�;'؏<4�H=-�W=~=L ��}A=Q�3���P�G<i�+x4=8.�<754<'�Z�8P,=78=�#U=�9�;ą�P	�;��nXܻ�<q/�<gJ ;c3����-����<"�x=�a���WC=��k���D<�v����;Ĕ<��J=��������)=�;,=�x�<���D��<h�����=d��<�5=7ۻg�ļ��ծ��qJ����=(�9�m�<*"ؼ���NcS=�=Z�6��BB=�8#=�����&<i�-��i;�� =C���hI=�T�H�{(~<��+=6Ya=����=�}����߼��N=~4=ӁX<�X=q����0�E�ּ��<kՕ�٨���r<p����n��c&=*Ub<��e=A��!F~�$k �d���;R=�y"��+=zK�Q�������;��:�<&�ܜ��36<1�^�4�<~��/F=�#��	f�.�9�K�o:�<�
Z;}Ղ�p.�h6�ݻ?=�I=0���<��0=�3�<A� =��
;� ��v��[�J=��m�C�ۻ��I=+;=�����(�F�� İ��g��'�	=㚬<P�$�L|�;��8��8@=�K�&M�&;j^=�-�<,G��/ ��
��=F��;�L$�ۄ��B�< ��<ãv��B�=�"�:!h�<�u>�>y<�Y�
ȍ�^��{�?�ߌ\=	�p=g�12p�\h��}<���W�=2Du��a?=��^=�m��sq=*p��~F=	�[Xw��:4�=����!=��C��1=�F���<l�<EY��ho=��J<}��P�C���W=g3A=%민HE�<�҉;�|=��꼫˼�z�<�wo�@�<�����Z=q��;�Z�<R><#P'��~D=ز|�x��G��뜱����"�7����<]#�<
W�e��fs��qs<c�=]�k=tV�<���:��*=�+=��9.붼"�=�U=f�K=�h@�L����3����Z���Ij�B�¼�/:���=z�6=2�}�e똼�T���R��rԼ�<�<�;L�;a|�<��R=�yt;HY��s���i\ =k�F=j�=m�=&��V׼2+���̮<�5�=%
a�� =�=T8Y�)��=�&���]�5�k��h���d;�n[�Ǒi���1��	X�ڬ�<��:�E�_`�~'�<���<�>���ܼ�μ����;��t��-���&˼{B�(3<를ka��1�2��N������*���"=�F=d��t$"=N=X_@�.Sv�K�<���K �<��<�7����4@�X��<�U<(R��m�D=#Q:<�;���P=@�ʼҥd���O=z��v�<o8�c�J��j�;�
q��l�<�e<2�Ӻҿ";���<�_=\������͉7� ��<��=�ڼ������0=�G�<���;��d#=�&H=�� =a�~=��j���Ϻ��q��j7=�3�<U)ѻQ�#���0�U�{<��!���4<{<Œ=�ւ��ĳ:�V=2mu=/W��v
��^�G=���<Z4��y;V!Ƽ�ǲ<?*��rs=\A$��=�_���+���ټ�V���<H*=��e<8��<)=�%T=E ����<=8K�����$��y�<L$R�Z=�K=���<<w���X������=xA�;�����<X�I=@�$=�38���<r⏼�^7�Rh�<��6=YH=߿����<R�s��;�c!��	 <��6<��-��9\<z��<�q=�����o<��E=3�9=���<L�	=B��<�uW=vk�JJF��[�=�������<�` �fv(=�~B�.�o���#=&��:����X�<�X�;��#���<���<���;�l9���D=�/�<M���k��-S����<0- �#Mp<�-�n��EO{=s��<o�"=����|�T�)_<��޼���R=	�c<�[��&^Լ���3�9�RX��k�y<Bb.�e�+<�m�<�����v5=� =O��~<�v�/=����<N;�<o�<H�=�	���/=�֢��b�:P;=�M3���&���R��R�<��(=E��k�F<�;���L�]�����;�+��[=��^<�:~l�<!��;OG��-$�mf��[UE;�*Լ�ͦ<�H(�u=.-]�\��;�j<䤶< l�;ֽ<zT�<���,�a=�O�<�=g��<s{=�=5=�ּF6�<I�9Wm+��?��b9=w�"=��h�"�<Rw=~7=�?껗�G�h�#=A
�<��h��~���~(��F"�n��=�I=��<�d=*�8���F�{��<�[a�2Y�#���J<jz=�P,;2Y�:=d�<@��;x�8��R�qټEI�7 �<La��,L=�t�;����iY(=9��;��$=mȾ���<2����0¼=o;��d��kd���3<%�=N0b<qw�<�Lټ��+<�A=�I;�I���U >�L�F=��P��잼c��<�|�ŭW=؂��iL=ޑ�3�=�t��!�<Q�=k��{��(=F<�L�<�.��U�<�=<{��<�<�Z|�<r�k<���+����F=L���oB=J����< E��5i@<I=�<�	F��C<?�z�����X�92�^��<Jo�9s�=,�=��:ݼ����a�=Ťƻ������-<r�4=>v¼�����!<hn�<���<���O[�;@0=߬��ݻ�H?;�x�<+���F�Ļ�*=�BҼ��<u�3��ŕ=D1=��W=:�2��X:cN���$�<��%� �B�vH=�o��J߼�(���j=�`}�
��w�<�}�=n�;�=2�<��<!�S��@��%e4�:U�<C��<#����G�d!1��d�m��#�D=w|�<hA�<�.5=*�,:��<~˃<nBs���L��<k邽�12=tR=�\=�ļ�&�;t�[��Ȉ�5��<��<�)*�}J��&S<a$=�8�m�=Y�b=9�h���a=�ҝ��5�<ۋ*=gw=&�:�*�j�����u��)=��<=yO��̉�;!(ȼ��q�ze/���X���\=������9)S����<K�=\@_=�4��@u=T��x-�=��6<�5=c���,��<ɟ<��_:��X���!=Y�N=������;���;`��;�T.�":»&i<�����!�:'��G�<��<�j�<��<�Q�8��;��n���L��Ѱ-= �C;)�����^Um=A���^<f�=g�����=�	=�^7�t K�� �J�9xټ��<ɨp�xJu<k'�~9��������>����7=��V=�Z=�f�<:�&�0�W��<�0X9WZC�(�=π0=�C=
��;$��;���;�� ;�fD=�Nü|~�<��8�F�&�u�/�П����W�e�%��gA=)32=�_	��K<��8�,�=�����-7���=SI6��t����<j���{�;�=Z���Y=ڎ<=
!=��!�CH��?q4�o�J��o���*=�q=T&��Z�;r�=��$D�#����^�X~�<f��ڂ\���<�Ng�8a=���:�N�;�%:�*�h�80�x�1=S��<�ˠ<ox���ٹh��<�J;� �����<���<��ͺI�K=��+�hN�����;�<j=.�9ϻj"E�I����P<_� ����<!@b�j�=6C���S;�;��s����ʌ3=D�=�̣<����+�cA�<���:����{=���H�e<;&��lQ��9Y]�j�<�仲(���s�G��� ���f���=&�=�c��y@��G��=0����l��[=X�<a�=^k��5��=?�6:�SQ�4=��=����m������h�1=���2_f�;%�;�l=��|�u� ��m%=�	=σ�<�8=��d<��;l�x�(xU��?� ����<
2�<M=�;N�<�Y=K�=�01�>B>��qs����<�}<�)�5�f����<���-�<�~m=����9�������`?��vY�ci��~R=�"<S�=���E��^����/�������o��;�W7�+w<�I�M8q���<=����"!�2j=V�-��=1�F=V�D�i���9�<���;m`	�x�=Ȓ�<y��� 9�����
�,�e���/�G=8�@�e+A�&���x�K�A��V�<8�%:��)���o<6e�;k�V=�]o=��=zb=[b�<�O�j���E=����C=Z��N�{=��=�/<{��7s�<�8��N�2;u�(�~~=��<=��b�_��=�����<U�(�I?��qϼ1�%t�<�R�C�n;��:�C|=���:�ݼ1?���4r���
κ��������&�9�Z=r�,=S,=*��VZX=5���L4=#�<�6Ѽz����:I=3���O>��P���4!����ɼ��`��FY��XJ<'���-K�'��cF=���������< ���E�D8�<�91�B�������YO=�m =��==J���!�;`����P%B=[�;�6����::�����f<6�*=���<�K=����=��X=É�N1 �Qn=~!ĺ�ͺ�=��h��*5���(��}�<�7��7BA�#�U�(�g�٩�M�c�м\�=�k =4W����Y� <<�;ipz�P<G����<Z�O�7U���oQ�@m=� ��(w��܁�<�$��Ѧ�<Ĩk=j{l����<�9�<T>C�C�#=,㗻�]��\�N=R�?�<�e+�J?l=!��=�K"�0<h9�0��ߚ���<�恽�&=��3�]<i~�;����ؚG���*=��N=k�	=jT�n���٭<q�E=�jZ=��^=�Y*��< ﻼ����`�=���<�g��=p/�����U=�Z6=�G����d=k�)=ߦ��̷<ȼ}�\�)�&�6=��k;j���6=�U`��c=�#�<��<�s���$���L�I�@=Dx8��	<f���,��K<O:/<e+.���k<௝�q� =D��<;��1��0(%�� `�V���H)��U!=�;B<�v���<{�%=^)	�^���C �$X,���6=�o��q�
�L�����=OK(=����e����$*�:��;�=�t-���J=_N�������I�[�
=�8R;4��W��*4��	�5�z�����������=��ļ>P5=w]h=9%�<��T=�`�<��A�����#�=�]ļ�4<��h;�n	=>^=��{�~=�8>�D��j(�<�];�C/������t�=T�h��ے��(]=��<����3��xX=r�����=E=��\�� D��0{<��98Y(=&Y���� =��<�>\=4��<_'P=&3�<f_4=��'=tQ��tGL���Ǽz�G=�|��ݎ�<I�G��D���;�6��L.�����wD�<P=�y#�Pa`=a��<-���D�o�'E����B�.F��+R)��ē�H��5y �	�=��s<3L�=�d��m�=H���=Ѻ������0�=��l��xw=�;.�
<���B&=�S�<���i��;v�b=�<�cH=�15<��G=&<�,�T=���R�/=xdW=�J�s�ݼ6��<
])=�з<�w<������:�����)�<��g;�<1�1� {,�i����׼5��<�����z=w�N��4=-����ɵ���=�L��<?=ɎV�S�<�V8y=�a\��ɕ��~�;��P��z=�M�B����aS=��<`<�_�<����<����@$H��޻b�ɼ�h���=�]�<j�E;�_\�ɺ;�%p<�t�;�u�����c�;B�,=]�Y��cY����<���;�5;�����<=�B4��Z�O=ry=�m�<>=��S��^��W�;�.U���P�+��;��=�{=�C0<A �<t��<���<��G�Q�=}=ϟ.=s���F<��㼉Y�<��<���Ɋ��	n�ۋN����T��<o?V����8i�<�6l=4;e�gJ����Z�<Jk=�i���t�9>o���Ԟ��x��bYE;d|��&��<�������ie3�ۅ�;��<�p����E<T�<a_<�!=�*I��] =��$=�V��=hΆ��&3��bE<�S��F���:=�����l�����V�+�&ļ"�<��H=����j���f�����<�I/<�H��Jz=�����r�U<r����Q<"��;�]�;�n$�q�Z=5�v�F��;_`�I2���O,��=��%�l�����<������ܼ��Ҽ��:GU=�U;��"=�OG=!,ϼm=�=���<�\�iW=� ,�(3� �	�e�
<���<e�w;���\=ؓ�<���<f�V=Z%�;�g���*��bx=lU���A='��A8*�\�Dм����)��0�<y�<=(�:&�ۻu8C�����pH=�����|���"=���<�y<cۻ�\=�mE:�.=7� ������<5��;�ܧ;eH�;[["=EQ=�zO�_�<~�8=C��<�7��c���*����h��;g4�<�oY���ϼ(X�
�8�ީݻ=n��kx'=i�%<�2�� ڼ��;��]���=?-���%�uۺ�S(<<��];�<I�\8�<'�+��<�*= %�;Hֈ<�&��=+X�u�@=	�3=U�6=�e�<��N=JF�����<LrP�$���*2e<���:�K=��R�� =�,Z�:�:O���"��j�<�:�f���ü�=�D�=O=E.������ā�����!��#����j:»��;K��3=<3
�92���M=�/=ۍ�<M:/�ߠX����<c�N��C�<Iol�P�c�O@��2�μn4<�� =�Xv��X߼��+<?xD=x���=#�a��?�<-�R�K�9��ἁ�^�p�<>/�h_����<����m<{�0=�l=w�=�I�<ܩQ<M51�a��ڑ>;$E���k=x�껶�/��L�<�̼=+�<S�]=�jX=񭒻�] =�k����<
kU�O���!=tF��&���4j=6�g�M�
����<`@;�V=M���<���<�pm��mY�>P6�t�[=��U=֬W=��v<�����e=Izy=/�¼��&=E���-�<-[�����<�	�����
)�Ί�<���[�y<���J�'���;��I�X��=����ļ[�<��A=��C�7E��G<7s�s�;�'�;��*��H�&μ����٨�~�$=;8=�P<I�����;
<���(��+�6=sAH��=�����$��@=v?=���<O3t<o���-���QK=�+<�9c=:Ds=S���[�Jm�LN`=wH=pa���>g=|D=�)��J&=O_�<��B<_hh�� �/�3�Ņ�<�Im<w�ټ|c��O�=�R�<�5���5�a�<t�C=�2=隶���`;Q	�9l�=�K=[�'�D/,��+<7.���8����n��<�Y�<$5=�<<�)f=HZ�<l�<�[���=t�<'����U'��	=�`�<�M���L+=�q�<l�q=~�\�7���.��6�H���<H:�O k��kU=9�<Pk���/-<��;���:�d���	;�|�;x�<��c=ܭ���k-������1=�`!��-�դA�D�7���f;�<W;��=�_�BqV�4�A%����Bs�Vś<�/h<L�m�E�9�c�k;G�;���������ںC~��];<��G<�i�<V�(�fo�6��;wrY�@�+=��-<�oL<#�������$=m?���=94缁�:�;:=
�7��;;�=&n�Gh�<���q}�������H��n<n����q�$5E�����(�U=^p����<-�<�D���z�rp���O�ѣ�<�<2��Q����;-�O=��*=��C=H\9<)�8���޼�ǝ� �*;� ��ZC�}h� �����#� M�-�:����G�	�FE���e=qP�J�G��(=�J�=�!I=���<l�;8���HH�[#�81#�C|ϻ�=�;=�$4=�ٲ�8Պ�dc���&���.��v}T��T=�
=�4��F��m�9���<=���<�μ{�;r=`=m,Z��x��+E���0�X/�:W5�<�4[=�t��aի�E�C��'�<<�=֨5=��<,~�<��w<�Iz<lL�<��!�}�4=S@<��[��.f�<� ��j����=�!L���|<����L�T�<�n��^=t�����:�L��P�<�lu�3�� ���jH��h��n]�����ފ=̰�r���2�]�us�;�J\<��C����<�'�<���=�+%=�g�ϕC<2=td�<�r߻F�<F��<�4m��=<ݜ�;;k=]q��,����d=l\(;��<Y�,�������6ڻRc/��eu�3R=��=`�������l���� ��p<Od��w�<�ԼG3,=�ݼ�*%��?e=\Z=^�����<�
d��Z��k��<u���D�}<����;�n=$h<��|=��͐=K_�<��G�F���஼���<��7<8+n9@�e<��=Az�;U����<"�b�N?9Z�<**��g-A�6���5=��,<U��b����<�
I�|�o��<�L�5N	<O�Ѽ�-�<�&�����F�<�Ｄ�h��L��4dJ��L*� �.=�T�<�R�)�<��G����<��L����<%=w��ߎ�噘<q��<�OL<?��:��:=��-��;
��~<w�7=��&�V�[���:�u�<��
7=��!=��=�W��[ߌ<�+*�)��=��c�<�-��8�V��;��=?�= ȼ��;Qc̼�ѓ�º��T���+��/�}j=\��vW=�1$=K�7��f�<'J�<���<D�=����Y=�>r��K���
m�"�$=0�`=�-Y�&����_��{<�<
=���<�@=�L���i�;|1=���ބJ��<��m��Լ��߼�)�<b~�ˑ�<���<�,2=$,\�'g<v>Ի��I�Y��<I�����To/<OI=4��<�P��̼O�j��pZ���<�:�<�=��2�?�t�%]����:<��J��2:<�S!���C��e�,�={<G=L'ͼ
=��o�;\Ԗ�]��<��,����<�8�<kyɼg��=� #�U;"�=x�=��	a=�C�;
��<�Z�q��������$;�$�9��D��(��~��4�2�)=B�z�pU�<7{�<���?��<��c��wM�=;&�G�P��]Y=�w����F�V��<�N�{V�<Fnk�
�z]�v�!��=Ӌ�;���<�,	<)�C=������<\P��:5=pG�E��V*���4=SʼOH�;Ϭ���Vo<[ �<{�<��@=x"=���:��=���<=<�<c��������3�m��<���;OG=c��<�.���U=���<�!���k��t���=�E>=�N:�s:"=
�i���ͼ�%F���=[(3=Z��<��#�Zc�<-�>� Z��&ļ��l<�;?���k==j�V=PG�зͼ~D�:G5�=\���C�����:�ż��;Ⱦ�<%��U�U���<�I<=I{�; Jw=��5=N5b=5Aټ�
�<"���v�;b%��È�q{=�p$;����"=�P��4"C=S�/����<VVL=�0�ƨ/=���Y
=3�=)��<�r���R�<��<!�b&=��!<�ҋ;�2 =L�"=��ջbxT<ˠ
�K4�)�(3����ȹs�j=]G���<P՛;��ؼzɨ�VES�Pfg��,�Dm�<���^�׼k�}���Ի�&=��<��r^��Ug=Q����邼��<�h�<<��©�/�(=��=�+v;�i�<�T�k�Ҽ$��<�@�:Iqt=c�h�N�\��=͔�:�k=3`A��:8=]
�&�<�=�<����[=;�Ҽ�9=�:3=�Y��0�3<A����	<|�A=��!��R#=8�b=�H���=�)=He=z===}��d'�;�B=��e;���<r4(=�����|�c�� ;$~<��{�i.�	�b=�g=�U��C=��ܼ��.�nu�<��=����<܍B���;a3���$=.̼�4=i\=]��<��＿ѐ�6I ��]Ѽ���Hhj��cܼ�b�<�y<N�Ҽ0G���<�f�����vK ���=",�_�5=�
;=r'���.<C��<)�<d7A=�P�<��i�G=�u&��|-=��<�T;ݱf==J���<����R��;��R�<�ü��Z�+H�;����ˈ���'=���g#�<�.Z��Y�9T�Z�#߹<�	�;w��<�:��Ë>=��(=� ��Ua= >N�2�y<XvM�r���F�k�5Rȼ��2� r���8ǼE�I=�,���qE=Y�;���/Q�<H+�e�'�y�3=�m��~�=��`�-�i<z�3=Cֆ<B�;=�^U���H=��?�}N����=�|�ac��N��ܱ�<�мG+^=��L���\������K=˛� ����+���`=��3��;��;<�?�R!�<�v�<�m��q���� )=8J<���3�= ��[3��� �yl=�o8=̶�<��)�O}(��m߼���<QI`:h��g�<OK`��9'�(���nw�;QA�:��.;/G�j)��Y��]��<$6ּA��<�I���k�=3�<�+����I7e��``���<�Ȅ<X��<�1X=k�<`�A:�M���l<|�%�wG��q~)���@=5XJ�1B�<������=����}ǼQ����*˻޶k=�w��ŀ6<Y4=��v��r`�#���hZ�<!�H��
=�<��R��zM=ƚK<��<6�"=�΢<~XT�kR̼� �	��<3�?=��'=�3�������=�\�<��AF�t�����X��=�^�;��=�����Fo=��-�;Z�<A�ռ�*^=�z]<d��@��:��n�:I�:=�<�e,<�݇�{�\���+;��T<�>�<�J|���Ҽc�6=*���i���.t#��aܼ���}	�w+u�9�<���<A΁�>7	=)�<�<r�9=v��#��o���]�:,�3�"r�;�� ǿ<`����!�ȼ����=�<����&�<*���=��H<��@�Aj�]�<���ݿ<x�*�b�=y#����<UL_=��%=$�p<�!#��g���}A����3�cq4=lo"�TT<H��<
Y<=��=E%��n|\=EU�=�'�9fU�<�Ǽ82=�=8=㏍=-�q=��(=�� ���<.
��E$���=���k�3� �$��<���=�~{��9���H<!�<<����7 �Q� oC�je	�P=��=�-7��ө<�케2<��r��Ϸ*<�'��y�<�)":<c+=Lk��e<���q 2���+��ִ����_��&=��A�GN=�<=rK�B�g<���<���`f�<��<J���:��[��&��%t��D ��E!�R3A���	�$�U4�V�X=�M~�lC�@�h=e]r���8=�/�Ǵb�J�x�=��L.ܺr����;���<R}Ǽ�>���~=9%�fA�<���7�|��=�&��p5�J]���"P<^:м|� <�|]=J<=�v��=r2<L���">�[����<��!=�HG=�'=��.�[�ڼ	!A�,�4=6�<���[�t=��O=-�=���޼?4�<#�|��5<I��D�D=�/�;zJ=ܧ�<���;��/��������.�=�<�q���=]�z��JN��l���%9��ڻV��;1^�:�7�<v�8=�J��/��Gnb<��f�?�=%�ɼZ̷:^��<�!D�}M-=F���*��&�I]=��=/��<��Q�,�f�t"��&����L=ч�?��<Ό,��\i=��i�F=��¼̋�<�i��8�<}\=�/�<�<��r��<�ױ<p�O<
ɖ<�<�,=��K<N �<y�ټ%.�<�~=��;�{N�y],��R�<:�Y=z��:�J=
�3=�sq=�$e;�.��d�L���P��L}<t�=��"=H2=#=��<x���5��<�
=�s-<{^�5S�<f/���8;�p�I��&��yq���5��=D�Xyۼ�b=N�<_�#=�uD<=�n��G�r�����ּq�;��<`�����1T�����C��?M%�E�v={�ܼ::=�ϖ����;uz=�����<�1�<�￺q���F<�N�oH�<���3Z��7=�W��Z=@O!=5�E=Vb��`�<��<$��<6{�<�:n=.`�J0z<��#=U �������<�w�==�%�̋Լ1I=���VN�a�<�<���<no'�q3;ϡT=�a�<z}=�Cw=������;4�5�A�WKA�'=��Ż''4���T=�8 �1�h<�q�=u�o=�B�kg=���<�M�<���<�x��DH�[�H<U�C<.�7=X�6��;!==�5=�1#�+���σ���=�%=�4��u��<�5�<���^'2�hF��w��[Y�B*=D�:ns�<��!���2��J�<�U���z�I��
�@=���<���"�=��';0�W�Q-��!A<B�V=�k"=�Լ0
O��Ԭ:���<7b.��8=UpY��h����y<.�;>RB�������w(A=�9�<
.S�3�,�;̼^�]��V��^1�<�ğ�ыs<^�S����������==�ؼ�<W�<-��1�=�*�<����e/�pWc<�༪n��֧.=\�l�i�E��:)C<=q�;��������ҳ��@O	���A=!~�<��9(h��,%^=������2�|�_=��1�R�>�zS�;��»%������<���صM�C=�=�)c=�U{=6;=X�+�u�]=�YN�����P��vyO<�,޻9�F� R�\�*=��h=��<�#�<��$<������Z%=�Jm=�wC=��2�qO��9���Y=�qk=V��@_B=\V��.V�c	=~�6<Mp=y�=M�|=
-.=��Sq =���<�S=��8=�A�J�����<��=�<B��ڼ�X<`���=��<��;�6r:6M�gq���.�<!�(=-֘<,%���G<=�(��,�_n=��l=E�+�&�@�o��<�)=>z�8���	h?=>��<%��<��B�˽�`~����ٻ��\<��~<�Z»�~{���� ��<�1==�lg���d=6kۼ��-=��/f�X��)Nw=�^a�ӑ���bl���1�o�2=9L=��h<A1ʼ��X��A.�d1<�8�=�3ټ ���5���?z�P}H�~��|��<A�3��vO��
�;�
�/мX����E����ٸ<?�U���==ж˼R�2�m-+��/A;e�l<�� =Q�@�H|J<�|�[�����<+����e}���"l	�^���\ݼ1����V>=3V��^�<�3�����nx�V�I�L��Et1��=�==lQ�;�o����5=�2=Y�<��м	��}K���=P4=2�<\Q�=��c<�8#<�˩�GA=Y+M�z'=)��<�l9(�7=�P<�N�;��=��K<�[��D�9IQ�R��; I[�
>y�W�Ѽ_��;�L-=1�@���u���#�\x��.)1<��>����J<ަ޺{O���d=/���(A����B�P]=gJ��t��<�==&a=}ߢ��,<�$,=�@�z��7�
��[;�*�<��߼-S�<�B�<�$_�5*6�^FK�j�&�l�d;?�?=��'=�ĭ;'������G��;2���xr���ܼK/��M��)1=�N!=Y�=p"=��(=��a�ް��C��<�s=��'�<�3@<�@"=Պ��m��F���3�<��b<���<	_=UtG����#���p=�33=��=AD�7?��N �:��<�*�G��sB?<q�=akw<��s=�_�;p��FԄ�p}"=�g����<�!y�/0G�6�i=�	h=6P=�h�=1�J=A&�<��qN|=�S��IR�tS��t�����<1:U=��K���H�>c<��N�������s�{T�7=^�;;q�<,����;�	�<�8��|@=]�<��%��\<=n��D�<�N����<i�$�Pe\���!;�+@���0=W���HAT=J}��1�s)��~5�=��<m�	)7�=��<��	�
m<�G�����<V_2������=�xM��j�<��N=��ܼ3����9��/���ͺ���<lQ=�M�=�~���# �1$�<�Re�b����Ҕ<?N	:�/=�=ڭ ��u:��ڼ`����<=��0�+P㼿6$�+�����;v P=��'=ȉ�<W���Z��� S�;&�����]�y���
�]<���U��:�	���=�wμC:���ڼ ��9q� �d&��p� <�����<~�����f�f���f���Y� D�t�<8�d��7�;�~�<�D���JQ��1�*¼�=����z�!�J�<�1�=����R6=�b$<Ɛ����;�]%����������p'<;�f=�=��%<��?=��8=d֒��^��~���5==���ćn��l~�7F���]��@ ;��L��\<��v��lk<�G��$:=
uG��v"=c��� :s��bb=���<� =(^�<�#���EN=�k:���;e��c^5�K,=�>�;Qc@�NQ���@�{��<0�"�~�\=�+�:wx=X(�ƞ�<��R�9�I=!�J���9<|<uc ="ջ7?<�d=�u�<�<���T=�(=�3�<2(�,/;�E�h<��Kd��O&=�*)�W={�/=��!��F*=�!x��,=ՒW�F)�X�����"\z�cK�x�ȼ�����9v��AV<�>s�N2�<�(=��ʼ���<3�.=ŊI=��g=�	=�}1=O�<d���;���<�i=+����Ҕ�sjc�1�߼s�=� i���h=l2�;��<���<�Dټ]H�;ֿ=�);0�'=P�7�}?����<��+=�\����<�M�𭶼?]+�Rx<��J�Xm<;%9=P�g=0�>=a2���d�< 0e�TY �	�'=�� �ӯ�<:B=I��<�>�<����?<�}=�~j�0Y�<%�=f��o&x=?���d;�<��:�j�K��<»0<�\a�����<5��'��<�}O�B
���q=_�^����;a�<%�1����;B��P!=������2�O��¤K���;=�`��]4s=�8C=��<��=�BU=�Y;�0�=>y=��o���󼹰#=4��<Lhf�+�2=#=��_������T<�5=�"���� =;<sd��A. �Q�<��F=�I�:�w��&Ӽ�n�<��;��Z���<<[��������=�U�<u��}̶<�<=�<^�|<|	+�l�==���;�h�<s����bf��u�������<B���j�&=�'�<�N=�̼����A�GH=}�<������7=�*=K8��~��;� �<7t��<C�K=ĝ,=��E�Tq �n�g<�U��#W=f�2 �;v5%����<�H=ᾫ;���<�L=3<=�8K=����XK��z;=A�j������=�c=�;T=�>@<&�ѻ�pɻf�h�A����T=@wY�{5=8D�w[=¡��S̼�8�i|#�V�1��'뼰+�<�^����@�Kz��$f�(���1o<P��<LP���<��9��s��'+=ɲ^����<*k'=��$=�P�<<�C�5�?=Kr��cX�C���:e���=�+=����݃:=���]%=ML<�ӹռ ���C=�4�:��<>�<X����R=/G��/=��=�-ͻ����[��<� =*!2;�iB���h�iQH��,�;�����ӭ��<�)=<�^=Z�l<��@�SZo;�s����޼�?��^<�/]�vY��ZE;b���><��U�{7=fE<�ǲ��7�;��J�W��xֻOuE��7���=�
�:`�^=cN��vF��s�<t��\+�;���<��;@���������7K0=uP�=Rdz���-=�U.=~���R2��Յ<�D=l<�X�<�ȃ;�����?<�� =�r��Zs=hmO=[3�=/���$��B���If=�F/=g��^�!=Yn=��Q=��<�i_��h,�lc�:#���ͦ�6�_=�� =�bG=.MC=X��x�<뿥�t���c�g:Qf��3缯9��!мc���=v=3� =���aһ�0=�����Bn=g5����F�;��V�<`����~�< TP�d3��$�<@R<�(w!=�����e=�ӹ�����	뤼S �<�TK=��Z�����Q�R�[cQ�F�nf;�w�n��9=�*#=���<9* �x�}���<��U�ـ�<�J=�u��p����G��]g;<D���<E�;=S%�����q�������<'�;.���c=r�C��u�9^���0��K=j=��T�˸�<Qļ�Dc=��4���<��R��3���=òU<�m�;p5R=üZ����|:��b����/<�+07����<�s�8q?	=��?<����4ؼ��4=�h}�{�t�;jD={�h=�L2�Ɖ\��.=�7G�n�:XNw<&�4=Zb=tP����?��Ƌ<O`M�	^�;�uB�a4���=CY�z�UK	��B�=4	�`FĻ軡�=b ;��V�x�h=륝<�؆�Ҟh��/=�*�<��Z<�`�=ۑ����r��(�<(����h�<�Pa���'=i�<�=h=� :=q�k�yJ�9bZ<�4�;���o���=�r��v2���;D����w=>�=!Br���K�AJ=������Qh��������!c���;����#.�p�/���5=ZP���� <�;<�d-<H�I�q�:)�<=g�+�?ԟ��;���d�g���?:g�
��	=��R�]���2=��a��X����a�3�EU�<#ʻ��غ$�<��m=Y��=�3g=iĩ�I/=���<5�E=�C�@=�N���fD���Z=ޛ��̈́���!�5�B�A$Q��W�>��<d�A��M�;���]�:*�<��D=J����J]�t�(�N��;6�d���Y��9<	^9����8Ɖ;�k9<az���=]��<�vg��w�=}�q={M�����<?�W���=��/���<.%<ZĬ�S���yҼrTw;�CN�t/<~��<��=��;�=�U#<�<��J�;��<==9R��- �'�ܼ|�_=�Z�=�8�:�1��>=��+=����d1(���=�� =_ǻ�=�$=g"=�=xOH=8ͬ�x0�=x9';;�=���)ʠ;gD�xܓ<�̓<�7p<�;=�y�,kn��R�T�M=4(<���0�N�@<�>�<KF�<_A�� y?���8=O�ռX����%��(��HFd�����Cmd=�.\�QK-���<��i< 
j=�<��ۏR�ItM=C�9�_i���i=��<i]�<��%=�=�����E(�Tp�����F��w��<���WDo�NTB<��j��E�8�2=5�|���	��s�<V��;���)= ><f&;�~�<�R=�ź<a�
�<�=�3��[f��ϣ�^�85�����};$m��"L_<p=�l�M��ϓ<�&o�$���<	|=U�>�_x�<"�@=���zz����<�ݖ�<ؙt<�dD�w�J��#Լ��O=���;Sb=7�v��:<�Ƈ=�L~��'��1ֹ}!1<ޣ;N/
=V4&�)���uM�z���Tp�<\҉��D=��<;��ְV=ؗ_��mi=�J=�X=�Β=�=r��y�3���<=A�{��^=,~���:V;��=��G=������$��D༌7���5�����R��e�����;���q=P�j<�	I�(���E��B�=���<EM�g=@����p<��,= �=x��vϼk�=y��;��;���`�]����g�}<3�<�]�;��?��g?��;��;��ͼ�z���s�<�xҼɂq<G:=)�=l���N�ʼ/�C�=<�:���~ll:��(�����?uU���@�YGL�m���S�=�+� b=�����Y�V��dC�z?6�(�:��R<�~���d�]����6��<�c�=� ;u��\HO�����N�<�:��T8<�ZI�ь�;�~�c�H��<�}��!5<�����;�-t�J�=��
��0�<�sb��1<�N<�����=�4�Jk<�a�<M�0�3R�a��;8���<u�ӼWM���<~�\�
#2������5����<����p=���<.̼)1N=�_4�n =K�<?Y���Fu�]��;��<[^�<��z<T.-;
G=j���ق~�,[��W�G;��:�*�;�<Ϩg��@.<*-g�@�b=�)�;}(O=:�ʻ*�<�p˼��q�<R�;�$��*��ka��k;=z	<Js�< �=�|�Ly<n�_=��ż��K��#�	)5<���'w�<N~���A�����"��Y ��+=H�꼊,e��iۻ���<�p=��q�L=NtL��Z�����q�-��ϻfܐ<��dVD�J뼧�\��k <I�-�2E��炓<��2<{l|�����S�Ց=lFU�K�k=t�*=رF=�J=��l=/B���~��g�<F�*=#��_<�o�q/�s>]=Y�_���<;<�<y��^�2=�Ww=��`�x�K�<�=a%Y��O�<Zց��<b��d���B�.=�<*Ȍ��ї��	�<[��<��<��X=�V=�L= "5=R�t��� ��=�Y'�qx��%A=��+;]��<�|-�rGP�� μI阻`��Α
<�Cr<�ќ�m�=4�^=(�G�P��<���ļ+#N=M� �*�=�������D�`�;;Be;������< ��<�eR=�8�=(|�< c|��p<��=ʴ��y��;�҄���C=��6=�(<�F�k�+=t�
=O*�<�:�<4t��:N��!���{2�r��<��=�K"���V=�:�*�<��f���i��H=)����|�^=��'��P���K�K]B�l+z���;W�+=!�A=|)o=��L�GG�R<1RP������K=no�<����n��=l�칝p�<��f=�,�8q	�'�a���:���`�f�L<c"S=�����뙻��]<Ki��U4�Tq�<�H�;N��<��<���\��7A��9���:<˔u�'~���!�8=�Rּ���6 7=���<��B�<.ּ%�Իs4��B=�����خ�C���E���	<TZ�;?f�=�  =?Q=m,a����<O)C��Ҽ%�&=�{`<v�ʻ`�ʻ[o�<޼4����9������~<�r��"���m=�`�<am�;�N��Q�:Ub1<"����w=q��=:@���+�;!����+s=C�s���ż"�f��7r= ��!7;>���>[L���=&�v�<�_�E�=�S�[��.�=��'��ӽ<��<��	�w�n�؏�<p�<q���u�;�q<K�f;b�=i�*=�=�#x:� =h=�GL<���݀�*�i<�J�=�4Y�pA�<��o�=�=v�,���J=Ȍ:.�=��<1�H=�C�<�us=�� �̎=<�0E<���ݹS�	�b�KI��vj=,A=�7S��T����;&�=͉ü	�2�r3B�G�l��=��H=5_��4�=�%L�<|q=�L��}=�*N=���<)Zݼ(̪��*���)=Xx�qY=R�@���<��*��!C���=TED<(�޼�ټ��=t���@�;]i)=s值<�����k�d�*���D=�m\<!|9=Em��*RQ=X���o�f�}����;$>u<GG�<�S�;%xż���<Tv4�Rm=�h�<-�4<�:�<]�<�#;�r�ļ��<�6��|uS=`pL�����=������[<���<X�Լ��Ԟ�G�Ӽ��z=�qw��/=�}��:�L���X�_�q=�4��a<z�9=	�˻C��<��v㚼�v�ݏ�G	=���/��<�`=��p=|c=_</<-m�<�r��Β˼ڿ	=��S=�ch=m�U� ]=����l��}��i�<z�P=�<<#ɻ. (�x#<��=v����:J�O�l�==�Hb=E�2�@}'=�]6=H)E=�D}�L|���)�3l�<��O�����n+�jz�;\/�;�_�<�:=�\Q<��<�:�~1==R��<T�a<=���hN=%3�<�q�B��:c���-C��o���p=n�=�O��h�:	[��v�����>�dwA=СL=�j9:�.W;�g���K=��b�q���0��<�Œ������5��y��;��#=Z+�aI�<?�a"=ݓ=�:%=_N���=@���(���`=$���p�|���4�wP� �Eo#�rj#�%L��h���T?���;~Y=]��Z�'=���4*=4z�9<P9=�Y<�~�����<�0<�F?��]G='��<|�)�5�N=�O��!�N=�����0=(J���f$�$VG=���H�<5�;��y=T=x��<B�<�u;S�>=�_<=J&�<�6���0=��)=Q�+�4��/���y�=:&	�Xb���+<[�4�&V�<?�L�-��<'z=��R=��K��b�����h�2=��-=���<��<�3X���z;���<�4�9�,=��ۼoQ,�(�=���k=��g=k�=똹������5�a�߼���s4�<T�f��h	���:=T	X=��A�xp*��V)�$�p<�=�gׂ��<�d=L����d<�;Jdw<�?=x+=��<�ZջJ��<W�=�R\��᥼O6�p/ �U@t;P']=Hܼ�=-7�d�=�Ga=6���̤��ՠ��|z=�㯼��<��=J)����hɺ<1�=������I=�~�<�c�6}=b��;�� ���<�?*��2=X��<��><���;����ǋ�C˃�ꟻ㐃�͡=���V�b{=TԺ�/���I�<���<��u;�n;��U�Ӻۼ��:�#���k�D��<O�|�
��<��2<'t<���E=8z�<2ɋ�h�E����Ϥ��%�<�wټ �-���<O�I�;P�w9X=�>~<���;��B�h��<
\�<�i����[=�����d��|/��~ӫ<L�p�;���"��E���'��H���9y<�L =�Ɓ��NX<;Ɛ=�"��$n�h31=�Y�<5`<=,�;��m<�47<�/��R��<4��<��]=>]��੉�J���]
<�1�mZ�;+lM=��<���E���(�t�ϼ�4d=��D=(��<��ür�C=��;���<L��5��������=��=}���1��R���7=����A?9>K=fi ��� �I��{Y������ݼ��0���8��9\=t��;_k:=��<��w�_���X-/�7�)���9=@|�Xu;�I��+jӼ�\Y�a�<�3Ҽ��9�򠼝��<UE\�`����s��vc�z�U��i�<�,ܼC����1���o����<bJ�;:������;Q&�N۽�n���Y=��>=�%����( �Z��b�;�z��5�����=Db[;u3s=�Y/<Q�D=��̻\)�<�����@��D ���D���=J�a=6Y��f=p�L;ؕ�d�]�}�4;VZ�<ta���O���+=]�.����y���n�8=���<V� ��K�<��=��<�û��y(���w��Z�;Qv��Ee��]�>�eG<�z�<���;B×�s�u��0��X�<�F=�,�Cs=��O<��/=��=:q��]�)�^�a=I�<��Q� ӻ��l��e�%wt=w!=|��<�d=9m=q�8<LUb�R��=���<k(V=eH�:��^=�/=~s<�w��:<��=���<�0�<�M=`��<;�=u����<�㹼|"o=
\，{C�5�8<�&=x.H��=�>=����UnV�*70=t%f��r�{@=�T�͚Y�OM��
k.=0�<�"=���P;n��:ۤ`=|�9=�o�<8F=H>N=��:�������j�Z��<�gO=�9b�,���VH�7rHA=m,=F埻�~�<��<�5U�Y�<��;m��<�R<"�3��Rr<8p�����<�����	�Nʡ<����3+=��%����'��i7�� �����<��X����������)���#=�,=�:��<kxg�ovL=�=F=}:];�nؼz�:��#�cP=D�O<�Ck<ך:��!;��a+���<=7Y<�)<��<�=��;�&=�j!���R�x�=� =�M[���a<&'=4�<��F����<��0=��=�ǿ�7A=ں�}j��ʊ�\�=���:G&�<#���Q�����|z�Ƃ��픻����3�4�%���<1��<�s<&��<��jU<5�C;'پ�=J0Z;�m�=�`?<�-u�u���2E=G="=�+ =�#��h90=u��<�NU<�(>;<�m��;��<g"=��Ъ����C�F\:���!=r��<��<
�<
T���̼p�P���/�˛�<�*��l�<����va�$��;��ܫ)=�;���r5�X�=Ep�=d6=a��;f�S�m=b��<�Vd<����^��d>�Ʈ<=�q�N�`���;�A�<�X9=�=��.�zt;�<V+�R61���;�Q��w�B�<=�)�4X��[�-z;=�d1<ތ�; y=
�G����"ʋ��A�<�N�E9o�1�<�,�!`���μ{�����=�Έ���<�\=;�;?{^=��B=[+=`�h=ﺻ��Y�_�<(`B=.���R<a�̦�d�j��(=�c<�@=�����&�V+�	�"=�%�;߇=tk
<�Cb�� ���R=�Lϼ���<�۫��w6�\�׼$��<�J>:	tm�C�S<�F��#�<����$�{��<vS'��p)�^lY<p��<{�<������:�47=	�;�*����<nd�`s��
<S^�<�E=���=sӼ�/�����.��H�<���;��\=�˰��U�VӼ-�<k:� q�<�蟻���<R�l���"�#�ּ��==`�&���<���;�oż�=���<¬a�z�*=�?<���<�'W=�μ�-W=1�4�m�&�=�1�|�U�Z�����f�â<�7<�O��ɡ�<��N=�r�'c��ژ�O��;�E�p@6<(��<@���]�H��v��&��<��!<�
ƻ(6=�f=��*�!�\��x�kgm;��<�տ<[��<�n�����~���hV�и���b�<˃�mE���8�</ĕ���μ��<�CP=�w�<H׍�-�?=G:��m+=�xH�[�6<�Q��E�t�5�<�.E�'s�[İ���^���R=�O��J����.<�`Ƽ��<O�J�wU��Ad�A�'�Z�=:_6�|�-<�=��MT=��;84<��N=�r;�2Y����>�'�������;��<@���;��y��Y�/�;�1�<J�|< �)��P<�_ۺ�2��c�<�:s=�9q��;�e=˪T=[��<E�黙���bd���P=>̉�[R��V2="�n�X��<���c)׻j��>����G���<�7=5
�<A#��UE��ͅ�0��;�J!�tQ��y�;��>=����7+��M����Y����<�����Z=��;�=�<�'�<�%�<K<�3�8ң��쾼��9��&ػ7}h=>�ü���L�|=�?k�����DZ=/7<�-*���P��;�y���u=1z�oU�ML7=d�<��=0Z*<sG�����=[�T=�����)��ʶ�m�G�)�<ʞ���s���<��l<�Tϻ�
.���=��<���/�e�;�����<�G=aA��}��o.<���y�};ڣ��Ͳ�;.����鼆�f<۴��=���<��"��u9=�z<L݁�>�����E.�<�#���@n;yB�<x�X=m���)�<�)=�Z�;#���4�9=��r=��<��=Q���)�ܼ��(=r�$�X�<5�D�s�='"=�=Y+��&�+= �;2�3�ۆP:�'<���<�Cq=�Ԫ�Bb�<<�X;���β�<�Y�,^{<#��;K�=�F�<���<�0�b�{;�/<�<���vܼ7T�<
"=�\=�-�OE�=�ݼ�����$=n7==ƏI=e�����<!�1�!��;� �;y�ͻx��_�����/��0o:�LI�������#=�b�|6*�B�@o��j�W<
�H���6�j�2=�KI=���9�i��}=x��'r=
�V���S=3|R<�:��J=�!F���; �Һ�p�#�Q=������Y�M�+����5!�=.^=���c�<�0��{���<8�뼦5<~�'����K�x=�D<�1m�3:��nc�('E=�K���<�`�<囻N�<=%�>Qo��{<��S��Ζ<��x=�=x`Q=��*=R��=�i�=ز�;���3�/=:<T����Ƽ-��<���<�(�VM=���<^���  J=�#=���<���OE<���<d�b=��a�xy��t��Y*�Q�K�S��<���<r-U��|�<U�N���`<��z<��+=U&s<+Ļ(a;�$�*�<�FW=:1=�J=�|_=ܸ&�"�ݼ`Q�챈��.�׏�x�R<� ���R��b�	�j�<à��L�!�l<��<�3���o��0��	���Ѽ�,�z�!���X���E������؃�6�'�I�9�0�<�J&=���b#��mH�yU�);�&�������=��<�"���׻�=C�����;�QX=��?=~�e<��s�����_��7w�;�N=M9��_������� =��<m[u=2ۻ(c���^5�֠<�D��W�:ĉ9='�'���;�D$�yzt�D_=a(*<֥�N?�F�{=Y�r���<M�=�=pny�$��<�R�<���<�'��꼯��<̋�$s=�^�<R�:{=$=V�DTT=aRQ<33����<���:o���|���M<k�0�b4��/�����Z=<��:�<
����V=���6T��%��Pn���[�1�b�h���ݼ�D'�4�R��y���<�g
����=I+?�9�F<u�-�:f��"S=�y~=Z~1�w�<�K��S�<sj4=�q,��}���S=9�<��(G���<�D��l=��;��<	)=Y��F �9M�;�A:*�;��H=�V��2��[z=Cq�<�o�f@�<q�<f7];,-a�RE��l�L�<�����Z�<	��<hϼ&dX<|,/:�D5<N����H��4=��<����#p��TA=h�ϻ\���p_=�J
=k?j���ļ�
�;2�R=GNi<��<���9?=�I2=2�U�=z���#�0�J=��<�U�<Xnp�	�/�E��<L��l�K=��˼9)=KWP��<A=x�Ǽ�ك�7C=v�(���&�'4<=��L=�W�ՇܼW7=����;L��Z �<[p�pm=�AN=�Ǝ;�]=P�C���y=h�=Wp��/�==LF=w�<<�;&��k�;3�d��;�����`=r#˼�1<08@��Ֆ<���;�[=���<
<N�R=K)e=e�j��H�����z�l� =��#���< .`��a�1� ���7���*��BI<�m	;�{���X���<=,�==�����:�5=��5�?E|�7v���fE=@=�c=��<��޼���<��m��r���W=�q"�,,d���K���@�"=��<<�<YE����=?&��~�=+=�DC������-��D��<t�"=$�����<AE0�Ԓ�K�;�G׼eF�%��;��k��NE<��ڼ�&�O�9������I�(B����r:?J ��W=�=KM^�� r����t�X;�F���N���%�U��P��<��v<���{�<m៼?m�<�uI�.=*��oB=�f�<r�S=6F޹oC� \=�\���D<SgȺ�F_=��)����q�;f	=�1=�@a<�m�<��R=ՔI=(�Q�� @���ȼ��3=��9=B��<r�6���_;�x��@�;<���Js�<k�o�x�}�<�<����;x=��,= 
=����;<E$�'W�;B�;����U�(=9u̼r��\wY��1�<8�Ѽ늟�<��<;Y�<��<Gῼ�+�<l3��
C�-����<=�W���#=�==j�<L������I^=�ʼq�=B滼�LK=��<�У<c?��?t�<�=�vܼ6굼J�,����<p4�<z� ����"�0�\�g=QV�	`�<w��<��<�d���=�[N=�
�F��<4���v@<��:��D=g<��?��c=Z5#��ys�vW��>��Gjv=�i;�	�;�� =��
��8�:�=ւ���%�=|$=5v�C�L=�/�<l�]<��<��@<$�%;��=,��<�$��w�<�߻��v=�.ü@�'��1X����:M�=����Wً�4h=��"=3e=�&h��Jf��`ּ��B�f9F=�E=�L���C=~��<����C����*���=�Z=�l5�� �8ں�N;B����0�^�1���]��<�-<��H<���d�S=��k
����`�m=��:�Vt=�c<�<�D�=�}��Eм�Q1���B=�9�]	>�G(��?�A=>�@=T�
�׼������<��<��缢P@�[8=^�#�5��;�伉vZ=}�=�<�������M��1=��l<��<�`��<��<��!��8�E>��9`=�rF=l����M�S)��Ys���Â�-��:o�!;��q�O`����2=8�
��a��=��o���/=�@_�{�<(O�`�;��+���,=��5=j�|���p�Mg�#����&�����<'!=��#=�<=�1"=�L=�ʮ<�J���%���;����������<�d���:=���:��;c�Z��=����=o,=J?y;�=r���\���D1�Ɠۺ����D@���z;D����cA�T0�;3�n�� �<&*a=H?<!�+���<4��)���%<0��6�Ǽ�Q�����<�@�;�:9��2��wV=yf=�輇8=P0=₍<�^ȼ�`;i�U=�v<���;���<E&K�Qr��م=
J�^�#����<�D��S�<��=
�V��j6�u?;�)�=�u�����w��;���<�r��P<XGG��������@�;� A=f��<�;����=qk@���=�P=|� =��}=���ҁ�*'�;�(=\�:h��)�*�����9�%�q��ҼE�ռ	%=󴦻�;��/=�g������+%���;sܼ̍t�HD=8f˼��<�����W��1^�
j�`!�<5��<�`K�B����M�K*���@<��j=&JD=��c�e2=�~����<Z+��-�<�!뼢�h=0>�<��ӻ��F����6���[=��[� �ﻳ��<}֟<�7=������.>g�v=4��â�U�J�U�(=?�=�,�O��N!A=���<�<��`:~���Ɵ�uTN=���<Jl\�ݘ�ћx=�W=kG��R�<����H�b�A<�r#��22�#�{=KD��(���< ��<Eʐ<���s =6ZJ���ϼ��&#�<�� �#�,=�<=Ï�<_�M�d< փ<������:�p�<w��<X��<�<��N�a#���<�b�pA��T=f7[;u���1n=����e�=Y��]7�:Oɼ% �<R�̼��Z=�e=!m��0ռ��ݼ�`�<m�Q=��뼽ʩ;�c(����<d�.=�i�'����o��(= X�<��	kr=�?Ȼ|A=C�C��<�.��BX =c�3�`�u�\B<o	�<5FK=��Ik��5W�I��<�^��#W=��=�,���n<w]=ς#=�V�ω[;۟<|��=�#Q=ׅ=�e�<��x<G��;̈漲�)<uA����u=��<�h�P�{���:=��$��7Y=��T<�*���B�B���{�<�'<����xB=�g��a�B�<��<d�:=bXh=Jk�9�R=+�˻*���rR<�3�<���!��$�j��=b�
���F;��=��_=��6=aa��=�6K���<�킽ǜA<�<��ηֻ=s<���<�R󻸂?;��k=بǼޠ&�\N���l�=�5�<P<���^I=y�^���=�콼a�ؼ��L=̬h<�=�<W�=􁽖�3�s�:kA�;�Q=oO�<(�
��04=M6�<~�=���<rj�<�h�;Ն@�>a;�*c�*�<4�F�=���Wp=sH𼞫ٺ�;e=���<L��<Ve{=��[�ܿ�<@�<v�;�����e=��(�X-�<��ʼd\=�����(<9�n��L���;�[��p'`�����+�=�9�<��E�Y�/=��$=�&�<�L�=x<��8���,=&B�gG;��ؼ7!<�[)�M��;SI�7���е<�}�̵x: ߼���<h�;v�{<�#��FB��}��{*)�E�=ǆk�gRn��(�=$=����)�b�hj<�K=U�=&�h<?)�0}�<\W����;ۧJ�t�X8�m��p����&��:=s��#4���=�����}�<~�=��əu<*9�Ӫ��X5�<𛊽-:S�0��J�4=�E�<����X��<T�v<�O�,��g$��=,=m8��o��΁b��Y$�z�g<M�?;��"��̸��f_�A<�[�u=w��;�=�=$+���3=d7b�2j<*�<��V=�)�<��R��/C=`���vD0:t��<?Ә�c�;�B�nl��9��c<�3�ļ�mQ�|up;cꆽ��!=�	=��9^�:��=ԞY�+�;É��n=������<�@#���<Z�o��໼i��<��h�1�o�C��<x4�4vS�@\= d�����Q<=B$=�e=<Z==�<W�<��C=�}��;<��<����B�RT!=�;�<赺'��O4����X��V1;�*��Xi��C;��O=[h(<}#=e�E=�h��p��|X<����;��	=�'��~�<�C<�����#û^鳺}�\�� ���=�XN=29[���<-?� fh������=��<�"J��\=������y<�u���H<���d��+�M����Z���c�<�,2=a'=��3y�<��;�y�B�'
�*��<G��bܼ&�H�e
�� ���H�s����xR��_z=��w�T�U�����=�BD���=��)��C&��$h��7@=���<]�<�_F=�z�<�	�Bm�/c�<�A5��T-=Pc;=�[��1f�<��R=͙U����<&��E5����F�Ɵ1�X�n= ��;ktO�Y{��x�q= �����<��󻁺��*]<��b=��{��h��&���)������#�4
����<~=�<҈=���C=��"=S�a��@g<P���뗼�n6��}���۶;���(=R8=�C��[�<���������E=U�T�m�'=��<�ٯ<F�Y�owԼ�^���˼`{Y:��<'�=��ݼz�:�� 
����2���V(=Ūؼ{La���<�D'�OYH�P�A�y�<3�]��(0�Ct'=L���5��oJ���9���<]��ӽ6���=<i9<<�2��(q�z�������ڼ�o���\#����=8ɠ;��e=�0�.�;/I�<8d��¾��0�<s�[=CNټ EH��K�9y�^ =�K�;Zxb9�g@��x�;p�v=b��<�����Ő<���<�ˌ��rf�'\���)=��=�?ʼ������<��e; �=Kk=We�����m�:�=I(<!t��6���'�<��ռ�0�+��-E�Y��� �)�6IF�g��ۚ�<g�=*x�;�=�by<�4;̒����E�f�ռ���+p0=)#=K*�=n=|BԼ�z<^Ȅ���:�W[<�8n�qUJ��=�$=����	��=� �*�.=�F�;p;L��B�<`��s�<��=�@�0��B ��N��;�V�9�S2�*&�У�<���<�*�@<	}�����<��=���	�	�+ES��<W- �}^<��5�i���:^=����g��%<���R���i<^�:%�;�>s=�G��ʼD�=4o=ƪX��L�=B�ȼ3j߼vU�<��C=ʚ:���(�!�;5&#=7�;�=�N<�R=a1|���T=.-�={.���;%��<�g��G=!�U�̈������[z<Qv�< �����P<�wz���%=]�3�N��`+?=,�<(B��ʌ�<͡�<Hhɼq��4��e�<�����r:�ܼ���-�l�}Ǳ�n�b�^#s=F S<au�}1K��K=�R=(��#�=
0�;�O"=�'O��$R<�g�P9d=3�P=�-?�A��<;vO:�i��W2;����<��O=�Vd�*3r<I�A=
��4?�����4:�I�=�D#=Z��<筒<��E= )=�k�<�9=)�<b�=�3��L���g�<��=;=ri���<���$V�G�vg�<��X=ݙ<Dtʻ�D�����)=���J'
<`O����;�O��[�<gH'���<0]�<�y�O`=u�f��⌽��p�=y�:�49��u��J�P=�/=��=��u=�m=?��;?޼ �=m�R=��<;Y,�"��<�л�(�<c
�;��
��
�<X<��]�<�=�2=ޖ;~U=1���"�f<�5A�}�m=��)���V=a���M¼��`<�Hk�;!y������ ���9<�?�U�*���[��I=��-<�]�<���<�Qr=ٱG�Gp��N]):�H�<��<z==�3=2�O�F�<m�[�pY�<H <>.Z��)�n�8=�������ٙ�:�~j<�z��u�;�TS�&��=�%��G�<���� <�1���.<�#����R�mJ�;w`��C���׼c~D�F��<T��;S�T<�ټ���쪄�͸�=5��(Ł�%#�U L=�=�c�<�6�����bCükI�=�{r�kiJ�=�H=7����9�<\#k�;�=���SyE<��<��;J^�d@��1w=Z�~��'��[P��u=؇�����<r���˻��N��	+�Lh ��(=�]_<�y��V�=\-�D�Q=s8@s�<�Ag�ס<���;�:�<q�d���C�y�4<_��F�<tov=g2��1=Y��<H�=�+�<Rq?=�5�ڑ��$=�G���J��.=��!�'VF;Bz;�i�� v�<M4,������W��X#=Ղ�M���=>�T����(!�� ���F���i=�ߜ�)�2=gn=��<�q6=��^�(Xĺ?�<iP	=i��ƼEx="�=[Q����$�Ǯ=�gG;�U��0���|J޼s�=����:�Ӽ�%T<d�<��?;��l<
�1����b=�X=���<��;����R=��8� �=�S���?���	*=�M�����<Ψ�<^9�q��<Q�#=[���<�E};<�<��<ί���J�ңi;
�<L@A=�y�;F�W;My=~�_��x=G�мE��<�����G�J�B=��T��rO�(�5�<4���a:��[<�1�<���<�P�<�J=B1�=�<�Y==p	���	=
w�����v~6�֒�<�;�����CB�<Ys\=��x7K=�/=��	=�d2�/Ց<�����*��Z��hż��n�bR�:��޼���[�ż�T=��a��al=Q�"=�źL>��= )E= =F� �"7Q��O�;�m<@`.��=�2+��;�<֨a�G��<�L=A��<��<z0����<	��<��f�!`�9jz���2��|X�A�&=|CܼC ��RP=&�	���V�.`ǻr8�����a҃�cGM�P���ཟ��g�����Tt��>0<Pn���T8=�O���<O݀�bj=u��:��N=f��_?�l�*=���-�� �<�q���~=^�^=��*��d��*7=c�(�F[*=XH=PJ�<*W���N����<�.�<����ܺ���<r�N�?�4�Z�޼K�=2�;�G�;�
n���_���]��M����<i}C=7�%����RC�<B��<*�&��;�����:��J!���;��=pļ�������a6`=�X�<�]=���7�r�t�<��<���<��p=ܱk<b3q=��,�����'3C�A�w=OM������Δ�73��[P�+<N�	�:���B;g��<5B$�q�/���B�YKt;�&���Q�b
�;uJt=���<����-�B���M<@�Y=T6�<�"�;�燼I���!����<K�H������v=0V�:�=8E��?�� ��=�0=�	�X�L��� =�"_< 5��o����G=�5���<�A�<c�!�@�H�� �<U�*U�<Z��;D9��
��Xx=}���,�C�7�<QM����=�l!�Kf����<�F��L����������|��5�Fټr���3aA=]�<�9�<�˻��b=��B�2�I�=��C<J<�=����s�=�#ͼ�� =��	=Pk1=�u��hV`�GO,��	Y���5�WbY�y�C=}Z�<��<�
b=Ӫ���?0�<�ռ|��<]����$=o��<6�g=E�W=��i�*l
�5wD�4�N��=Z��N�;3�W��3�<Q]@=��E=B�@=r
�g�;_��]2��ǀһBt�<��??�<�����x����;�~Q�ߒ�Q��<`-@�_*W�~�������);�S�<�<-aL��D=���;��"�H��<�z=����q�<�bO�&�>�){��U�<v�W=�mA��w�@�L=�I;@��<#@c=�Fż=��;|�g�0C���z��ՍH;l��<'tI�A��<r7��n��<��:���ɀ�=��ڼ��"���<lo�<�{F<�Ѽ�Qw��S=#���R��7�'=��0=V,�<mg);ōH��`�<�N�;��l���"=��b=��~n�MK@<�h�<�r<2nc;`�=�5=��=�AP��S��X>=.��ס����<�v��z�N�I5�������<:$_�n3=��º�޽<�Ӄ<�NK=�;��^�b;~���+���ۈ]=�f��Ƞ�l�6=d��boa=� <���<�N�����`)�u��;A�<��<���;��o���X=Ԣ�<�`���A�<L�i==�@��)��<=�sP���<��<5���t�1=�$�<�*^=d����w�;�E���MB=u�<h	�<�l|;7�i=T��<��@<^��L#b=��;#���~�;@��<g�Ӽ�ⰹ"�L<�I=�j;����;<�H�o����(��=�GS����<��<��;=d&G����<��G=�%��Z@��>=�q�<�f��A�E=�r<�@r=���C��<��E=K��<�?S�q��<3��/�a<�G=�z|��1��X=l�*=m�l�����ֳ<DJڼ�<�[=��<=u�	8ʼTY�<�(,=e����f<\;>=���;����f����7��F���B =�0�J�q<*B��U-�Y8"=�d���(��Mq�<(\ּ)].=X�z�����<���<�W9�N�V�Q��<Y����g<��ڻ�Q�<L�52+=!�9��+�Q(=��q=P��<<�rl�U���n��9M�~�Ǽ�Ϙ���2=�a��l<k�I��Q]�k(�<0��<r�<�4=��<=�\��+4=	l�13%���$�ҰϼՖ�ӢS��;�<���<Z~E=�@.=��+=D��������P��$@`;�h�<����е3�y�\=��R=�D���ü��=��n:Mz�<��Yq����K������A=@`g��`����V=��;�={���Z�G��BXj;[e�<��;�%�b1A�o�t<6�3����ցY=*�E<y����<�VN���<B�<�e��I)=	�8����u\��>�;��R;�@=!�L=I�ռ�SZ���D=�c=��_K�)w�<��������Ǽ|,$�dw:=!���pi�����<��z��N�<w��<2�
� ��;_�<��H�<ir>=|�4�Ʃ=Ҭ�y_;=`P���缃�,=Vt��Ь�/P����<3N�<8"|;���!�; ���JV=g�����Q�z$< ��<B����}��('<���K��K���7L��3L=�[�߉�<K�6�oN=�h�;;�<>y=�>/�����<�&=�o=+<�t������,=�^i<���<f_<�ML=ѷ�<���<h%Ƽ�IE=(�=ߙļ�2=���;�����;����B3*�lo=�3�ٴ<�Ѯ��%���=��L�}e�<�C=���*�
�D=�s�5u���̻���<�|���"u=�H0�O�j<��ļpD�;ڄ��դ��5�*=
�P�"��u��������<���s,i<�6=����k��=6rw<��
=�D'=%a��s�<e��<�`�<<�\=�o>��	=��39.�=�x�<L��;{jE���<���;p�)=�^
��8�H�/;�'1='ü;��d�
=�tS�i8S=�`7�]�@<�#�nH�����;��<Q^��T=�<4Iܻ�Qu<�4����e��f�<��G=#��<�Dw=B�h�V:H�\ܞ;�	�<�v!�.��l�.=�q������1�0&S<�|>�<�;�-=e[�g�>=2����=��`=��;�}2��;:���$��<�o<˕I=�)=e��;y��#�0=�fǼ3�X�V3-=�4��b�<.���'=<��'k�<f�=�7�<���<��O�Ę���wI�� *������C=g�=�a߼%���D���[<��)��<SY=��=2�<s�=��C=h��<wL<RBF�/���V<$6���=֕m��7q���]�l��;�K]=`�'�u�e�hP$��C�<��=�|2;�P��s=��,;��9cϼ���l������G��� "<�z޼��=��r��b!=��<��*=�,6=���<�����ڼ��h����;,$ �&@���P� OA=�n0=�hN���;<:�'���ּ��=�	��ż��Ἔ}
�=�ּ�aJ=�����
��3��=Lk=�=��#=,>ļ��x�r<&�ۼA�U=���=r�;=���N.��� ��`-��g�:-�w=܂H:��μ� ���p=��C= ���G�<��'�R�޹8i�;M�	=k�2;�� =4��=���<||�����/׎��vg=��&<�P8<��c�=ʼ}���� �˾=E���e8�x��<1���O�<H:���Z��ē�� =��H<�s{;�q%=�����+=�6/=�=^E= F���=�r���=m� �� �aJ�<>%Q=}�s����;����0����g��E��nb=�/�<Y4�vE=�eK�"�<�Uh��9^��%����<%u"��[ü��(�@=6֕<�(T�8�%=�(e�ݝE<nAǼ\�l=��M�c��<g	�<�<�<�H=dC<h=:k=��Q=s�;=��<q$Ժ=5��JL�]�*���K���4=W'�<��V=q˻��\<���<:�*���<=hP��;�>=��^�O$E�+�6��i�<z&=��F���'<����dh�'cH���<�y.=�e��7��N�7<�i7�ק�<��;z1T=1�<M�J�k=��Z=|��G���<1O�<�輝�^<�Y�<�0�>]ݼ��7����<�r<,v^=L����F�;@&�<�W�O=�戻EJt�)�v��؂�/g���:�<��6��x�<vko=�jH<ɏ];�мM�=�#ϼ���<��d��ڐ��?޻�������<�1;/f�<��<���<'�<+��7U�;�����e=�~����漻=ew��	y=�=�?z<�+:=��=vO���0X��=w] =�s>=�<���c�]m�<I�<y�<�<=�"���=��<x�w�b��ll=�V��.��W(�<]��<����*$��I�:��3�M�2����<�A=c�m���Ƽ�gQ=������>�Z=����#�;W��hx=�'����{=�G���]=������<���!=�iͼ�4]=&4;r����^=Z�]<�#=p	����<�g�;o�$�	��DT=�n�<���<w��<L��<�(~�S50����KH��!߼c�B��<��r�1B=������=��U��S=�i|=�?�<
� =�/����<�i=Ж"=.F&=�K:���U=r#=�H��㚼�K�;8{p��F����f��==gϻ��<:G\�hj˼��3=����(r=��<�i=1�z���:�
;����Bp=f
��:=0�	=^OG=�B�<��?��=jO��,�����==�Iq��Y?=#�.=����L<�ü��O)=�ϝ<�S9=8�a�	k�'�3=�-���nV<�
|<�s�����g�<�xb<�7G;��W��i�p�r<s�'���=�!V���:1>=��=T��ǽ'���<�QO��M8��e`=/�����	0=��p�e�3=��<3�C=ڀ	��7=瘠<3�a���̼���0�ሧ<}�P�n_;�)ۼ�1>=�)<r�����}=V�2=�6�5B|�����t�;V����!>�&z;%*h<��"=�~�<�hO��L-��҂���<�����<�^H=�~�;q�����f�R|�<V[����<~1�<i��<��B=��<U=9b9�(��!�k=U�;_+=��<���<���:����;M�<|`=¾==��;��Ż�ü uG=+^�oQ��#�Ouļ~Q�<o��<IF3��4U��^A=�N��u=�nO���n;����3t)<�H��T$=:�	�%͉<..f�R�ټd��</��<�ƕ<��9=o:�����Ƚ�<Ť�:l;A=�ר�\"�.E?����<�Y���I%�'(�h�6��<�O9��r��i�<��~�������<�h1=��5���¼'X�;H@�;ߩ�������7�h1]<�eG<$U��"��W;�)N<��T��dN��k6<�b~=![=�J =�-M��.�����F����Qj��C�7�ںxW�<@+�;	�Ǽ��=�%<���=W�<&'��N=�K=Og�;�8T=��<H�����p��{g=���HV��ٻ���x���=���>��#G�W����}F=i��$Sn�����<�; �S�ͺ�<��=�r<��O�Z_m=y#=PO���=�<���<.��=�KG�+ga�l�ؼ�(�74=�� =�ټo[.;>.���<�<1%=$]H�� ׼7<�3=n(4<M�Ѽk�3��*=tՐ�7�"<�(�s��:f��k<�k=Y"Ӽ�������M=�=�#ϼ�:���P#�5N=�������<7���aA�b8n�y�W�gs}<�*=(�;��!�<�m��݉*�y������<�F=���XFV=YB7���0��t=�A��)S�?W=I`z=��Y�=~=X�;���9u����[�ź�Ss=��<LD=�<=syI��=��P=��'=���<Ț�=}]2=1�F���<YC޺Tng�����r�zv��g�F��Oz����`��<l�|<!7�<�.=B���!1=|R+������<ƱJ=E�,���H�~�������3iA=	���/bӻtx=A2t���<
D=�ż3�=|U�f=+-o< H=�������J�=���D�üjAD=�A=�ኼ��&�Vg"���G=�<Y�m�z��<;��,��<��=�w$=tz=L19z9�<�l�<��
�@��=�;ֻ�L0��5���-��/�Y�.<�{=�C�4z��3)=ax@���ۧ��x��黼$�;R�d�E�4=��$���c<���<6����J=��L=~�=�b��I]!��񣽡擼�����U�*r	��E����Y��U����<a��<�De���=��==N�;��"����<F�<�Mz-�p�?��;�L���LƼ�=��d=�w��:�<��&=�E=j���L��R�?��<��~<��L�W ����ť�<F�J�bӼ�AG<R}[<H�?���s=6�&<t"�F�C�<C:<mK;@/�;���<��4�<m�T�U�]�P:<�C�<8h���G=�W�;�Q�<d�=	�#=��t<o�'=�5�;]=r�(�w�(�dЖ<?��@����;��ϼ�GT�Z�O��=��)�#G&=��=�S2�N�����o=�M�,��a=3�ڼ�|<.e�<_<
��|�Q��4Y���X=}v;=o��<�*=�w[|���ؼ�Q�E����=?��<��ϼ���q�<=�;����s<Ú�<�n�� =f=��@��+x��dC=}rK��'�<T =�
X�ۋK�C��<d2�=�w��H�Q<���<�?�;b�˼�u=��=�xc�P�1��d�<�d ����3=�������<ʤo<k$=nY<"�ʼ>�׻wv�o)���Et�Gf�<���<y@�#u:<�Z�;�mT����5u���̺-����I=�89=�z�=6���o����&�+��Z�D����wkJ��y<e�y=�+���$��Vv<=�:=Qe��{�5����8�<�K;;�� =~�\�3*~=��I<�((=%����\�g�A�dj�9�x�9x��s�8=4�=��=c���R�K=�7=��D<�мC��S��q;�G�F��2M�����C}=���<�����=/�.<n���5=*D�=k��<F0g�L	=�_=���;#�=o�_=��<R��B��F�O�;���*N=�rX=����W�<�sﻦ�l���-�/ID���_�?�6��;[�:�=�^r<WY�<���ǫ�;1{�ys�<��U��JP���=���<Z��<W�<x.1<��=�����#=�TS=ļR�|���<����B�n�<]`:��*;�����������<$k����<�g�<E�=��<5@�=徼��ܼ�y0���߼Z�<�o�)H#=�\�;�?��FX<ہ$=�=3��;��N=���s�𼮺:�T�C=ݷ �Y,&�,�:Υ0���򼛱D����:��<�'���0����!�S<�="~ռ�LC=ѫ�<���<W���\�;���V=d�<�$��%d���:��C���=e�ͼ���k=ن_<��Y=9�����<���G	R�:�Y;��K=k1��1=Q�;=�,���Ļܖ!�"�<�38��'/=@
Ƽ:�Z�3<�2����k��;Y��<�ҧ��c2<�����<'Ӽ��"�m4[=���<�T��rM�<J��'�<�>ۼD�s���;;�B��Ȝ��n��1�˻�q=�}��R�V�LR&�����*=傽��5�5�l�]��:#��<#D��Xֈ=<$��0}-�'�<i�=B=�(M<�|O=1�<�9��"��-�<�I:�(�����<t6��8��,�
������J$;7:1���L=}Ի�*��:+��\=���6�^4J���D=�M2��z<��;	�ja���uXA=��<B-R��yB�f_H=�5�|�%��ZR;��|=>>=�=c�x<�>=1>^���t=�3�<+�<Ep+=��S=-�"=�<X$S��P@:��< ��;�O��e1=Ū"�⤄<�����
1�]]Ἇ��3�D=��_���h�Аk�5H�<�9ȼl��<��9�PV<=��L<���݃����=L	��_����=��(�y&2=M���{��0=L'¼��2�k1!=kh��Eռ\[=�+�<T�$=P�%;�mp9�JO=V^,�~g�<��ϻ�߼��<�2K�+��<c�i=k�6�XJ2��3*=)7Һ�������Cw?=ls��ˤ�OY��5~<r�8=�.N=�m����n=�s)����I�n�-�0� ��2;E���K@��
���-�x�	����(=�����P<F�Ѽ�3R<��
=�f�=|�;�����Z��k=��x��J�;	Gܼ[p˼$�<= �#���H=�=G=P�;X���<����5��ku;�=N�伧�I��Ѽ_׼<���ٍ�߁�;M�<��o�t=u9	���(�2�(=ӥ���>�MS�;	&<l_={�J<��=���~�F==I�<�5�4�����:�Z@����9��=+�)=fi-;������������;����<�0�<��<�� �X%�<´z<)L�;R`6<F�:�Ȩ��#���2p�Á[����x���QΩ�#2�W��;o���5�!�l�^��<�'b�8V=S�=�$��ч5=���<oPY�␼�I�<�l[���<����;t��M�<7YT��K����=��ٻ�d=͈!�0i`=�-=}:=��<��ś뺜y��h��<����/��<i�C�&l<�W!0��w�<]'|�x;�g=��U=��=��<��<9�W;��<a"���v< �㼪�=��U�;�=͍�<"�
<{e�t�<fPR�+6
<�sm��2���$W��=?�|�f=	dz�Z\<��ۼ�"+�ܼ=���HTҼ�j;�\F=�Sֺ�2<<�q��=_{=�'[��\�:P	�$ �d0�=%o�<�D������vD=��=��^�����#N	���;��ZZ;�%�:�Iݼ�@=I[<��9=���<��{��k�(��<<�T=K�85"�ud��ͼJѼ�	�=TJO��)r=�4�����!���;�j)��\%���<��<�� ��)w<��<�������i���衛<툩<f�<v�Z=)����6��=�6���]���<uP�w�:=��<��= �J='�-��J=��l���:=�M<<�1��-��<k�M:^*�&vW�r�w�v=+\�	,/�(P�;3��c������1�A�ô><Cڇ<}{�����x�Q<��2<�
���}=�j9��5<;��V�~=
*=xO~=�XA=�g�;A��Z�C��<��Y��=T=�ߍ<~� =M��;�=K�l�flc=��#;�z=ҕn<�4o=L��.��<@�<��;ӌH��RM�'/���*�u��;��G�V?���s��W;�=�ý:�cc=rfK=-r��4=�0X��,=CWC�)�=��=����D.,=^&�$P=�x<?�{����:B�!;NȀ<��j=>>�<w�i�<m����L=��ȼ&��9��<�F*;�z?=�n�<��<r/=��r#ʻo?��=0���mu$=k�=���=h��<��7=�̼����혖�5�`=�H�<�Sϻ��=�@3�8=*�=tI��HW�V_��銼�'`��|o�IEH��r8<�jg=��&�y�`;X1�:��p���ϼb�Լq+�`c,<R*A��	�<ŋԻ>K�<�L,��購��ü�������f= �<b=�]r��5!=�W8��<&�]����x'%��4�hS=�|<N�B���=<��<L�I���g�=��/<� C��6�<d�]��A�f4�<�Fs<r�������W������<�x]=���V��<�[�O��<��"=3`3���l;�j<�)�R�;�R����!��@���~c=.�ӻw���n=�'=�o=�	�,�;~�<bxg�+�=u =�g�"N��p�:�T�;1���@�к�v����u�^�<������
=�+;�AB=��=�<=��=�����=O�<��t<��#��e���<��t��2<��Q;r񹼯��<?*1<�2�}��<�D�<?HA���=�ɛ�<��P��ĺ��@�;d�=��]�Ų<>�@<�����q�<Ə��\�:��̖<3u=P�0�A,��<X��j�}C����;-��w<
Լ�f��<�T=�k=����V=hy==��=*�<��#���P=�%[���=�B=�{��g�Ҽ]8L�	L��j(���8=	�I=� �<��5�`E��豻$�P=��ۼ<��M�&�<T =�r�!A�<+o �o�:i��<v��=��R<�e伱��=jQ���ռ	�Y=�`*=;V �����*0=�@����.=�b{�ѽ�=K���Gj:=w=2�=O�!=a��������n��=:	%�4<�o�;M$��Aa����^g�<$�� [μ��.<�i��=c�<��,=�'�	̺�V��ӕ�ܜ�,�#=Z�p=�
��sY�`-=�j�F�B�</��:�h��"�;Lm.�]5&=g�g=ț(<B ��h�ڻq�W=Z�E��S�<e'�<�.�K�9�vL<iXF=��(=���q��=�xJ�qV9=|�~=*.�����Y� c���X=���<�.�<a���p;~��<T��;���<�6��9;���!H�H��<�����Ǽ�ƻx��<>��O*���ȻF��;���9fQ<C+�}���0=�_�ʼ���;�$<ΓY<��*=:i=�C߼�>�<�M6=��º�=w&q��*��_��<����	T=8�=o%�<	ڱ�1���l� I�<ʯ`�/G��u���g=��y$=T����+(�jX��N銼�~d="�`<e�T�6Sk����[��<�9���t*=g�^9����s=��Y�]��<�Z={���'���<~�4�=�(<��g< �D=
��<�� =x�<o]ļ�>B<Q=��^��;�a=k3n��Y�;%�N=��<ȍf�&�㻟����f�`Wм*��<�9~<��lC�U�A�2=�G=��=9���+={MM��4=�y"=�&b�K<�<ףK=Bni=�?����<ߨW=�K�'�f<!B4�ᨒ�^,�=ū�<hB���a@���<��;#+=A\A��\?:O}=iud="��/�<�(/<+��6�};<ӌ����H�3=�C�<lDJ�RV��D���������;�����4�d�;���	y��K^;�x�:9b8���T=�Ȼ<ӕ)<���k�&�!��;�!<&4�<��S���y<K�=�j*=�r(=�=�Z��0><,�'=��Y�����1�<�=(޿:��>=ꇜ�E3<1�,=,D��"�>�aZ"=�jl�UA���o(=��%=N>a=O�<�60=�C�������<4��;��h�/���*|Q=h'=���;t�R�ɖ��N�=;�<<ը*:v�9�޼-QW=�D=�O5�Ra�?q ��S��܄�xX=}�=z�<�wټ̍���O��>�`��;��1\@���(����;�m�MA��g	���?����<�F̼s�N=Ə�M8Թ('=�`��t�J���8@=x��~<=0<��>�C"�<����kG5=/^~�[.�<z�3���<ֲH;�_��(�<��<t��< ;=��ٻ� [=�w"�"j������Y� 3ʼ^=W(:��{5���=qc0=f��<�I=��2�><������4-�z��<&
F=Y���x2>=�^=�!�<[��;��g��t��I�H=��<������=9Tr�u� <�1��V4=�D�4
�=ը�;n�I�C������6>���u<�M�x

��rk���p�}=���<ߑC=��6=<�t=1����O~�<R=�ӫ�Q��b!=�ͫ���!��7����C=V}F='֊<�i�;�-�oz'=nA��U�?=�7C��:=׊�)S����:�S=)Z=�-<<��Q�;<
�m�:�����z|��z�<.�=�*=��|=�R�������tC=��<�m<�l�>83=�=���a.�{�^�D�<�qR=S��v�<Zt�<�h=N=�=HfF�@�߼��<�~л(3�o��^ٲ<�k=�� =&I�;t�r<1�<6�<ٔ�;�R}=�qL��Լ��`�9�;�T=���<���(~6�Qc=��r��9��c��[��<JS<�V#��,=�2=w��<�1��)C�;J1��)��	U�����`K=�q�;�G�<��=�mI=�p�<cf@=�=�o=+!6<􊮼7X�M�X����<^�"=���:Bx�����9r=��=��	������	y=�uQ��c=��޼��=|���>�<�+<�Ǆ=W%�?��F��;���N��IB]�@F���f=0�i��Y�Il�l�;�����=��&<����"�:��/��1�E��<�
<�wS;�g=C� <��=	_={��;�?9=��;*�<5�/��Γ<5�2=絩;}8=��<�+�kB<� <��d=�]׻�F<�<;߀<�7v<���;a�=#��:'����_<������;,==}b��6�9���&U�'�;&��<�^��M=��J;]ռ��j�������Eؼ�R<ACؼ��2�&Uk=��F�����7@1=K��<�0�<&W��j�<�~x��{�ll��/R<3�'=�c���=<���<[���P=t�v=��C=�^��@7f�����B��<�;A��7�<��_��<�:��0=�J�<�,*�ʳ���r=c^=�H=CQ��`/�;f=c<W��=fT��"�m=��<[=�;=�]?�ɢ-=����<���<�u.=8=�V�<?1M���g;���=������m�=(n =�%�<�x�@�<޶μ��:��=��+;}�=��9=
=D��:�H���3��~X��
a�+ػ��W=Ff<��;=�*9��Q:YǺ�1�k��=��v�����Ƽ�'�i=5�ҼlFc=�ˌ<�����k;��Z;���=������RI<�4G=!�:�/���A<gK���6�<����xK����]��\=,TB��<�Ru<@Ԓ��_�d0K� ��\�b���y�Nկ<���@;� �<��O=��F�a����%�?��mN����<SNu�u�X:�S�gu��qļ�P������t��OB�� �O���(N<���<5�=`ᦼ�=�ʘ#����;Cݪ�Y6<۳;�� ���E�<�F)��y'=�=3�i�����ż�a�C=(n��Z�K=����t�M<� �Pbx=%ٶ�Wi�
�:� �� �#�b�m=����U��8 �;�٨<E���D�=]�=���<X�7��p�x�;.+�<8�=�ļ�<z=�YF�
�.<=CG<&]]=�#[=�̬�0����<4F�h�F<ժ�:��=m�*<�1�<�kɼ?���Jcn=���<7=5��
�;��<�7�<F�G���-<��
=�7S�PEH�{W�<+v ���<z�m�m�<в�<:�.=(/*���=\A/<�L\=�#*�I μ�(�<�e&<�뒽.;=@���=�j���,�����w=�獼Y�A<�'v=}��j�a�E��;j�T=�N�:��P=�ĵ��U���>��V=�]y;&�%$���Xc=��Y��<��<]�,:�}L=�K��$�,��E��܏<&/&��d�<[O��N��2!J<�s	��)="�=�`Z=GM��<���؂�e�< 2=����̮�<�<�;\�"<*?$��.�׌i�&�c��$P=��G������Au���.���q=�/<�3�<4�<�19=���)k=�7���#=]�4=-W����<6����}I��c�<U�h<Bfe����j�
=�됼�R!=
E==���<��~<�2;y&"��o�=(sT<��=p��r�p���e=�lZ�x�6����;�~*�^9x<�g�<��=�y���`�ˀy�i�l<KSy�Y�|�'3<�)����(�/|<�À<7�=p���Ǡ��Y�<��4��h�;�Gd=��T=�C��#A)=A}'��~=�E<�	'�[�<c_=��;��=�{'<&�,���	���F<�=���
�A=i�I:��Լ�&h=�!�Z�c:�=^<#��<��X�<��\��;:Y�8�<ݧ���yQ��[H�Sż��=�1T� ���,��Z*Z�KV�;P.�=W�<R,=�00=zu�R<�<�IT:�=W�9=^(=�T ��:=��*=IFS�e>Y=٬=�Rq<  =��5�����s=���X�]�1�ż��<g��	�V=,�0��/�A��<�C=�٣���<�V�=��z<�c,<`c)=�򼣏�<Wfi��*!�|u3���.�K��<����`0<3��n�=>�Q���=��B���)��<�3��;HG��V�o.��}n=��]��s>=��<��r<_�I=����$�<s�<�-!=�\��C�^��5���{=a�79�#�.׼��/����<�ʀ��:=��_�'�t���T�܀	��
���1���<�t|=��9��*<Ŝ�<3-=�]�����</}ƼH�i;X�=�W�<e=�J�ള�;[��d�k=�'�;��#���5�݇=����@�k�!:U�C�;���~��Rؼ]?�;D>?�1�Q=�o<��Ǽ4��8O��<�5=�
�:#�0��μ�e�k�j���<7�1=Q�Ƽ��߻=�S��Hq�fǝ��_[�0�S�zs|=�q;�@5��fp=|���˄=���FJ�<hX� `)=�9�/�s�R�������N��f)��ǼE���F%&��m��E�����K=����c�	�@�'�x{C�л�<Z��;�R�<e�(�Ǳ=|ܼ��+=��;���abi��5 =�δ�^�D��3=Cث<E!�<m�==��5=�z�?�<x�,�����1<���=Ԣ˼Q�=�W�#�="S=���9�H���R�L�i=@Fݼ�9��t�<��U;�c�<�f�<��2����9�'�w�O�!C?��(��	�dP��%(�<o���Z�����="�m<��L��r�<�5.=\�~=k<@��:��W=�J=	�����U=47�=J.�<��+�UZ�<�������z���=��ߒ= e�<��H7I�x��5�c�L�b�o��Ck=�`q����ԃ?��]A=S�<Ho<��<�'�@<��+=+�D=b��<I��<T	G<X<=���ؼP�;#���7=��d�p�ؼ�H;S< zs;�@p��.=�H=h<2=܃�<S�G�� ���=5=���<D94�������S=e�_�!=[��<B�#�?Q���I�[W*�0I
�4�<��`=(!Q=@�_����uV�<��)�}�\=�:<X��:��μ2�Q=��Y=0��K�T�.���R¼�	c;�"�|�==�=:3��[D���2<N�#�D�;=q�&�J�Z=V��<	0<��c�Os�<�޼�V�<9�L�@.���ʼ8�{=�7d<��;�xa���Q=�n=��!������E����;��%�\0=�|
=v�<;&��S�7<c=��[=1�X�0�<�G{<�۶�Z=�R=��;��k�<�"q=@ټ�rw�|����d�0�<WLD�Hl�<n!_=�4����.���߼l�<�s.�_U�<���<��ɼ1m6��m�=��j
= ���,+=�C���]�r���(=�hD<��m�Jw���5)�L2�<z�.=�׷��2[<[傽�=U�y ��ܝ��ܧ<Q�n��ye=�V��-��=�l��0S�;��o;YMҼD7O�tK��2���"r�t���-�)x+=�Z\��--�`�r=_�-=�0��� �o�=�j�<b�1<y����������R��=�[�<�J;�˰w=BE��3�<7s<^�<"�|<��|��X=�r�<������м�N���Z=z�u< B��F!�<�<�&,==,c=��<���!�=��ּ�7�S$*=?�;ĐH���λ�u�<	�<l��Gz�<��=��W=x�l�jm����b����=�Ԏ�t�0�,v�<4`b��wO��g<��*���;Y3�U��<�ӻW�1<��Ƽ~��\غ<��/�>pZ;Kt=�yE=���<�h|�\��<��9���<F��<{��;C�2=Y�m���	=�tR=cNd� )�<$7�!��$�I�6�T=z?Q�\!��n~";o�j��l=��R=��Z�;K~������ =�8=�8>�9�!мHb#=�f]<����A=�r3�]�޼��:=�rS��<OS= ]Ǽ���g,���K<����ջ��s<��E�x�;�Yu=���<ncy��x�3�==?��:ǓL�[�0���#=e��<��s<�H�x	=���j&4=�b�<��ļ{=] ׼�s�<~�=iB*=��X=O8==��0�KW���=� 3<!�1�:;/���=u��^�r=�r���J�ΘQ=�=��S�>}��L�2z���	�b0Y<��=�G��:�;�RM���%=U��<Pz����ӧ`<D�м��;��N=v���y�^�=���<I=�9�<Z�%=�Nx<�ܼy��[�6=.�=~�Y�:0=W��=Qx�;���	�; 2;&��<��j����;S�< N�<U��1�N�^"c<�.J��L;R�R��=�ͦ�k}ҼR��_#!�|n.��s&���Q����=�Ɋ�r�N=G�)<Q4�?f���"	���!�?=ќ<Z�a=l��v�==r"�<��=F����;�G=�B�;b�<ޤ�-��:6!��ތ<�o9=�W=�_(=B�=dr%:�<��ѻ��b=S���38�b����;\Ѽ�N�e�O=���<�m�L��<$�K��y~�{c��OH0��N:=^�@��<��w�<�P��A�<�G8=���N�	^�^����:Q=�c+=�(<�p�:�S=7�<.D=����3_޼/�]=}�=`��;��3�:rf�/�"=lB=��$=�A<|$4��qk�u��{�+���<@Y1=E�|;e� ����;����6=�M�;�Y���=�03:��μ�L=��;�E"=EX=�,����1X=�~=� �.�꼊4=vEu<�*�<r�6�纾�<�kZ�
���'(�m��^:<� =s<T�~�廳v=`��XQ�}�t��l4=�<!Sd=�B�Va==�#�<=���.�<�T���<������=���;H����)��ܮ�^�=J=z8�h��%���P6=Gi����<9>��iC=��i=C����/T<J*=͏��|��4,;zu&�6�K=n���L�ݼH�<�g���1	���;�^�E���}�{�Ἄ��<�<��V���
<��Y=��<4g�vj��=�"=i*Լ��I=ö<�J�����<<�=-�;A���9e2=��,=Ƃw;�k<�<�r�����<$6���7�Zxs<~U=^73��ࢼqz=���;��#�z����ƥ�/w)���=ui=��L�#;�=b�T�Ac��D{=����ټ�d�Z4�f���g��u�<����[�:N���m�L�=|�8��i�8e=���;��=1�6<bd����e���:�<�C=�m=�B�;���v8=�V<��׼16�t=3�����=>��<��[��$�S��<Nsl�@�o�C���X<�@�B�B���<�Zl=��F=Mvͼ��[�����J<]x�<.p�<�1D=�l�:�'к�1�<wn<ق���O��o=�P[�w�<��M<䗘;!����+;�+;�� %=��7=��`=��:=�k=l_=�ϸ<�	d��Pi�qd"=�?
=T4�:�<F�{<
��<K�\��W=���;�Q#���"��0=�R�0�==}.���1��;q�'�f�9MF�goW��Le���>�q�=��<���;C��=gBo<�J?=ޔԺ��=�E�<��`�PS�<8�?=V)� �T=Igs�N/�<��.����;��5=ґ�;\�@<ڄ5��_��62=�w���o\�@B��C=��(��M��q=i�L�;>s��5�<�\�<�= =$)�<SVv��i���
�9:R���<�k�%�x��Q$��r����<]fR=�\9��}=������<@>�bO��mt=zI˼O)q=�]M=�2/�^3�<����0�2�.={�	�:]I���w��"=}��<�:�_���'���Y�\;Y�6��
�h����:=��U<`,H=��N�
b�Ĥ�;=,�;@�i<��-�Iʋ=,ܵ��mP�D�w<��-=$Jo="�<6��z��ro6���z'G�/�<M�N=-�<BV�<���<��J=��<���<�5=C�<s����_���B0�i%:��J»IH3=łx<��Y���^���<	�V��!�����&=�H�:� �ҩ�����<v�:PU��M �8�u�U��;�����:��s%:9�=���+��%=ϲ6�������Ӽqrȼ�n<w!����;�:4�G+ü`�9����8� �+(��Fkw=Cl*;��H=�C�<d���:�w��5u�;
/	<�Qp;R����T�<p��^�=;�Q<�<�;�'�*�<Af;>�<2F�i��<
��}�H=U<\;]�b=��)�ǵ{=�g�<�Z=0�0}h<�q���=�՗w:��Y=�&2�/��:؝'<��2��di���8�:P2�;i�<$��<���ǈ�2��<`->�H���#ʦ:;'���9="�<L�6�&1�<4��<���;s�5������<=Jj}��c��/� �^�,=��<�����
G<=;�<T6J��A���x<Ѯ|�E=��3�<bZ&=Gh3��Rk�&���@F^���1��|��5T�F�=Lq=����#^=��ۼ��f���!=��$=S���"��=�Ҁ=4�$<�NM�Ѳ��xL/={7����<=>=Im9���=ZZ�<�};>�c9�sѼz�U=<!-���]��ヽ.l5=z������<���<�E�=�Hx=�X��.j��`����<��޼�g&���*=��%�<*�<���<�<�[C=�es=�?C��>��A�<:l�<L�<�Y0=~@�<$�<���&=��ü%V<�^D=��s<�m"=u�X�`�弿��y�������F��DU��Y��<)V7�&S*;�姼QQ!���6�ɲ�<�}n��9=�=��<�u,�l*S<9;a��<�ֳ<B���M�`I=��<����$�h=N��<�v/�@p�<�� ��ME<:�ؼ��߻��=�܄<v�.��۾<��e=vW=��%=�)����P=b�'�=��;l�c=��m<�mI=y��<ߘM<�T㼹�=�NZ�M�+=Ӽ55켄 �u =wͼ�Y�f�=>��<��e��Sݼ���5Yƻ��H��P9=Dtɻ�A�������=DY`=�=C��5]1<���<E�P�I��<���� =����Ԙ�<�~�<Ou=�ym�Q�^=�d�� ��+ָ���s<i|��;�������1=Q��Wh=7{ϼ�ʹ<$��<{���;� =�"��4�F=���<H�< ���5s��]�</.=��=ߢ�K�0;��(�	�!��xY=�\�&�<���F<�ڑ���8���b��k@��gt�2��Yt9��8=���������dJ;<���R�=c��UR�;	̗<�nc=�t1� RZ��+���w=���9(켲��:r���%%\<�);]#��k;�M��p�G=y~b=�o�;Q���6��� �<{*;�Z@=?��<����M��9q)8�O�m=�,=�e]�7�#�N�o<�����9+�	=�w������a=�ْ���ͼ_(ɼ��=�)=s�Żi�=Y�׻�R�@����*�]����]�?X��,=�v_=U�f;C"=`7=�9�<�	y=��;&ϻC�A8E��]b=7?Z�ᅽ�x���a=H&b=������~E���<z�$=)q;<�j�<HSU=�j;�h=�-N��5b� �d��p;�a����Mδ�����-�;�f(=={F�$�?�HPd;T�D=�t	�aG��v:=j;-;&7�i�����;rK����V=$����=jou����~};�r�f�2��%<�2�Ģ��z}_;
dT=^	�<C�q:Z=[M�׫@=����<Σ<~.^�k?�]pK=8�<�U=�ZE=?eN=�;L<=vI==�?�����f�<2r|����<B�^=K�)�u�N���L=O�U<h�g�?���t U��
n��Y�����<;� ��:�M�He�<V޿<h ��2��s;o��wD=��%����;��f=�<M;�X�������d�k�R=n �;�EY=M�8�Z�<X���4Ӽ��\=i���I�p�X_=�,=�9�<�>����6��.J<÷=���3�<gN`=v�&��!�#I9<"�;���30�3 8���<KQj�_�<����4��]�U�kS�<��v�b@`=�ش:�m
�3�,��;�<ХI���ؚ<��<[�<��=�'8=@N��	�;�M="]�	�@�/z<���-�0�=%�;��<��)��1=W�p{ʼ�c��$7=��6�-�==�������<j�7=�$!<g?�u�]�NmJ�c�;�v.��¼�\�"�=���+$����^���Y<�2�<�ā��Q��H�a��<b=E�ƹ�E=�P�/3���y=�:�<k�I<�����b�<?�=��<���R�����3}��T=��+�m޻0�\�NPW=:PZ�?L	��=����"=q\�;z?���V�z�X���+=vY��dcC=�n輔,�<vL�<U��� �a<p�л�:Y=+�ll��+Zl���	<3c8���ۼ�� =�-�s�$����<aZ<��ջ!B <N$��CO��5"�-�=���<��:;]$=,Q�:(��5�A�5=m	;���<�<T���C�W<����L���׼�����*�EQ+�r�U���u<�|2=�C���;C��9�.\�S5I�'�!=�6�<��Zl�� :��q =�}y����<e�9o:I�+-=��;��<��=ft=i�b��Ӆ��k���!h�����c=�`W���=i�=J�;�j��%==8�<=��=Ӛ$���(=�<U�*�̻�=�l��o=��=�@=�k�<�v;yN=�S�?�.zI=�Y�<�D(�e;��K<9P`��d6=YRZ��B�<w]ƻ����r =�<��eZS��$�<PcP�wW���8�<�!���̯�$������ a�K��F�:�_�����;�p�F�Q<�˿;\"=0��M�HNg<歅�'t="��Q=�_E�N�Y�!<��+���<�A����<>0�rjN��#���P=����
�<P����O=��;��K;�Gֻ�&��<=�V7���B��c켩��r�$�||4���H�N?�;�hD<�h<�Y�t i=q�<����Fa=\��P�ݼ�M�=�ӭ�Jx=!�<F�G��Ɖ��Z�0�p=���<�W��=GQQ=A�$;��S=S=0t�g�<�=<�.}ռ[�S><�l޼	2j<�]e�*��0^Ƽ�8<"�\�wμL��u�G=}<U��<�����+��\��8��_��۷A<��5EQ=e�Z=� �'�`���R�%�[��@=�@�<����wwB��� ���<6P%=�nԼ��2�����఼��=L�j��y�;o���ȔC��ys��>@�����fQ�<�e
=nG��H�<&n�<�,��=H�Ƽ<tpq=�����<V{R=`=��y�_k���j;"5�<��B�PQ+=�CT�6#μ�	�gF>=`f�:0�B=~Q=����0 <v�
<)b6=s�z��ͼí�<�@=��=m/=bh��uJ�#T=�ƭ�M�'=F��v��Œ���F��<�0[<�e6�� ��ꟊ�o90�s��<9�=�PY��B��B=�;1�� cq�gT<�~"<�h���:�m<��<z��<wd�6�����=����Y��$f=Ovջ��c�7>�AF"=���;nm8=�V�Ϻ�<�tʻ�識֙��o=2�l��:伛@��h�<>�<ɽѼM�E���;����)����P� �ڼ�C��f'=��
���(��8!=q�_=)���w�Hf�<�.=1@R�n����;�cF����=f=�ƃ���O=��7=��<���<&���t�y�<�_�<�1=a�=�Ce=b ��J������1=Yy� �9<f�<�,#;�#����0;����ݧ�<�ż��=;ZT�������
<?�<=�:<w".����<P����=@\`�{O���p=K$=n[<c�.�] �<q�P=�G�<_%=RNX<�=�dL��=2�{<��/�%t���}3=`�z=�S�;y�g=֡<=�C+=�wc�&�<GZ�<i�R��8M=������<�ն<�ch�Ns3�ܺ8<��4<�I� �=�l+=/P= p��_;�#ڼ���i��<s�;�jI���=5$j;E쬻d��@�
<�+$��Żeh�<��.=�Ṽ��3=N�=��O��#:�!��<|YZ=?*�;�n1=��<��<`ې��=�FN�$�=��黚-ǼF_��_<,��:*e�����4�M��<�G4=���c��<�o�y��<)>%�4H�;��U=T_H�*R]=K�=�h=�$l=Kn��Ϲs�r3�e�u=�Ot�T�G�Ds;H�<L�O<��a�D�%=�k;�_u���j߼��`�=��bx�<�����cs����&��a=>=,W��S��be<�F��<����P��gX=�r��?g=�8�<@@����;���<*����S�<�m�r3�<M��<�C
9�I=�n3�\Zy;V�e={����^'=����K�k=߅���5���=�c�;S���&����[�,=%u�i�t<���Y���&=�7��<��7a=2<{=���;y.���Z=�%@��8���ʼ,d�IO=+��&��<��=
?y���;�������<�<�Iu1��a=��黽�<��S�!�H���k=p.]����<����㾻�3m<A+R=�(Z�?�ڼ�"N=�=�ܼ��E��̛<�
=�j:=.b���dl��3����<-s4=���<*=8񀽍�j<_�@<�����i��2�<Ty�=.?�<Y��IE;=[d[<)����}�<��Ƽ�𐻺�=A:=���)����c�����nJ�-[�z$z��L���o���b��� =p���ܻOM�<襸;�s@�XT��<D�ɼ�b =�h��물~L ����<�� ���u<�:�p���=y�)=A�����'���\1�<Q���*;|�������������;���s�S=�>n���"=zz�������!=�=�<9)=޴M<��޼�8���;'鹼!c�*�3��=��#"<�]=�ML��s]<�-�;W�L=<�<ʤ�<��5=�U9t=/Z}=?T=^xC��K���2<��<�yK=E�T�dh=F��n4�<d�滶N2�بT=���K�l�\�/�?=07 �}Y���<փP=��<�R%=�p}�u2$���
�Y@n�Lt�<2�1�Y�	��C=c4O=��?��-��#���Z��&���L���.=I�U��)���P]��J�0|�=��¼�pt��3x���"�0t���J�<4M1�Đ�<t����9=D�[��mf�ő����-��Uc����;��R�s�̼?�=��<>"F=R�7<�Gмݎ�� ϼ�v����8�k��<�0���i�%��� �Ǽ[?���(�<��-�y�R��`,�X\ϼ�j	���+�D�P��`
�y�:=�Cm=ݕ'=ߤ1��\=X?<߁F��xN�! �<�<�<�p=}-=<�C��6�<7u���>�f���	�Cx�C�@=�`�<��<�}~=�*@�(�輔7`=f�����;�4��j�6�>��r\=t�]=f�C=k�r=�.
;�TR<S��dp�<M�A;p�~�>����=�߷�9���&-=�L<�b=l�=b$R=��e�|�4=��=��'���.��j<֥[=�ȼ��_=>�L���6=I�I=a�(��ҏ;K=�<�X=L�=���<�8*�`�<ừ8-�k,</?;�0=��=�|8="[�s�=�7*���9��l}=W��2�N=�Ku��.�f���D=��=W�!��!NL�o��d�L���<�R���C�m=;�Z=Q�t<`�4�q[<���}�;�q�d����Jǐ<�=�ܼԽ�<:�/�|oM<=�#���̼{�j=��<�򼆰g<h!1����<g:!=\,�({%�8I<��;�|W=W�^��A=�=wi����ɻZGA�?Ϣ���|�6D=�%�<��*��^�zR��*���ʼ]�K�\�H=�2�xvR=�3ͼ${:=S��{���b�<O��<��<W��(V=���<�����<e�*�
Ѳ��t^=|$C�8<�b롼}~�<����=o �<���<VW���R�)ʀ=/�ĺ �lz�<K�F��A=ox<}+b���y���<�����=^|޼�zA�m�8�z�]9ߦ<�R��,��'�f�^�d�F:a�2=�~�<����<���<�< T��á<Zkʻ M休*!���]=�K��[|<=(����w��-���}=�3��O����@��&�<`���
�y�% =��4��=�#3��9=�c�;CE��u�w�-=�Cu<��<�Do=2�p����<�����'�W�:�ޑ�j}�g`�<-+9���G�mz������*%�ׇX=K-���3"=<��=#C	������8�F+!=�e=��"<�|�����z��<{=(E=
�ּf
`��|=��;=ψr=�毼5�[=�vD=�-\=!޼?�1<���=o��fa=�]=�6=G�<��ټ�pj�������<�4J=W��CZ��PL=2���q�;F���-0~��#�4/|<cT���&<;�$��J��t=���O��K��<�b^�EF�����<6��]K=�E�C���g��{���i�ǉ��X\=�6j=վ�;2�,<Z�м*{�<�#ͼ��=�~ֺ�Q}=�U���;=.˼�:<�Z�<�1�Jͼ��d�ek�[���H=��Q=y�<h��<��<-��;�o;�Ҁd=��w�^j��}�(��y���d�ĵ�:�$'�Xf=�E|��@;\ɻ�v���oZ=�l�<�2=���g=�뜼��<o=rG���H�;6�⻗��<�D=�@5��aR=?�-�}6�!��<F�7���8e���E=w/=��"=)��<�=�UT�؅�:@�<"T=�hE����L�;� C=M��<��߼{rżqs�=4�<�&�W=oZ�<c<��N�;��<�;�;�L��ݧ=;kY=��V=�ֺ(-���\=��=��<�����%�$=���<#��nF�<�d���="|�N���M�<�[7� =f�=r��k ?�i�V=e�8<�E��d⻠����<�%=�R�;�o�����n;=�=�9�l�W��ϗ<~�;5�<M��Z�<�=# ��}���ؼ��2<Y#���5Y����<'"�:(�E���4�<��<�#��"=_\c�Q�8��W=r����==�%<x����m	��Y#=!c�<!U,���D=ݒq��x=2S�<Ma�y��� �.��
J����
������K��e��W�<ǂ���+�<X�O=�����k3=�����"����< F��
=�c>={Қ�T�`�����W��ŉ��I�=Y"3=�X�~�~�%dL9�ݎ��c��~� �8�W��<
إ�|(��0ʻ\<Z<���<�^<�]�<i޼%Lc=3��<ue=�j�� �;<wm==|���'��<)"w��=I��<=)�<}�);��n��������v�ֻb>�;�-#=���&\����=�뼻�$�}?<�U=���<��T<�j%=���Q!=a�=�0&=Gk��ۚ�<�Y�Ҹ�<�Ѽ[z���C�_�ϼ�=vO<=���ZA8���<�ϼ!=�֤=��=�S=k{9;���5Ip��RG=��<��<��=�E4<WAN<N�i��򼨱T��1=�܉�]L=l�=U�i�
�	�Z�t;����0���:4�=��~����U�M��d=������)�U:B=��ѻ�,=uU�<J�<�=�	�qZx�A���f�8��<\l�<ӫP���R=NH�Ȑ1=�K1�A�<����N,=���<�~�;孼��-<�{D=PH�d�1=�J��#C�2L]�-��,���	t�<�<�!�=��hod�/R�<�k�<�i:��AL=ce��h;�X)��)��;��<��K�4��<V��<�?C<�}����r�B=�ڼ�t�<<值w\ۻ��F=R�<L��u<=�=��m=��<��;Q=�C���b<hո�7�����;ї�:�@R����WK�$<�c6V�#p!��D=m�S�8WC����n/=�CC<A�}=M��=���[7=i�g=/�<`b�<f�Z�H�z<����N<�:Ҽ.�;_B�;����M=��B=ӕ%�6&(����G�,=����Jr=*��<U�<bPv������=�'��^Z�l[m���]='ݼ�1?<#1S<�����D3O������r�;�c9{N˺O-d�`s�;jV�<A�^�{�=�י<�D�Y������C���;�k5=�a#�3��Wb;�c��F8;���2:�#Z����;��;�[�����<�_��;�k<�c�<o!�5���T��<���id(���,��Ѽ��<��/<�L�<p�-����<I̊<T�$=
0f���ʻʄ���#��{Q;X��=�;�<L�<A~~�۷!=���w�E�ϼ��<H(B=5Ň<`b<�û^�=x2?�E�<�p�<w<��M*���=�e����^=n�B=��<=R��^�<�.9|�]3�����5��ݷ�q)<=�������)=��ͼ�:１t�<`z�B�0���=�}ռ��&=�v�;S��"�&��7D=pĦ�����r$c��ڙ<�\t�9�*��$^=��4=0�<���̐I<i8��͈M=8�U�|5�wD= �c<�>=F��<����/<�6g<�@��<#=��5��}9��z<؀<Q���]�}Ϸ<BW�<+�+��4=�L<6`�;�<��[�<zl!=�ȃ=��鼸/o<dS4;�/��� =��)<ͺ=}H�<4C�<�$<��<�>|</;��QL;Nd��8�)=v���EG<�J�=�GR�ӊ��΋4=��W=������7����6�J=9 �<�R�<����0=�H< �,�Q̤<��Ƽ��,<��ȼo�1=O�Ǽ���<.Ƽ6i�;J�<��$�����37J�1��;CI<�}`s�м<1b�O��<r���D���W<�9<��>;i��<IP��Aj�|�=��r<�H-������1�EA9=�=�J,�����Mj�3�༘�`;�w4�OcF��,�=�r������4E��K�<�;=��<tC|=mu����xyռ��6��GL���x<,�>��v$<��<y75= �V��G+=�q�<��n=�Q�k_�9oZ�2k�<�@�<��~<x�:B�O�KI=����ȸ�<\hS<o=���7 =؆��[=�pj����<���(FӼ�� �XT�<���z�c�1���=��=��<��Z��ݼ��/=��(=��F=�l�<pj�<��#<���3� <�t����<<��y��x=^���d�$0�<F�L=Nӈ�6�i��M=v&��Ҭ���A=��
�Oe���YV=���<������=��
�M?Z��\=:��iV�;�8�� 4=��q<L;R%z�����<����"�K���"�w��A���Y����<yy=SI�<\��=XK=˓�<T���ع�:�=��0<*_d=�+=pn�: �a�X:8=Z�[�E�����*=�)-���i�ǼU�)�u9J=�x�GP�<'nr=N]N;_�I</��< fj�z����<?7�<0H�<����"ջ��+����;ld.=|s�j�j�٧����#���<�IӼ�{K=�����$�g�E����<7Z=w�x����<��D�[�N�h}�<�Qm=/%=:TQ=5��<3�;�g[=�RV�piY=����Bw==�n�s���#k��gּS��;ך<T�<B�K�F�2=�X@=�7B=A�
o�<��T=�C]<�ۼ��*<$�J<�=�4�˳��6z=�z=��=ѡg�s���/<��6;Eg=�=��[W=d/=P7��ы�b��:ϔ�8]�=��x<w�;=\l=��<��o�QD�+��H� �<��4�	=��ʼ��X=�	"<�1p=���Ь��b5�i�����]�f �=-g��5=��<���<��h��;�㖻,E-<��<�:p=��z�����<i=���dɰ���U���#=�pl�p�S=�&�;�.��5�<��;rP��û(�G��K2<�<Ήn<��K;d��<�r<��=s�;j� �k��l������m�:�'�<��A<��}�[��B����$5=�޼/�<@T#�A;�����7�<��C=d�a���m���>�C���m<�r��;l��=˝�<�WV�ñM��v��c��Ǽh�=���-�b�
�=�3@=?%]��94<��%� gO��g�;'�1��0=�����h)�
n��1U�;�PM=s���,���y�<�,=7�η�;��<�\M=�Y�<c�<�^=�	=�=��<�8=}�#�z�(3>�vh�62+�޵��i�T��A�=	����[����<�U�{��V��=�3!=�)N����=���Y���@��[<n:�:1�5��y+=��J<&��<l?:=�8H�nn�:�����ѝ<�3�<ʶ6��N^���#;|nW=��~�E���U�R�V�/��ʹ<����;R��;���<;����8�O�<�J�<I���Zf=�Q�^�Ϊ�<��C=x�e�?�Eaٻ�&=�N��H�G����wRN��u{�R��<�gX�.X3=�5�<1�<�=%<6�l������y:/=��<���닍<���<�B=
O�<ls�j>�<T��O#=��%��B�<�+'=�ͻ<A�D��,�U�Ӽ�i%<���;��I��-�м�G=/���W�In���=ɍ =�K�25j�E˥<�<��v�#�;����<�J����n�c�[�d�U=��qS�̌0=�'>=���;@��,��I�<=,�%=i= �<(�
=<�*���%�?��|����ż3={����%=���<u{���3�;l��<
�=����B�<��=�^��<�<?�3�!=�	׼�~
=��[<ae�<"���	��X�=�d鼌1=`(�<�� �qG�<~�N���n=�d=L=�x�D ����!�b�`:S��F#���=���Ϥ�����XT��K�<��"�2��<m:�B;��޾�A��<�K�<��|��v=�=��3=+~�;W�=�鷻��'�U��.{(����<io>���=8(Y�5=��6=���g7���ȼ"�#�C◻$/������m/����|,�:�QY�@1D��<yǻ�U=P�ļ���;:z���╺d��+���(�<���<�I�<b�c�14P=|Z,=���P(�)a<,{׼��ټդ�"<B=$=�rL=eS)�@�1�,�n=�@�<"�伃_�<+�<h&#=��A=ĩ��;Tt!���=瘦<��:�
�l�[<�nټRC=uY=?�	=�i��=�u�;�~m<nx=f���cA=�=1�U=�?P�2aB���`�p���t�7=N�)�Z��ʼi^��C	���=1bJ=K�M��=��N��	�<�\=�Fp����<�ͽ��Ub��*g�.���2�ȼ^����\�Z�9=l�M=i˼���X�<ך�<�><�xZ��?=O?m��qR��a�<`}<�By��G�;��:�g�8�u�:K=@��=p@�<�����/<y��FD=���;��Z=?J���̼2�,=n>3=�	?�Ӡ�<b�[</����<���</�;an�;S�r<�>�f+��ON��ϼ�c1�=���k��<�ۄ<޶I���B���-=���;�
:۟мFC���/��7<�*=�e���<<�l���(:��<��
�F��;d|~<��)��<(���S���<Q���)@���$*��#�<X�帟T�<�c����*�a���=n7�<}�=eûձ�</�<�+�<�&�.�B�g=���jIF�g�s��1<�^��Y=<��ݼ��);ʖ��4;͘�<@|�:Џ%=aV�<~��<�c*��ӂ;,���*=;���k�:��`<�Gɼ6;=��P=�K���P�U���+�.�����м#9��V=���<8S<=��_H<�B=Ӻ=����ki=���V�<u)=�V};�N��HM$=�� �b֒�������B�Ƽ�M=�j=�$_=M\)��V=,C=�3���7�m��"�1�;�=�=z��W�"=c@�^�!�$�;�h1��A�U��<NBP���ͼ�[�<�Ґ�R)H��^��'	=�F������&a<:�����P;��λ*o?�켋�.=�ci��6=�� ��i�<K=];�.o><Ӳ��5Za=�Y��wE�TK�<\l=-�= �B=�P=��;j�Q={լ<![/����;\��;
3�Qw�<��=U�<c��>�<!.5=��=m6�<`�<T'��r�<*=��l�� =;�+=s����<�UQ=�v�:ID�< M=��=(���L�H9=�,=�T��2�?�<k�e��^>�v�^<~S\=�%�<4�ּ�s�<Q���HB�<b�;g#D<r��:� �RDD��˖<�,>=���;\��lb=l��<f:<^W,<料<~fļ���<�����>��<Q���7V=�H=��1=�P�<����T��ss�<�.�<m��;=�;��[9=9�<�.c��6-=ܫڻ��)�n�x[4<Sm�;�16=v�G=C=��3=>И<8m�_�)=0���KP��@|[�~�M=����x_�����������<giw�d<��ż�����Y���|=3]m�*p�<��p�UO�2���5
���g=��c���:���z���^�1�4�B]���E=���<*%�<l�_�hb�<��y=��B=RuA=�8�l�`=��(=� G;�48W*�~#=�r;���<�0i=p�M����3=v*F���E��*h��Ӆ�R+(�k���^�;r�<�f��I>�;ވj�>�(��<��ψ<Q��=�'&�(�8�M$���3=g2E�$�<7B@�;�y6�.���}�̺�ü%?*���.�0�i�D^^;��@�9�D=z޻;�f�<y6<��i��I=lA�:>�<t�,�@-�D�Z���H=��*�����Ɓ<@a==��&�B����5�KP�<ou�8!����<i�A�o/��}z�x7�<�^+�B6k���+={�<1��<>ĺ<�Mӻ�Y:=�TP�%"t��⼖2��A=)�1<_1=@h'�8D=H =�l	=13�<<<Y���Ǽ�;#=��C�|��r�� s*�}�f�*RE<_o�
���1��<%����𼖗��ȴ���#!�5AW<N#d�`�"���;U=)2��F��r�=�g���<j ���켢�$=u��<J`���e����=�����vO<9�]���`<s,6�/=�<��1��-=sF$��2�<��:=z�<�s8��F =$&=�K<^� ��I�<���<[�*�f���O���/��J���G�=��Ǽ���<-_=�0%<
O�- Ļ��<�W��m�;�$=��u;Y�Y<�+=<d �I�G�{;U���h���<{���z3=��m=[4���;N?�<4�=ml=E�p�jV�ϣu�eQ=��<P��<&t-=��)�x�1=YZ=�\��c�<^�]�3�����KkN��vx=�D켬%=<#�=9Q<=�+ļ�T�<��.��MX=y_�Q��;k�5=+%|=g��=��6=iLU�"[F�fM��c'=���<,���6�������#<���A4 ����)�#������b�=��>~��̼�� �m�=��<\Qi��=7=�a����<�m+=���<�=*����/=��<�rD��%=��<Ea��j���ϼ��z;�����¼�n�9T�WZ=�Y=�^V=�d�;t��d�+��s���w	�yZ���GƼ��n;;��=8�|<���<�%=��V�z H=l)�����<�,�<nl�<g�,��q���Q��R�<�(='��;,��n�ۺ���Fj
����"�B�.��;q�;���<�(j��# �aks=���Z��<>�=����Vs=���<��-�¶	<�$ɻ?�L=��<k4�ǭ�<~`5=K�~�gi7=�=�y�;<h=I��]t�.�+�7�I�XH=Z���m�;C*��G����B�#���\=R�9=Н<7G�z�A=3X����ߤ<}f=u��<�u\���=¹)=�=�I�pTi��̆�� =���<�Hr;4=����l<P��mԼ}��=�q"�r���:���=A0<gє�j�/�k�*������i�<���<�wQ���<ˈ�<���<6k�B̺�꺍�<��&�uL=�d><��+�"�T=�|E�:�Z�z
e<>S�<|i#����AВ<'��;��<L2��64=�H�<e��;�]��t�F=9�׻��c=��?�I�*�~����!�J=�j��ߋ:c�M<������<G<�E����;]�<&�_=��<��^�*�Bd̼-Q=�j��BO�o苼���<��=�!E<@�̼��m�+��<��d<ɬ����4=Rc�<8)�ۈ'=5{%=�9��\U�D��=�J��]?���=��;�Б�YW�<Y���#���w�<�E��}��`� =�8e<^�5<#�<r�Ҽp���%����9<a=�<rʙ<M����<3��=_D=�#="�=���0��<|2���=���/<=\m��-= �ڼ�E�t�<��K=n$Q=���<��r��;9�:=�H/�E���?���(N><z��<U��2����R��k��3=�l�<gF�c�g���<*M>=�}�<��)=Z�4=�O=�`v<u�=
�<�>=�L9�"��r@=�4̼�����<=>/8��I�����<�I-��ff��r� �d=�w�<I�a�,CM=æ0�������<c;<���[6=���<��<YP��J�c<3c=�X����D��0<d��<M�z$�<�0=�߻j��6܎��6Z�ƛ�:{8g=�qK=Su=�Y�G;�TҼ�B�2'+=|�4=�
������R=�Z�<Q�=w�4=�Z=�;�
<!����=Dq���ğ���!�h�F=&�C
��sѼ��1�g�a����<��;"�a=�M=�W�_�<M���=Z�Ӽ5s�<��n=�a4��گ�|n=�&6=��<T�=}�m=�y�T�$���"=p�,<��{=6ym=)^�<ػ=ӓQ��ۊ<�VC=,<������<��F=��J�<�$=6߭�XG�8_�=���9�<W� ����;�����O���<u�H�tyU�0&T�͋��P4=s]6=pE=+�	<��0��5/���S�Du,��>���;J<<S0��JQ=E�m<F)0���<,wü�o�=�J�A�K�>Ŀ<�%�>]ͻ��<��;���<�#�<h�%�<4ν<��5�/A�<�D�;/�$=Ęm�\�g���O���;�N\����N<��@�������<�Ύ=}�����<X2����1�<�@��
�<�c�<��_<�`#�ō7=��e=t =*�7=�h�<�Tm����<��+=D�P=��[�#�x=�{��ج;�X�OB=T��Y<=W�8���^<�̻	�=Uk:��2���2���	=�BR�L{�<ͳ`�u�C=�_R=A�I�����3:=��B<���]�-�;=�N�<�ƚ��gr=����l����!�����!��Ǽ<�H=��ͻ_٠;��9=r=l��<��<�a=�����?=�u>=������=Hzּ��
�S=<�&�P�P�ZE�rQ�8��[��s�Ч�;]=�E���,�<��"=y�J=��<N�E=���ȝ����;"F}�ڼ���X=���<P�<��
�n��:��+���_�)'��sF=���l=���E��x6=��R=%j��ݚ:��=ҫ=����D8=��Z�L�'=��3�mߤ<�d�:�-ѻ���"���0S�1�~�^<<�]��xx �kY��RI<+78���.=�T]=��=��5�t1�<�f=D�����<|��pA=�^�;�8�<'}�<uY:��-=9�F=ޝ$�,]�����O�<����=�g=��Ӽ��E<U� <��ݼ��R<�<�����x=8Sw�"aF�"�-��Pc�OrG;q�g�d�k=�8=��ϻ��ǼrO�4N�=
v3��z�>�|=
a^=@~e�h�n<;i��q:{=�U<�E��a{1<��F����<��i=��<¹;=HYo<�
^=93�*b<D�d=��<�?���=��H���G=, �<+��<F��<�_6�E�,�n��}I��nk���*<����,��%�=CD=�������<r=<)��T=)7�c��<J/C�5f��J�< ��<;L��`I^�
2n=��Ҕ�<�[�;�&�;�>W=��<���<fE=�N+=��G=6���œq:_�¼)T���%=b07=&�=�-&�w��� �%=}�d���$<���Տ�<��]<ǣ3�4u;=�۬���O<$u+�<v=0��<İ�<��&=�϶�Y�^=k�<���K;=9�&<t���-�l�:W�G=`��W-�<�,��QBмnR=;��u���t�:D�Y<��x=��Ƽ0-P���6���ȼ1��<�2��[oE=�;=�;85�b����(=��3�j6�{�;P�������p����< B�D�5=��;�ڼ%J��诼D��<��A�� $������a�Mӕ�9��n�<ξ=}�;ZA�<C� =0Қ<*i=P�/=����YG�=i"_={|���e�FgR=GX������<#1<b�9�c�r<����.����6�,='���R�SG�:q�ʼ�$=hT=�ZQ��"�ћ��gT
�F�3=_�<��=�;�����=���zQ��ّ<Ⓔ�?!�t9_<�W޼�+<Da==iwy;�8;6+�<�K�<GO��w(=�E;Ju��m���	��KQ�د�<��B�h���£��R����<�]��M�<�J��'<g�<�m=a��s<�2<^�ټ�4�����9��͇#����<�k+��:;����7�<��.��f(=�q�v�6=/;R=Wy<�0"=��g�=���gd����<"�e=�����<� ��2]ջнX=-�4=��<�o&��p����J��46=�*A�7�:=�{@�$ſ<@A<Au-=Bm=�0t��O�<��o��=q�'="�<p�I=�%��
�<�r�������p<��;�8��LN<��a��()=L�:�?=V�X=�<�iƻkE�m�=�K���(������#�n��k�<�2<�:ʼ�e%=WP=��o�f%x<�}��]n�� =بڻ�Q=� B��9=�H�<}�'=D�;�S=؝�.=�೼|(=�4�(=�Q)��*����Z�%�<�)ʼ��a�P�X��=���E�!�Ŋ<�,T=���;^�ɼCP�`#�;����ڼN�Y��7= �l���i<���<idp�sQ6=�5��w�e<aH�=u�o;S�t�װ����7=J�\=v���]=2�	�g��@ 9�²�<��,�����值d`���V�<[�J=��=��:=�f�=��<A�T�����<)Ⱦ��<:ލ<�G�<{�<�
�<��2=p�M��Ψ�>{=�D=��=&+�=����1��g#<�V��ydP;�A=��*����n�μNB=gp={t��G���B�<��R=_E�O/��f��?Y=��<g���ù=����P��<��Ǽ�Y:�=g<��ܼ�<"�k�Ap���K=Խ��1�:�z����<��������Kll=BG�<{�;�Y=�g������3=_V��	*=��=ġ<���<��= `�<�g�<$B�;�6=!�<�$=��t=M.�(���ź%�9C<�ݎ�.='<��j��1[�.&=]�=�s:���P����<�����^ɻ�L=���<0�K�_<B�=)ͻ��[������<�^.=��9�FfI�ΞZ=-��<::�<�Q�Q�O�����m�ػ>���&pǼ�@<8��<��<���i�.���;��^a6=aK?�,���7����B�p"0=���;�&����+��q9�%-�m9=�=��<�g��0.��=�t"��L$=xj�<��ѻYU=s���!�Q���0��7";z�I=�
�-:J���<�n'=�����&=���R�C��'�+�[=xG�ߖ=������X�1$1�聼{���ZH���X�)��9�j_=��'���S=���?�%=��F���<O�J��J��ɉ=�=UoK�yp<�I�=>l�&�u=	WP<��l<��=x=��r���@=	ˉ� �r��<k��cj=�ü��<�)?=��мl�=#h=�������<��W�����L�sǪ;��<n>�7<  u�ES�=��A���1�7[�<�RZ=�*A=��\��<q>=�u��1��� =%�:=<R$�)h��>ż���<�K=��3��گ��-p�̮��ڡ<1�P�/�<��<l{7�ΌP�=t6��Kt�|f�<����|���=�8X��k"=�B= 2�<�Z{<;���²<�7p=z��;�A��e�<=�z1�t�l=Ob��9
��=?=<F/|�����h.�S"?=�d���4�<^�m=��8=Gf*��ﻹ����?y$=��@=Y���L*�u�<8/ȼ�D�񦊽�aܼ�s��m=�F,��|<�J=�ߛ<g�E=�9��@8=�	=�F�;T@�=4&=�b����c:�W<�	��=�L=��
�	�,= �C�:W>��T���dl=d#�<>懼�j6=()=$"	�@� ;�=i�݀l�J�C���b<*�	={i�(Hϼ�1�^��;T�t<
���:���;!���o��<��_��k>��Di=�N=E���j�_�}h<�?=�/=�J����:7=�J�<�7�=؎=�ɧ$=�LF�l�<ۮN=��A5=�?�<�V���= O0����r�=��=Q�<X$����;��8��oD�₽����z���A��;Ej�<�Q���>�j;=��.��<Ha=��("�r���6<7�[=��� �;�6t��:�SW�� �<����)=គ:��<��=\�!�LF#<���;�/�?L�D����T=^->=ђR�KÙ�/׮<$�<)��<Z�T�=]����N��R:0=�6�<�N�%�g�M�m��ּG��lX�;T�(=�z����Q�5=�*f=���<�A;5E=mIR=�:�l�=l)=��(=+�<M�]=c�<��='�C�V��Q=0��3.�� �wY��ܥ`�� ?��at�<{�;J-���K�<i]g�U�;�|��;An�C6��<=4G��x�;=xw=Q<�i��uͨ�\>��==1;�
���eۼT��q;�F8=+'X��I2=����B���l�ݼ�2ռa�<��;؛<��4���.��%&<qk���Ӽsr�=��F;T��R�H�0<�.��}�b<O�E<n{�<�>�^/�=��?<&SW�4#8��W�K�����<�%W���k=!t-=k;=�2:T��˳:�!�B��خ�<�Ij�a�%�c%�S4<=���=">0�k�=�k�<|�Y�X]F<�uq�rڻ�D=J@��o,�<�� �X�j��r;��HB��cD���`��
=DP�D��������A9!�Z<�z=�W=�$�8�"=��/�Г��o�<�=�ܼ:��lz���E<i#;�#<HѼ�<=y=,�<0�L; (��$�o=�;O=�!��N�X=;	�̅�0�H��b@�RoV=Ý$=�[=G�=�j�<(�w�p��;�$��K<	8^�+;���;�;��N=}x¼��;���N����<�9<^��<�d=�\=�~g<�z;���:�`< =7��=�[ļUׁ�=
{b=q"<�}=ٳ�=D��F�O=��=��?�
 =0pD�χ�;,P<Ԅ���;hy= �k=�6������p=�<쐱�}Z=�ˎ�0u0��$�&R_=��%�&tP=`�},<ܣ`��{;���8�j �<ml<#��;��9=����Xs�[�=��I�T�,=�Ŭ���ļGی�L�*���<��b�*i���p�<E�D=|$z�c�f=��f<�债G�廞�l� ���!���R<�n�:�u=��ʸk]���,-��Iz�n�=
�����</=Q�B�B�1�����@cD;�==ۻ�O�0�vL-�2�j��z=@�;�L�U<��<�Tf�X�a�A��<u˛<�CT��V+;�%=�+�Td�;&���S�!��&F=_	����׎ڻ��=�E���֠<�j<�h���!�mU=����DK=��#��4�;�M�:!ɏ�,%�<=ݹ<���;g=��=�i �Z���'~`:�q!=�_�<�<�;�S_=�W�<�*�<Ӄ�:H�g<��,<v ��*=��<*;]=7�O,=I�/��5=�'=`x�M1��q���R=���y)<�1�=��W<�	K=`+=;$D=<�纟�u�b�W�F2󼰁
:=�D��D=rBH=4d���^=����H��<�Dx=�<=�(�S|=
c�<���I�)=�׷;��=B8=�!���!=1	<�o�<ܹ�<�x��i��(�2=1�
���;;��!�D�#./=�L?��}�<p��<�T6=�n#=WO=�eu�IRl�j1=��X��C� =餫<��S=m�=Y�s=���;��&<@7<<�>G������=�n;�>��:��b<}��@�Z;NF=��|<ȕ	;h�'����<v�=�2�<�b���[��&�<��ysh��T�$�O��#<�$=�7�;ꎈ�>�=i��;���<���;��:�<"[F<������F�:(=�o==�)�<64�#<��U<"1Y��'�;iK�9��;��9��=��r<���;�>|=1�h�M-!<s5����c���e��3=��9=��:Y=�?=�3�:h��D={,��
T=O�w�ޞ��x8==�?��x�<>�&�UQ<���1��`<��dب<�.��u鼶�'�M�;��\=-�>=�,<4|��3��k�<�R�
RO="�/�'����<0�ڻa�5� s[<|,��7Z�ȥT���C���"�W=�:I��<�rE�L =k�7�gZ�<�d<��Y��u=�%�k~�;y5*���c�B�I<`� ���S����<$�M�0�%=^3���1)=��%=0��<�6_=H�!=�!���[����<�tJ�mYx���Г9;�::���<�z�:w��#)�����$/���-=��l�p�6���x<�:����`=2�-�l任!��.��oD�m���E�X�=�($<)���&��$�<ˮ�����<�A�=�=}!K=����h?��2=��;e-7�@�<�Z�2B=9Rf=���:y�D� =	��<[r�<|�X�C��i];�ٍ@���<꼗g＄ɟ��Hj<�,1��>=�X���e ;=tǽ�C�Ƽ��*���:ׂ<4�����=�Վ;��Ӽ�^�<�}:=��R=�-�<.�6��E˻�%=M��<d�F=�=Q�c�q<����ֿ��G��<�đ�$�4<��:��e�h�<|�T=Q�޼?��<4/@=$�����ڼ��; 9�}5����<߮|���=	�F=BǼ��<RqV�_=j�V����;=�+� ����%�+�ռ�C��==0ʿ:1AļR�j=ތ<�C�<{We��q1���G�H�;V�=x�<0~��S���ջ���E@�<�wn�?Nq����<FM'=1*��TļQ�S��)=�q�;IE���v�	,<�*��R�M=��ۼ3�=_c�<��%���J^�<7�3=wZ�<!^�QO���K=���b����<ۙ����:��!�ibB=�mA=�$/=:��/:c=}��<�f<_���k-=Y5��Zn<H���>$��|�T�S�����y'<��\;�~���ļ���`E�C�|��n��7�<&t��^����<4��<���f��<�L1=$y�<-s�<kaT=�j�DI=��=Rݰ�A�ּ{������;�s;=G�[4�{�|�=��
Q=aEu<܅�Ĥ9�t�=���kn:�Q��<V��;"���^��㼥Jü�==j��Fkn�D�7=iP=�<;�a��W�7=Kc'���<e�X���=]�n�L�A��/�<�o� ���$=']�=�L�<՞�;��'=�'/;}$=Etg=e}���q; �B���<��y<���<6��^_\���<�x�f=^���ż#M��o?=%1�=[�m�~��;;��;�T(����<�췼�Qw=��ռ��a�kG��3�w&=�q�<^�#V��@�<�2���/��$�<҅=g9l=��!=��V�����߆=c��ܡK�F"=�|N=rl?=R��<��r=r�< ��j�<L�:<9^��c����[��&�`�GOr��"(���=UV�<3��T<��t�ɻǲ,=R1=�]=W�<~�=�8,=��z��@�<P��<tx+=|=��D=r{"�����<i_�<�KK=�=i���Y�2=�!=(iA=(�t��&8��z=g9d=��1= �<�&�Z!�=��d�<��a=R0��vt�<	�r=��I������껜M˼�A<D`��z��<!8 =J�|��j<=�y�I�L�(�Gӥ�ۭ~=�c=b=�lǼ�6=�X�E��<k/�G<Q[���=
~<l=����!=�==��'=��ݼ�0���=ְ���q�;��w�4% =k<I�J=�h,�lڻ�*�<w&=_����F�<ø�T=���硼�KN��tL��2�*�K�����$=KW�<�<[��=�f��K�S��|�3޼'�d<��ټ�-p����I���e<a�T�7)W���;����3=��G��},�j���к��a=%�=	+D�O���=u;=Ld�����;Z��;z"<|э�5{=�<Ѿb�T���V�<��G�?B)=�2�;�4�<Jm
=:���e�}!V<��<?�=�/.P�]�l��-&��6��J=�d�~+�<��h���B<ƭ<Ax�-�׻��a���=�2@=@� �<=c�<�*e=��;�?;N�=�Z�;��6=X�)�!kC�T��ø<�== W4=qh:�>c�<�r>�ǭK��D<V�B��d�<��ѻ����i���0=����)=�k�;a�=s7p<�j��u�\��ts;���bk=�j׼O����/.<�V_��$��j�C��$=v�I=�L���=tپ<�Z�:I>���켧��< � ='
=zU=9�=�>+�[ˏ<N�<��*=kU=O|�;���~��YO=�P=���;��ļ�(��<n����@��_�<�$h����;�)=��P���� }<�k&�*Jf<���t�P=��&=�nX��������U���]�Ԩ<�w�5�K=a�c=�n�'7���o=J�<��<Y�=�m=.�<���<ɠ�<K��#��<��ּ�2����}��=U�AW�oY����<��p<��:���-=�#?���=u��<Q�y�d��<y������w�c�L�0E����.=��J��t����:5�S�s>� ��`����--=v�o=�:=GeU�\F���ۼ�X�� �3��.���V�̈= 3=a]�<&h�<��:�.�w�Ի�w�^�ϼ��2=��4=��d`����<��==@H���z =�!��b���(!=C�f�w�<����<�c]���=U]=�=@ڼ��r=Ò��Nd�ڪ6�G��#�=C�f<kY�<�?]�u�����<��!="*x�=M.=f;9<2G<+�|=/��U�<�7�A����[�g�X=�������Ђ�<`QK��%=�G�/=�=��<S�<w�=|���C���c��/i�<	M�CMI;^8�<��������ѩ̼��0<^X���=��\=F] <��2=�Y�<�>�M^�3������;�:�6�M�h=�Z =)6���
�Q�E<��f=�:e<�<����l���켈��<��,�^)�< *q��U������[�ϴ<�l$�<�
�lT/=�{�<T�t���@<5><k�������<��;Q�
�>���?�0=F��<���<Θ,�:�$�M0B�^Y�~r <H�]���K=l=�i<D��<�:��Z:L�XZ���<��=� 4�ǈ�<�@z��?k=��=�l(=�Ԏ;vd�:�7=�8�x�N��ֿ<t|�>��<w�9JL��Q/�1c��2#�����G�;��P=�Hi���[��G\=�%=���o��A�<=��6<���)s ���0=Vuּz[ռM������<C[��p§<��*��8�<�?���؝<\1s<L^d���c�to��Y�X=�<�UL��qP�<eD��U��<:=�
\=�`�g�T�d��x
����
=1���A�<!2ɼ�Y9������ �VtG���=�'<r�h�#�˼�=�Q�<y�=��=���ݓP���d���壼��<Α�<ఄ<������#J�;�d�<u�U<���F=�(Ӽԟ;{�<�lL<~2�X;=Ɣ5��2;�v��J���N�<t־�χ^�*mV=ʟ�6J¼�:�G�jO�;�:���@���z3��̎�[mԼ!I!=R�<�X-<��Y�'��<��1=X�j���K��NO=F��[S <�<��K<v`�P�=�������<a;<`Z��L�<�T%=� ��m�6�<aRd=wm�<h�<�`�<�';=uh�ť�c�üF��<��Û9�3�����=�1�<E3=7ɂ��KW=+h,<
"U=�K=��<�����!<�)���'=���:�<:�����<����0=˫�<�a|���7��~���%<c1u�ﲴ�2�<0�H<��s��(�)����S�~�DMc=��'=U�L<O縼�T�<���K=�)�<��m=r
=���:�o&������?��&�e�j=U�y=	�ּ~�7=
$�-�<���VW���r=(�i�iT=���O�F��1���̼��j�e
,=��<B��<PO<�9�~����i'=e�6<����@=�n;/���^�<?C����;Ϸ9u1K��
���nv=��=�3:�s�9�&=�1w�N���§P��l�<��\�;�S=��"<�XZ����:� w��(Z�e��W׼j,?�J/���-9��I��>���a��QD�Ն�	��<x󶼐0=���TD=]��:�.ļ��V<H=f����ֻP��<.�켵z��#Q=ȺK=�<�5=�c/��!d=�n��:����z�J�n����<���ڿɼ��1��Q=�0�<��<�_�N�i<R=�=��=��2�\�D� +B=6L�<�f=`d�6:W=#�����<j^��Zv��,=���<�,=�a�<b6�����|A=���=�|�7�C��PV��u�W<�������㼲]=���me����;8J;x�ʼ�=7�k��=�[�7S=q&!:�
;�8G=w�{=ve=�)޼DU��μ~-�<+�'={����H��e�;�O��wG<����������3�Q�=|��4�L��=�M���a4��2�(#><&/=��:��1�~�E��<�4���a#�َ,�	<r˃<���<�f�<Mh�v��}�9=y���T](��r�3u���d=OѼ�h#�v��;Dk,���9=*mq<�|L=P�2=��D<��<��˼���� �Q�=��a����x�*��&K�#Vu��?=�TC=W�=P/>=B�.=,:�<�=K��<���5�i/�<�)	���G=b�P=�k=�,��3�%)t���A={7���L�^ټ���<��,�� =F�=�YT�B�����<��7��	��Z��v�-�њ��μ���;�7����<�O�:��<ܧ����;B�>�i����= ��<�C�'�D=c	S��C�,�%����<.���ǻ���TN�iZ5���;:�<ط��_�)���dc�Yĭ�E�J�����wb�䐃<�5^<P��o<�>����;��p��*���<y��<���>��;�L"����:ߥ�<I+9�70���;>y���<���<Ӗ ��n8��ۻ��9�-�.���ἂ+0���E=n�b	�����L��<�ͼ] �9x�"���_=PB~<���<w1=:3�+#��	=�U����<	}6=�8��sԻW���=g���X���J+<y�	�2H����м/Q� X�D�;�P�!���>�#j<��+�s����=./=7�<Ƽ=��EW4�J�< '=�'G�<tT���NA�~[�N�;P뺼ЗO<�t����m|�<v�G���8<!Ũ<�a����!��<0P�<����u!]�EQ�<A���0��$5a�	`˻��%��$l�梩��%<��Ѽp�<�RK=���<��(=Fv輥3��i�<([���^�� =�v.�2��M��鱼3�=�.=,�*=�[=�5=�2�A.���=ٌ�<{�7�a���ߣ;#�<U;X�g�5=����x`�_��< 2�;p�<_S���N#�����9�<H����8n-M�m%�<D�����"#u��;=��F=V��{�A�H�M��zY���;�H�՗̻�Em<v�=9"6<o�[=s�u<?XW����}����;���ˌ��M��<"�����<�+�� �<ߊG�zļl��M⽼H��;"�����;��Ҽ��U=@�ʼ����g�=cꮼ�b<�Ð�]k�;��O��;>輕1��i<�s�={�R=ڍ<�{;/�=��x<�!��V�LO?<K�"<4G=��q��t����;���k��pC�/�-�Y������7�<<��=d��C�1��
D�o�:&�E��=9=)�8��oT=�;�a�ny:=�ߔ��J=��<HO�Z7�W�8<���<{g?�J�?=ϴ=�J�2�*���������{Om=b�Ѽ�&=ʼa=�����K�b��<l��<��5�j7Q=�3�<
����^D�\ �<�N1<��=Yc���!�;1u=����$0���=O��M=�T�<�!�<D_<�߁���:J#7=��������;��<���<߇;�Q��鎎<��<~�Y<��h��<=8I!<W:;*-���h��{=;׻��]�=x=m�p�mQ�<��e�{=�n�r+������1ܯ�}��<5�/��Ba=!�Ӽ�M`�M+�<޴��=3��8�$= pA��s�� #��P�j1=r4=Gf��	W<B�<)=�<�=��A=�r�<��9J�H�_�޼cs��_U�ү��Ċ<�e�<O*ϼv�R<X Ƽ��4�wӛ��Ǽ��!<�O;� �l(�:�;�<1`=��V�m��g����x�<�B��l�<�t�<L�;�p=.Q̼��Ѽ�"
��6�<x)=&9Y��3�Hr-=4�|={�<�w�<S�[:��0=`�;
?�<4��<��.=�! =��<H���V�4�ko<��P��WP=Ĺ<���*��23=/��=� �;>�]�FL�=�P�<�L@;���<8�켯�<������P<���jT��dE=A�;'TK��@=��ݼ��=�:ɼ�EO�W�-���Q�@6=p��<;4�<&�e=�=������A��;cK\�S��3G?��뭺ja"�`�;�m�;�Q���:z�\��M"�P�:�/<*�ż�����'�H�0=��"�+}k��\�5��� S�;�<&=P<Y����;��<�_
=��<=��<ۮ$=�wt�䙌��0��9�<$��
�B�^����v�I��<��w<��;��	=t)5=[���h�<��T�_�E=sS=�'=�^�Ox&<���<23=�,=k=;St�����=����%;0�<�@=��i�{./�@��<�؄�k@J� �h<[��<L.�9��<�N%�xR3;���Y��E�<%��ȵ8=�l�<0?<��R���ʻ��ں
C軄��;y��:;�=&k=<��n�`���V�� ;��V�Q�f�ʱ��q>=������+3=���<d�2�j��s�z��d��ce��3���x����v&C<��=�::e6��qo5��a=c="�=:>����-��$�������;��:�+=5=�����$:d�=�ON��ԃ=���cB�<����'��:к�s�� ^<���<�_{=,d��7��z;>�vy=U�%=��<��=�H�~�;ef�;������<����=x��z#<g�%�� �䱸;��o=�xz=gR���1��ma���<��Q��~e=��O�:�L��EQ<�hN<2�|�wD��pM�QEn=:ۙ���z��!�r���jX�<U�a=��G�����I��1���]<tA�4�J=B^��F
�=�
�;�o��+��<#�R�Z�Q=hu���W�Y���RB�����m���-�;��Y=��A���O=�]<*<r�p�Jh{�s�`=��Z�W�<�!�u��1��<�����I��<T	q=��_���<p�=a㫼��<�4���X��(	=�=�~�<�����n= �?���)�+a���~�P&q=���=�uw<9���)�<�V=�e��<x~S�;m<U�<�@��'M���<\��tJ���Y{<�K���T�;H\=�^2=���t�}<�[=�=_2Q�,��<�rQ=��~��Z���=al����=Wa0�w�8�٠1��Dջ_'6<W{b=y�w<�A˼.Aຓ�;�0��G�<�Rf��I��1�<-��<.]=:�7��=g�5�݇Ƽ�#=��=Yխ<Q�����Ǽ�Z�<E�źZ�E<�P=�m`=b�<�k��m����p<���<l�$="AF�����9���6�)>��ҙ���=��=��<�<�x���q=~h<�";$=ø���2V=l
A=���3����[�t�\��1=�����&���6�C�=��<�/̼X<|���{=!�<=Ӊ�N�=1ҺJO<�V<�<�u�;�Aۼ��.=w�#�b�ؼu�<Ύ�<ͪ2�)�7=w)��p�K�`�]� �3���e<|�);��3��ch9��U=�=���|�;��t�<�^���=ۧ�<�����<�mA��]��?�<�>����F;�1���?=ƺ=yS;��E���=��<����?��:8��Rk=��R=(H�s�~<�&�<7�=�d~���n=D�S�K3��];��=��B�H�k��n;��*�::=5w���;DS��Q�Q=������6=�,X=���b�0�NvU=��?��y�<��<���]=��E��2�;�?W������Q���c�e+=���kO��RL����<�Fz=P�=�����M��k��)a������<�|,=!3b����j��=�<�Ӽ,@��G<�=�;z�L� �<��\=�m���ep=���΄��=��<̧'�g��+p���<�J�P팷W[X=�R&<=$��"%?���?��m`=��*=���<NGU�֨�;L�<i�Ǽb��:k<�
>=�|=�%7=��D=���<�pu<��<�6=�㊻sv��	��<�[�C��<Ɋ��ۏƼ���i=��d=j6�<ó�)��<�E�:c���m=]g
<�9a����:�����X���_i=o{�=�^��1������5j�
{3���78]����N=�m=e�v=w��h�<#�#�68=[�p=?a8����<E�� �-���=��;=��;<�U&=Ji�<M4<��P�M˚�D��<��A<;�<��c=�2�����==��<c�=4֯<3I�7��<�̼@�<l,r��|:���/�2=���A2p��f��g��<:�W��v���W=1kF=��a=$ED���W<&k<��t<�:t���=ԏ����ֻ��/=""�ϱ���� �HCZ�,=�Γ<s�ƼhK���>���*;Ȥ���3�Q ��߼$<˼�3�W�����1�;,=�ہ<�R�hx6��G�<,��" *��T�;���W{Q<V
E���a���"=��<=���;A7q�"���4�;�=��rk�'jҼ��ܺ4�9=)�_��
7=ʻV=2PW����d���T=1���*)��K�X'�D\����Jo<��v��]~=�u�<��z�*�6�Ϋ+��ĺ��>�¼�a)�.�i=oB�������
�JK=����@�;^˼��=B	X<)R�<?��<oU��|���c<
4�<V��X5���=��q���X�^��;/VĹp�-�����:9=��;;����X���l�<��=sS	�~;�;$Dg��1���<o�����e�dW��J�s�h�<u��<M+��Q�D=s�K�n���}+��qE=�K�<β<�ʱ��=M�`�{ܸ���n<�oA=}n�G�_<���<
�<�Q�����T��;uP����JA����z�<3��;��=�=+�;Ԝ���G=`&^��� ��.{=�=929ɼBp���g=1���j})=��9=�����<�i=DsL�D����<M�<�'1<��pN�<OX+=J�
�5��N��]�@=N��=��J=1���X�����J��;��=���*x=���=��׎�`�V�	���S�<�ؼP�=�=���AżFH=kMK<��l=|�u=ZP��g{�~�+=X��<p*�:1o=�Be=�)�,g�J�8<ό^���v��!��F�<Q�'��}R=��Q=K\7�d9=�޼Q�a=aH=s����K�u���N=�
b���Ҽk$=(&�+��:�<��������O���
=ro�;<�<Io==:�{v,=��Ի�gf��Ǉ��I�7o�<�O=ӯ;��<���<*�=�Ĭ��==�!|<j���<�!���)=.���������<������A<m�y<��N=ne<������	��'���<�����:ļܥ�Իû\_A<
��<~h*����}F���2��fj;�=��|����<QR=�
��o���(l����$>=4g�;��\�q
-���:��3�<��O����<�@"���:
`Y:^�ɻ�c����m����<n|���W=�`��/U�1 ��LeM�G$.=7� <T��G�F�x����(=����� �,*�;"\ҼaPX<��|<}J�;�Y�]P�=��ټ��m=�.��5��a�F�#��JP=���<��=1�4=�y=�tu=�wJ=4��<Ά`������uV=��W����hT��Dw<����o.��l�\��A�+;C�=�jU�w�:=���:/�'=��
��9ʤ������1��\$D��	ɼ�d��6�-;�b��[�<�hY=�B��è�<K��;G�$�Q5=�Sh=��C=1�p��.=a��;dr���<�E�<<��Ӽ�R�< �%�+���
��=IO�;��<�ե�]q:=;��0��Ԕ�YH=�4
���==\l�<v��<Ew�<7�=���3���
3=c�=�&�<m$���8����Q�ͼ �̼:��<���;��"�G�;�=��4=0��<ԥ�<��˻��/=�l=>b#�x�Q:�+=�E<p�2�<Y6��k����<F�a=�+=g$�<�Q^�UjP��������1����<�'=0��V��t�am�<��{=&7,=�e1��e,�Bބ:,�q�yT���I=1�<I�,;0o�;���<�aϼ�|�<�S����;̠?<CEݻZ;�Ӥe<���<bc=̷�<_��M]o=w�R=o��<2��`��<�)���j�;�^*���<�l�V�����v�䚍��o�<���<�.T�P!=��R�6Zܼ��><��<��λ!:<�IM=��:����l	�9;=�{ ���n<� ,=~�|<�=����M�<�!v<"*1=�C�ssk=J�<�r'���+�wwA�7�<#�=�W�Ի�%�;i�q;$9<M�P=ve�5��<@�=Ϧ.�cP��O�r��9\�d ���cb��w3<�uл� =-�;�wㇻ��＠$&=��!=�����_��Fʼ�Z=*?=�b�:�0�<b.�6E�GG���h=��\=l���B��T`-���W=؀=:uJ=��;m�����18����<���`����n|�L5C=�"M���<�T��`�A=�ʪ;�x��sA=�r=(���Zļ�����*=��<��<R�4<~��������'<@Sf=�&��A2=au=�AA=H4<��h=[�1��q�;܅���a�����;��=Hh�j@=v�F=���;mqP���?=~�.��ym=�\�<�F=��`<��{=�eY=�0���*<X	L��^C=̢�����$e��9�9�@;w�+=��C��j��z =��/;aK=c"�<���?O=M���=���r�pPA�U!��ͼ9�=��d�=Ƃ\��;9AD=oֱ<|L<��Sf&=�^�t��<�R����!�U�<�'�������ʼa���[=�'=��=I=ҝ���J��d8���
�9�L=�7����<~�<Њ&�\�/=��<��0=��O=e4��� +Y�o�<>s%:�E`��ů���y�D���$�I�,�?7�<��M=Q�6�Og7=ѯ�=�z(<SJO�o�=��o	=�W!:��d�,a<� =K�&�T	�<B ��<��[Y��(2=�Ї=���<��٘�����=\��< 1�;�
]<X-=<��=��/=�Vc<�:�� ��΁<��<4�8��K��:ꕸ;���<�E����ݼi^X�V=����q�M�==�Մ_<J휻��6����;��^zؼy1=�1G=��K=�C6�T���V�6�@�K��^=`E<a�;����<^V	���<��z<$�<��ἁr==�Q<�1=�Q==���!.�0�d<;�U=�eQ=u��<�pp;5��;܃1�z�r;+qV<Փ��X¶��{�<�	�;6�<�P<
C�<*��;�:��r5��s={��*]?��:X=Oǐ:��弸�<���)-ܼ�ȱ<���<W-<kv��\N�<���<~�i�E�62ļW@=Ld�<�H�<�l˼(T�<
w=����
	=�k�ߌO�]�����"��<�S<�yF���e������"S�� =��h<"X*�ַ��2E�<��<�v�<w�\���8d;�i�<z�<.�I=���y3�f�p=�����鼫�<^��h�ջ�FK=�1T=o5=�ĩ��S�<�h�"�<E^�Y�$=�ⷺ,�[<ln��ݼ���Z	=�l�<��>�2���Y��zb=�?���Z�P�H�0=y�v�SJ1����=�-=���;}��`���;�s <�^�������`D���5�%�)��J���h=@�:=f�<
�C=$��;\��<J�E<%� �r�<���;K^����=��1�[6�</0'=�U�l]x�Y6�R?��4=��=12.��X:
�o=��鼯C��5"��<<ԭ<R+<���$���߼W�D=
^���˼�IS��O=�g�;(��k��<��I=��:v�5�Ҏ��N=H����p=��N�x7�<zW����"=?p漥�L=~�k� ���r��T��b"�<
aj=�̇;j�=V� ��Ϻ�=��6-C=i�-;YC��Ӧq�"{H�_Z�`��&��<�2�<��C=�W���˺pz�<��]�<�XP��٧9@2O�&�~<�+���c��I��<o8<�=�	=��_<ޡ�BV�<�5�;�7f�3�XF^=�鼓�N��$<�䰼�a�}�V�J�;�=��Z<pQ��i�<��9=D�Ѽ��=t
�YL��A�<&Lb="�:o8F=�5+=)4�<aIj=�P�������W`=��=�6=��ۼ[�<�oϼ�p�����켯vN���6=�Cl��9ʵ�#a"��ۦ���F�Ǐ9<��U=-�}<�7=�Mi=8_����ɕ<�`?=�~ͼgr?=����d(<"�����/LL�y�:�������V�j퍽5F=S#X�������<�r��=d��<��<6H*<֛=��^��6��ݺƷ7�''p;d4�<u�2��D�<i'���A=�/�uĻ<M"=�~A=�����
;<�d����a���<�vw<�Ǔ�-����x�<f��c���2�Я�<~S=�8�J�Y=��?���V�~���!=�tY��{�<�Vo=�0���<J\>��L��+���]�<6�_=�\�<
m=���'��<��<\�=;{.;�I����f�Z�+<�<
9(=9J��?;V��<��!$�����n�t=`q<^��<7Z��
��;�ж<�R������}G�wp��A�B;�g�<�lM;	�6=�<�C=EJ����/�1<r����?a�rS='�i��/��~�`;�X=:��<)[=}B0��ph=��<}��j%�:�vB=G)�l,�#W�2=-驼� "�8�<��:�����3�b�!�jպ��K�̦'=۹���:i��}s=������=�S)���<o����<C��<��<>��9���;&�<F��ysW=�'����ϼ�߼��
�c4=M�<q�<�����;�� =��<�7-�s�L=��K=����9�C=��0���ݻO<�<
*@=��@�4����=X�����(�PĀ<t�<�~�;(�M�G,��T�����;u�=��Y=�ړ�7�y;_��<�/��x�!=]w�<M����u;��;A� ��S[=�P�B{��$�<C{"=�RQ=����D�a#�� R��mb=:�=L6=Y^�<�D�6C��ʟZ��H9��H=��;��;�;���<P�[��Va�Y�<µ�8-�=+$��v�ƀn�p�����;2�<����V���˅���6��J�2���[<���� #�+,e<�T<�$=�c��~Z���&��3m=O5��MQ�� �<�L��Cf�*聽�C�<����K������`꼋���kM�g�@=l��iw<,�=A�-��6Q�<��V=�W7��uJ=��<41�����<6�#�)���޼�6ʼR�Y=�쵻�m=�ā<}���`=����� =$�"���<t.R=��-=�d��V�f<}�%=�!���8y��-'3=��P�#�-��<rw��f�=)�<��=R=,˵�:Q軐��<�O[=��������;t !=6��FR�+��:����ȝ;<�4=%/��M�=93z= �g��Qy;뿝�?_�<9n�<��<��<hi�!L=_X���4���*�<O��39�;�3<��A��z���=>��C���<-J����k!=kr=BlҼC2�<� ��*�󸺼�Ė;�7�<�&�<�G��6*<��D� -�hH=~xj=*�(:@B&�%��q�<s[�<� �����-I��Bu^�-g�<Tb�罹<Ƭ7��O!���$=|7g�Q�[=q��<h��;H�ۼ=��`�=C� �Q��;�N=&n	=�2;�F=$��u�I=�_�C�l�<� ��i	�����ڦ;�"�<9CN=
w<7ve=D�� ���:+=�lN=��=�V=<�s�o_m�o@�e/��eӃ�3��;F)�<��������J��
P�:*�����;3\�<2�~��،<�dA=E,=�dg>=��<�ׇ�*&	=�2O=�h�=�8<Ѿ��t%?�T_�@`�xϼo�!=�*��76��`<��"�#�p��<g,����<ki=2�=�Z<���۸<�-P=4�}�w�I=�p��gg=��o���U<��ռc�P�!x==��4��W̻�¼j�< a ���<��&=3���:��;b��<DƼ��|����;輼>����*p<��y��2,�]9=-Hj�����-<v�"��3(�&),=�CS��@=�+�;F�#=b��<G����5D��$�+�R�M�A</�W=]�˻�C2�.u>=P8��=U�;̴<�O�7��:VI�<[24<���UA�TX����<��:
f&=��f�l,�������f<v��UN��U&=A���"=!~1�B�;��=���<�Lu��*�����#�<N7 ��gB���<��;=b�<##��<�|^6��,��{�<��< Z1=M�<)ޭ;�?��Y�����������<_={��@5l���#<C�=���,���K0����V2���:��J�c&��[y�:u�;u Q<=%Z�XZ0�t<�>��K����M����<VR��\=����n��< ��J_;�t=.�;tԔ��F<�~�<��b�U(>�� �<c?$:E�=2��<~�ؼw���p=@f=r ��ʿ���<�:�<?ǘ<7#��ݠ�L:<$x�<�
5�Q��{5+�p]�X˂��	�< ~:o$�<�?�<�o�<��==�����O=�0=�]�;w�<���:-�?<�L=����h$�eE���%=���W2�/�:9���;u�O=�'q<<��;M�ռ-I<�cͼ�),� �"��<՞<5�$��P=ҤW��*=a���ܽ<W����4��(=�}��[�CJ�9�Ka� �F��;b����K�r`��+�M��`e<\�|=j<d=DSE=O�U�xo�����yt<�"��fg)�}zF=	<�5]�P_�_}==�,=�9S=c�<��S:�5P<�2��/�.�N�E�@��1����6�<�>ټ	���9d�[KP=ww�9�h��=��\�X��=x0�<�U<��/���=��<��;�;ڻ,h<^}#�$�=����?���<�9��oF�aM��*=���<�hN��V���T�;{�-=�n= �<=V=c���9Ɠ�;��<��|��$�<8�<h�!�nỄD!=~|=�<I��r�3%ٺ9�s=&P�.}H=�}�<?�4=s��슼=�
�2Q�0�<�;���=ҡȻ�d ���O:��ݻ��`�P��<�-�p� �s�$=�y��:���V�.=���c�ݻ*�� R1=�-=�;`2��]�\<}q�:�/ڻ��I�F�M=�a���I��C�¼��<�py�#+�V�^�X�0�TI�<��<j�B<B#
;��E<p�E=W�I= %(�b��_�,���=W�L��<<��F�T_
�i}��ү=j��G,d=��ڼ�[���=����A����|=t�<��{=�g�<�ͼ<e�V<C= �}=?�����7=g~�<�!���8���<�����l����=Xi=Ԫ=G x=�a����<��Ǽ<��U�	�X3� ����2���ᴭ��թ�=|v��2 ��	��}=�.X���j=�
S;��/�~j><�o�Caw=��<=c=��<��ػM���	(�H����Q�9<�EF��2=�l=nf!<#19�|�G:����~�=X�Y=5Z漃6�<3��W2�h{=���HP���e���VF��'=��<<����<@=Rt7��)=盐=" μ�X���e�?��;��r=��j�%�'<��-=���, <{��{�=�K=�)��K����d=ϼ�h�:L���}W=e�;J}��� =e�W�*눻��/=:��<{>��+�=��=.�/��==�<
\t=sT=�a\=��r(=��U���x��߼+�E=��^=�R��X�<�K�<*��=1V�"�}_=0��<��<�i=�Y9=ny=�fy��}м��*=��O=n�=�����߼'����ݺ��ӼB����I��=h<
�<a�W����s���`���W<�����<����O�>�=$��;���:��<т��ݻF�h�4�k��׼�C�#�<�m��]�ټ�%<=��;�_'�����=���= �ݼ��mL�<)��X�;�(�#�a��8�j�<�	��;�����c=��X=�+A�L�#;�{=gא�%��<:�=�y<=�� =N�-=�?E���&������=wG¼S�;�;p��^q�V�1�\}{��	��$�<��=��+=N�켐�(�j[ڼ�A�ė��S7=a�IC=�f��.=��_��	�'�.��&�P�2�M�=F��H-ĺS�<\F4=((=#=���@�Q�]mQ=��%�P��x�����=�\�<tߥ;�-<��X�{�$�`&�<\�Q�T(v=��Ҽ���
$����E�e=P��;v�<���<�NS�(/�G�=�󠺰���5�p���ԼQ�=�O;�;��=,�^=�C=�OB=g�3<��<7� =ݕ@��,=�Q�aے�pnQ�s,���c�@�Z��<�0�<�����Ge��a��ox9�Ы�u���+�w���B�(���6O<�=���%<�J�<)FA�*�-�t�߼N���wU��!꼶�=8R����<��5=�r:��*=K	p�]i1=�
=�5���z?<�=a0ɼ�E����ļ�<[�{��0�<�-x�d�J�=�)���<Tf=�g�<\c~�f�s=WoP��r�˜�<�닼��7<�ݘ<P��X7=�7����6��9=
Z��2^;�'f=#o��2�;O"j=����߼즖<��l�xx���3$��<��ռ3o]=]n�=�Ӝ���V��('��{=����3��<!�!��r���|<F\�ܶf��l:0��^�<|Vh�'�P���H�����Pt���%�A_<�#a��M6<�"���<:R�K��<7�%=�=HY��>&�0cV�?�Y=`�=��<�@�=��<g5�����ݓ}=7�:-�<��k=�՟�䊰<���<��Z�yF=��=���<��1=vF�(�4��*���A_�x)�<���;^��h����S=�Ӥ����<*b\=�<=0E1�$��<H�Y=D�<)k=�:>=�V=� =�i>��즼��a��:9��a\�<�	�_\�<Ba��=�[=�i=?ܥ���	=y�j<�&��k����<��V�o�#=)� �H<�AǓ�.o_=�����`o;��=��!�������X=X�󻪼==�<������d6=�S=<.���%.=�5�<�Aٹ��A�`i��V�
o1��YN�9�+=�L�+@���(=!�V<�<v�z���������&�C=̀S<�g�;;�z=�c=��&=NvҼ�^=����˽<<�<d��<���<y䑼�+?=N������"�ͻ�V=���<�q=�C�̫��x�<vX�<Q�s���q=��S=�.c<ٳb=
�=�[�;�%{ļ�� <�n=I� �I�@=����j����3�ǧg��4a<{ɴ���3<*��;f�W=q�u��(�l�üN�Y���	=��{=���<"5�<�����V<k�?=��<A�G=�Hĺ���<B,�����F.����<��;KL׼U�#=�l�<�Dq<VN��=�k5�O��<T�f�W�!;}c'=6MC�B�=SzX=���<�2/<�dc�Es�<�(��d_9���;I�e�&;

T��:=�a-=�e=;���Mb�P�m=z�F��}�<����L*����r��/���#�<~,=;���pQ��� �E?=��<�}���{H=��v��CR�k<7=2U�jX��h��n#=\�V=<�<%=��z�G�#Vl�g�Ȼ�a��fh\<M�<�����������<�����=��Z�1@���H<̱l<�*����
���ż��'��Y&���I�X��D3<yLz��"лjX$���h��IZ=Y�=#EH�SU�< D]=]l�<駁��?��qz�<8'�<Jt=^Q=��=m_�a/��:=�[;r4����O�%�o�'<��P�l�C=cw�<���2�=���;f�0��b7=+N-��G�; =�Y�<��ؼ��O�"j\�:��4��F�H=6a*�0������R���E=��Q��VB<��F��:5=t��<E =�7ü95�a��<�w���<v|�fyT����;m4ü��Q<��v����;�;��8%T�Z7���1���<	X�е�#%��=�U���$����<�D<��=�t%��H�_~=;��;o�,S;�?=��<�q�<kX|<��O<�@�U=�p�ݙ
=����v��MKd���!��0t<�G�<sg�x�޺vy^=q	G��E&���8=^Z�y�<r�	@��sB��S����<P� �i���<;~=�ޫ�����;b�S]$=�D=�k�1�,<N�$��<_���].7:*E=����pO�� Q��һ���;����
k�������xw����=�
�5V=� -=c�=�G����w<f��(zP<��K<���;|:C�ZV����@�< ��<G�x<�-�<Y���f���7�;�f;�=���<������===I�S$s�
��N�L=�{��~,==�G<��<����<��C��3==��	�r)�<��=���<�[T< t¼�_:=����S�K��<X�⻢�G+�:�XU�]J��M�0=�-�ʡW=��Z���H����<i�:��!=G'}�B4r�!=��<@�<�H9�g�,=�]s��qr����<8��}�e��m��H=Fp�<�^�<�F.=6�[���k=�+�<���<��/��&�<'N�f��<��;6�h�O�[=&y<�L���P��D8<y6(=d�L�p!="���~S����;�q�u�
=�,e�ق"�}�/�>M�<�,��h<-7���S�<c���A�<"��<MHw<��;<l]��K�;I[�<��F=}4��q~=��'�P=�A�<�P<6#l��B:=�wP�I�O<�[D:₊<Z8��,==����<�n��GYk�	�V�T}��A-�7~<�K1�9�[d��	B���
=��<���;'��<�im�K�@<@�/=T�G=U̞<>N��ckN=�n:�3�!��`��<�x@=���<�;=��?��	�:��i�����>`D=椦<%�R;|�=fo�<�3b��3�;X���n�=���;�]�:s=�Z'=ZrY=���<'IO�CP���S<�2�0I=n8��|-5��x<#�^=S(��e5��쨼�%s=�� =�1L;�e�<5W����f=c��;=��<#�$=�%�B䛼�j3���9��a�,��D'��::=��C�v�?�S�<��6*+=�����vl=4J�<m���w|^�H�<}_��Ņ�	�A=��<�i�<�1�R�D<�bS�&+��eo�e}�am;Dc=�#t<2$�ܡ�:+�H=�S=죖<��l����<&C��3s=ƽ���)=���<b��;O��<|�����J�=ر�<M�_+��� =Cu�-�=�Ă��q��9��X��xd�<uN,=&o=��(�ƒ<-줼� ��R�;=�;tFR���%=#���l0j<]U�<�G=ڂ��
Z��_E=�]��U<�B=����<D�e,3��$`�!�F=Y����/�<���<Xb������L]=Č=6�A=L[=������O=?�<�/ڼ�2+�X�D;��<A^�`<p�D=	��;u
�;����c�,=�[=#Z	=��,:Q�%=m�:��żX��=�l�;D/(���ɼ�B5=KH�MC��9q���=���<Xk��Y�X��Z�����<�cP�&*(=�.�Ǖ��p�?�Ԣ����=�<o�(=X�W=M[���c9���N�W����<ܕb��Y�J�	=7V=k��;W ����J�G��<�= �X��_���l<�"=��=�!<����]�7�0�ɼ��(;���<p'���'��1�;V�ǘ����<d"����<;]C��c��<y��i]<ǶQ=/AD=��="�<Z�+=�/�XS��7�E<�J���;H�;������=*�GNY�٦���ͼ��ּ'����<��`�c���q��;�"��b=��E�a�E��J%<9�A=Q}g��<�G=�!<��F=�߻b9/=�4=���<�*�<�#�:O��Q��R*ʼBˑ<�<=_�;T�=�b�<);=ļa6�:�¬<۠�:C��;StH<���<�j_�UԻo�K=�l:���חo=�#m�v�<E��A��������:=�GM��ہ�fɪ�pO��Z�<A�<�wb=	��.��Xh��O�����|X��m$<ֲ%�r�<�N5���;��$=.�4�q⻺ ��m��<�BF�"?=������:=��U��9�E�^�>��^�L�o�A�G���;=�{'=���ՠּ��`��)=�$=�Ub�l?�<�yּ��<&w9��gۼ2ׇ<C����޲�K�����J��-N=�(M;N�����D=
����Ʃ���rx<:&_=�?G<���b'��ɶ<$8��c:�q���rA=��=䜼<};���3{=ƤW�W导�>Y=�j=@��<�ݻ�B��<D6=��=�<�;|�$�uT�<#�-��#=�	�:~�5�SR=��*�B�f=@ �=ȷu=��'�f��=�U���w��c��<?X�<b�>�%�`����<��#<���<T��<�'<�ZO=����a+="�=�$�:_��<��i=���� ���=J�ؼ��<:�>�po�=}� ;�W�����<N�\=;-=���S���2�r"=���<��"=Tlx=��<�1J=x<�<��	�۫�>9U���9=��	=kѼ�	�<?OV=گ;2'�g7�	S<-ij=���Mw��l��I+=̚�Nk�L��<pʧ��c�;@D��v==h)=��;�C�<�0=��n��M<3�<�<|e�<���<C"B=)��;�X�����]c���	=r9���맼G�/=ц#==�s#=>B���*<����9��ވ;�YR�����������R��C3=�Ƿ��Y�"�<]
k<�=����7��7<\��b�=���W�\=�ǫ<Q���I�<�P�P�ͼ�Ze=o�<`'=��?<d�~��F�����)<m�F<$K���)��5�=w@=�@=�,�<C��<�Ng=۞%��.g�c=�帼�/�<
���c=��G��'H�<�;� < lż�ʟ�C��;���Ò=?Dϻ�,�<XfP=�_�*8h��A�<7����<�4\�m�D�
HY��^�<�\�ЪJ���9<�	V���V;�G�8B����������;K���XW�<̟*�pMH;5M������=e�:�J�=q9X=B�7=�*=U��f����6�<��<k'B=��ϼ��u��3"��=�_��8\��m��=��,�$������;,@ =8w�j�@���<~�K��r�<�pW��j��u~���<w�:=<T������*�Gְ��
ڼ2`�&����� =_�:.`e<�8=�������� <!gz<�ق�s��}�y��9�=�S=zEƼ(�<n���\6�I�;��=��h�����p1�Q,g=���/��9^ڼY���d��4���/��>;�H�,�B��<�ټ�CC�j+�<R����[;�M@�!c=N�<��;�wS=*��<'Z$=
�;�$=�UY��N��f�<u ��bA��Z<\�#<��\�$Z���B�;2�5=��k=�C!�}o߼(�e�;��<ݮ��l�<�L=��}=�� ���=�t^<�;��k�<Q� <K�U=�\���D�ߦȼ��3=2!��~�<�_<��=<���N<���:	91��V��I.=��=�9=j�<j��Ž�<�H;~�:�o�|r�<��?��?4�L 	���[<�T�<��e<�}�L���^�������3ϼܡg;9 <�@���(;c}���j�<GL�:N�=�%n=h;Z��<w\R<La�<�9�ꋈ�n�5���6;ҏ����{v�k+=�0)�z�t���= S�<N�0= �6������0=�D��7��^���,�<�\R=���aF=Vt}<c�N�س�<z��;p`N=b�={�n= �d��úB�q���8�;�4���1�@m�?2=c뾼=��<!�ٻw��;|G＆P==%F�����T#=�!�`)��DH=[>=ymE�!q=�vA=>�*<�B��or<t(@������=�:���W=ru3����������,Y���<����U�Q��<�5�W헼������;Wx�<�	=�CӼ'Je=�@P���-=������{'T�D�n�7�j�R��<t^Q�I�p<��;=nXʼ־�<��*=�N�o�o;ˊ8�h��]x�pů����]���@=�X������=պh<���Z���ZS<|8I<��;�9���͇��S�<Gt<)�#=���C_üJ<�<�o�s�?��ぺq�;�/~=�� =_�_=?~A=��ڻY���$<G��=���<]��<{e=:5o������`;�������'B�ዼ��m`�;]Ja<�0<�	���y�<?��;�����=�#	��f����˼QX:��	���.�H��l�<=\8�\y�;��?���GR ��I �q�ǼK=��;K�l1(=�U<�gҼ�,C� Ǽ�y6<�rB���<��<=�n<�D��U�m1l�^�!��\�<b7M<̗<��<�雼I��	u�<��ѻ#�3=��=�����#=gk��@<��N<�~�;Yd��	�������o�����<N_�:�4=%_��=��9=��O=��=��%=æ�M�C���n=�����P =�=u=�<�u�<���/ `:(�;�`h���~�;!熽�
=�ܠ��M<=�V=�8m�^߁��{=�_(=Т�T�
�@�e=��r�&�"�ʀ&=E/�8N=�$o=A�=.�=p���R����;Ep���ڧ�;�W;E���,�< �׻{����} =�&:���_=KI�<_�H<@Z�<z��<�=���E�:4/� �z=[���z���\-<��P;�y0������������ �;6弑�=l~�<@��lj�\�;�=(=5�i���r=��<�˻�I���=3=�k���,V=T��lo��!w=#�:;LV=��V=�� �G�V�cWr=���;Ca�"�=J=$�=�- �����<�u�*���>�]3=��+=�vT�.9�<
E.�q�P=�&@=�u=�U�<�9��=G���A�sH=��;_
.�n;<а�~*��4鸻\��<�<����6=wl�<��k=�R�'T�;��>� �$R��WE�V���v����:���<ERZ=>_=�j�<k{�<�����,=Ȕ
�1=�V�;�#=���Ҏ_=S�5���'�BԼ+ɞ��e%�(	<�^t����"�_=zrؼ���m&#�{�"�y�;Ir)=�j+��I����ʼi� =�W����0<�պ�s=8�I�8=adm�ْR�R���NS:YW=��7=�AR=i�`=CmK<mǼ��;豮�%V�;w��<�~�;k��<��M�|0�<D=o=G�A=V��;=��:�G�>�;�-�H=G����	=55A=��:-b=lθC�<�+9=x K����:g7=-��� _�p�%=�R<�b�<ҷS=rm<���`�Vt����9+�n����b�0=�w�;��M���t��V�<x�=�C=���<em��Q5K=/ȝ��
�aV��Wo=*7i;��$=`��<-.�T�{��ܼRcO��G�;�r�<��4YD=/׻'��<�'?��;�y6�e	�󩶻9\B�::鼛�B=�S�<ؼ�Wi9=�_B��b���=x�Z�ጅ<0����L;Xx=3���gRU=�@�<2�����<�B-<G�a=��3=��ź���;�YV���.=#/�<���S/B=_��<��;����?=���<QO=���y}�Z�<���<���tڕ<(X7�ǎ<\�^��3�F>��Ι���<߹'�.�<AYZ��r�=E3={���T�;�db�*<kg5;�>��>l�_~M��/=<�*�	=�V(<���<����p���1=�i�*I^�3�y=�.��|=����=&���p溨�	�����=d
=3�]=��d�kH(��a�<�~=,�������e�;G�x�򫷼bu>����~tw=����Cּ>-���9=�m�j�w=�J���X�x�<��^=��)<Y,�XT�<c����I,=��&��{:����<z�I����<�B=oY='�<�P�<у6=�[j=.�=h&�;�L:�Z=���l!V�[�/<��b�D 9�G����.���>��!V���;f����!H����<Y[�8kȜ�B��1��s'=��x<M�¼	A�&�<�h2=�A=�e=��<>-��i�/:p�����y<�'_���c�Z_��<"=zu=��<T����̨<J
��=�f.=��<��<�����[=P;+��I�<?;<n�����
���=y�=�
!=,��<�q�Kп;ox�<xUj��6R��Y��@�V��ћ<F,�<Al�<G��O�=�΃=$֑;+?�;9=>`=��������;����f����<,d��;,��7�<��r�E�6�f�w�i<�'�;�n�9�7��w+@<��?m�^�"=��a<��|��k���f<��8=f!#��>^=O���X&l�Q�D���_=Sz=�l��Q�(��<��R��m^�P{�*�X=Ȩ/:2=��<�js�n�n=&�)�?T?=�-��٣�<詼^� :�s9�u�k��Kr=V�a=;��f�"=���e����dN����z��<�0=K�K=S3^=�$�<�Z�5�5=t�;���<u�=�6k����<�7ݻ�y<Ku#�L�Z�@j=�N=��<c��<�,�=��<\F7=�R���d�<��3<lJ�u4y=�9F�i˘�����|��E=|F=CW�\�%=L��<H�<&�؈{�1?O=L�H=%��ėf�:�7=��-=/;\���=VG���-`=�!|��g�<rݥ<�Z(=A�«��<a�h<I�"�=Ͻ;���< '�*d���j�(x7�\��<�0�����3?�<���<.@<tP{�-G=��d�Z=� ;$�y���%=�;J�KY�<�ǻ~=�l���VL=��&=z��<�F�<l�/��X=��F��'¼���|=��Z��؜��M{�0,�;�C�)��4�<Qʼ����C�(��L�p�+<�DA=%λ��-=m�=ܺ=1�<j��Ѭ =���<�p=��O�TS������X=Y��Wm�3w&<X{���߼��J�:?��(���ļ���<p��<��<b��9-Z�W{=�dȻ\u5<���C�A����P;�<��=	�仴��<��<� =�p��X�DQ=�c�j��aIl=��U��S<=PC=PM>=.�\��P����2=�{�<U�<�	&<��=y��<ފ<�CW�*:c��Go=���ŻX�_=��$�ݍ�?�= =�<��=܊C��&�0[;��&=�����b7��D���-ʻk�[�ǐ<Dd=�R�����F����<�vn����<Vg���b=_����9����;�6=ļC6'=��=o�<		<!�J�Us=��T�%L���Z=�D	=���wy��ɕ�e7==ٺ9=� p����9w=�~h=�?�Q��<.oc�X4$=�Pa��6�=J-=6:<<��I���1=���;�t:�b(���==�EʼS.y<�1H=�ռ�m����<!>4�0A9��
��+���ͼ{�D�97;\(5<ǝ*�:A=����R�8�7�x�ۗ��ZK���Q�1�<a��<7.�<3�^=�:�}��p��<b*=�~�t�hTE�8��;}]=��W=�_!=�6�s}�;��<��<�;"OC���<5"=7"(��<=kbm���A�'�6�i��<�R�����!�U=�|��м�ǎ��\�B���I;=�e=q�J�0J�<�.=���<�"�2��=�z}<ج�<1K!��m�<B��<PID��M<���=v���(=6�a=�<�V5�O�<��L��hH���9k���>�<&H�Т%�����C=j<=;����=&q)��G�;c��<���,�i<󷲼{rX=:�<�F=vSw�$�ż)�8�������<�0<�� :R#=�*���

<w7���<C8��Fz���}<�=�f�<�
#��f#��C��.=�I=�\-<�&=1�<�0==�y<h�s�w�]�@q1=Of�;���/+�2��:4�~

����<���<׎H=�90=�DV��1�<��ʼ(�=L�Ӽ~�=�[����<�wV�#�3�FѰ<ş�;O
 �7��9�7�� |
���<e#�\j.����xU��2=�b�<`3(=M�=<S|<��e��Ӽ���;�;,=���;�25��s��ؤ`��}<�� E;H�(��Y=��3=\e=��8�v=�xܼH�<��e��Q=�5��=o<1_<{'0=t^�Ȕ���V=�Y=�v伤A=!%=�!=~�-�ĉ���B�&����<�$�0 h�w��<l�9ig�],�=����d ���d����;��(��f=)�H=մ�<��<5�����$�8N �z������=P�=Z��<��&<��"=&�];h��]@7<A��;=��<��9=l-=]/��
ʼ��<$���"��;��f��;=�2�o�)=�-==ݟ�g��d�P=Liv<`��;��2="ڮ�$8�<�=��)=�r��"�����/��IT�2N�b���$<GPD��E=-><WN7=���q!�;���<�I��1�N��<��=rm�έ�<G`�m�s����\��K*�#D�!?=�M/�j�.=�!�<̲
�҂�<#?)�8⹼g��w��<v_<���~�<$��<-�9��/;
b!={�ɼ�*���<����M3=�RR<���;��5�/X��x=��=�/�i��<�[�=hr��Fr���@�&q�2��q�<ߡܼ�gt��.M��9����d=N'/��=¼�@1��޺����<LGQ=�<X�Z��PC=h�Kμ��G�gE��T����ֺ��i=���<H�;�l�-�}����<A`8�9�	�)��J�P<ꇍ�� ��k`<X��;���!%��@��]�+=�L�����<�s<=9�<��N=x�-�
I�6�;iUK<���y;	=�iE��#�<�i</��y����W����<`D�6?�<���<BL�<1�P=�6=��<����>=t3���u<j`#=�A=�=a�;��rFf=��<��<$�<�5=��i�	H��?�J<4��<+��<��v����uҼ<��9��:0�X=!�$�U,�<`an=��h�K���=l�"�~��<a|=GӺ��#�1�=�s�.D=�H�<�T��9W�<H꣼<ۯ<�;�] ����~�;�S���Q�$A=�@r�A��;��<K=o؅�痲<��=��;9Q=���;���F����Y<���<�%��s�=��<�+K=���<B�M�;\��%�x:<ʆ3��w���bI$�[�g�I� �ރ#����=�Q�;�S6=�҇�P��<��=+b7�c���d�=R(��3�����<��'�)w<=�l0���X����<R�J=�ӹ�2,/�QCû{�J<P=��9=K�<��<�뀽e�=��=�z-�Y�X����/� �bA��k�:�ء<;N:=�@��ն�x6<�3=b��<hTJ=�E=ЋH<���<l<�y��Ա<};]�j�==T�J�Xϼv�1��;���I=Q��#ɍ<k�`=��6=zfG;8W<�2�<�ۿ<P�<�=!OռO;5=�,=�H�<�6��@>=��=m��=X�c=���0�<� �+ܛ���@;���<�������߼��/1��;��IT��)�R�<�㼼`^�<>/]�p-�a�=ol�<w#�;��<�'����2=�^%=�f�<�a":}�I�d=.i��!�<�1}�9!��5�%����U�P�d�^=��8�+!T��S6�9<W�&��=.U���� -:'�0=z��ժ�<��_�K=���<�=T�6<��D=sC=��*�ېu���b���-=өD�j#��j��P���	j�E�>���_����0=�ɼ�
�!=�W�FjN=#��}�?=s �2� �� <��=A<����R�,=���H%!�w�,�T�7��E��:�E��Tռ��>;�8�KJ5����伓R�up�<�nӼ�SM�!e8��z�<�w;�S;���Ѕ=6��)��������p<K	a;
��d�<J�}�<�5Ѽ����q��ObF�%ȼ	b�<ɕc=�fR�!��<Pp@��h;�V���<Rk��2)=�N)�h����=���<���9u,��p���c���F�d���.T=�?<ɒ���A�?�,=3���F퓼R��:,��OO�=cT�l;_vq=���<���<1D!=�7ϼR@��:k���M=�{�<��\�L<����jػ@�����w�_��O^�r,?=>�5<��w��qϼ~���{�<�?���H�מ�$9��\X<i!=Dӆ<����<��+
ɼ��v�&)=͓@������&�&��^�p�<�m��Y=46`����Fw=��m�@����L<V�;R�ӻ�)���
�{g�<2�ռ��=��F��Ӥ���<���<��=��={ �R�4���%�����[�p?=̷l=��d󏼓�(=�w���K=z
c=N.�;j��:@5�����Ǽnsa���ϼg�4=$�k=��=,qN<<�����V�VY==6Ng��c�Ic?:�_�<>��<� b��W!= ����¼W3N=*ZU=�=�*|����n;��&=�4�;��2=�0��>���d�,g=�.�˃�<��=�(N�qu(=��-��6��?
]=�ƼJ��<5s�7�<)ڨ<~��1��r<�<�j����μ���c�]=J�t�fS=%T�;a7L<]?2�DO�8�<�s=\I�� �0�7��}��.�<�u�8�L��<�'�;n���j����<�o'<�/���aȔ��g:=0u7_y�<�z�g^պ���<�8�u<:<��p�}<�:�	��S��)�D��<UT�]z�����I<66�ID`��� =�M�J_����֍��γ��� =-`"��9[=F ��1�=���%�t&l��HG���=H�=�g黷 �;cd���=��<Z�j=fw��A=�=���<��m=%�T=ϧ�g�p<���a�v�W=������<�BS�u��W�,��W=��;�=�1=�<h�~�h�q��]-��i�F�*<'�;^˚<}�$=��"�8�-�:WH;�=�8G�=k�8=�]�2M�=�%0=�������Z��;fdX=y�0=�*<s�G=�&�<������[���<��<�k�<碢�����י��M�z��{��<�u�<����fQ=�u����Q=\�g��{<#�a=��
=]��<�����*=d`�:!�:���<�x=��J<K��-p`<|�<+p��P2����;�8R<�I�'�+=0�t����_�j�0�Ҡ���=����S������i�����=/�3��g�;Z=<=s�3=�y[��?��^�D��6@�WR�<tcR�)�<x_�;Ap=����}�V��e����<���l��<Ca��%�K�=��<p�M�c{8�i0<4a�zE�<�;=g������r)��/��:�m<:��<�}�;+l�ӥ=�������A̰<���<��<��m<�ĉ�ߵ%��d���9;=�ϖ<��"�T�Hw=�ѷ<�+m�m:=|\+=5�򺭔��[�W���#=�h2����� T�Z���������<����4�=��ͼ��=�!�<И(���/��ѼVi"=M�=�'�i�[���9�ћY<!P���8����<I�s=���<�o��%T�Z�C=���<��l��`=������ջU͔<G���"�-%���9==�K=zp�<�<�a�-5��핼���w�e�pG9��""=�E�{��<�4<U�<f�=�4�;��N���?��qP=�=��F=BY�<�c�Hg3�y<́Y=�0h=P�:灃=��ȼ��8��mh��qм8��<��=1��"�<�.���E=��	=F�Ȼ�G�2򔺽{!�H�<-�|��Lٻ>�x=8͐�xp ��d=��!��}Ƽ%�=�V���,=Օ;=_�g����,��pti=�꿻�� ��zkr�oS<��+��zV=A�	=9�<ucw=5��<�z��Si�<,�<{&�˳}�m�D=�n�<��@<$�,�2=�}�O�H�p����d�Pϧ<+�%=	|�h=�k�]�D��C��a+�C�
;�<��=��g<�9t��]d=�BF�����J
�;E���:=��=��8<��F��C����+=<�<�rY=ZL��:A����׻!�K�e�=:&���i�uS;�t	X�GjW�^�n��}=��d=�z:��Mj;!�~�Jr/��vB<���;ZT���<�=Jg�<���f����<��=�kZ<l�)���<��=�	�����<7D=�iL���B<��==��%=8
i�m�4=��3^=�q���G�#�4��/�;�b<�0r<T�	������L���.�V<;�<�=�?�=���<A�@�i�<��Y<@#e�� =8<"=rO=���<X`2��w/=����A=�_T���K=w�2�6��M_<3�S�;�<n��H粼�Qn<����0[�QO<=�dI=�}���k�;B=� u����<�P"�[�R��$/�%= �<I��<j<�Og�ױ�<��}��y�?=:@��RO}����M�����Q��,� �<c<=��==����n4<�A4�ה�<�K���Y�cX%���H�kE��2�u=;���#+�b��<¼]�Z�<wNA�����qB� �U���H�hY(=��3y5���A���=�=R�O3��J�;QE�FĊ<z.�(I����<�R߻9�F=%<=�r=m�(��z@=�u���xu���Od=M�<���<Wx9=��;<���i2;�=A��B�C�^��<.��<�M��W<jg �6��<aX&;G�h=��R;L"=���; ����4=B��<�2���zC�UN���J<�A<*i�<�E8=AN���C�2��<F�;�?
�qt#<)GJ<ζk�� n=Ā���(H<3=*U�<�8��0�\�_Qܼ����hq��~�;����S!=ju/=<���d�<�ZC=j7�<�+<�*�;-��<<��J��2�&�L��a��2W�����<��#=(.g=���Ϻ=��\�c�<�,
��6!�z�<I�û�t<�`�<�T=L,�<�酼F�<cH�<.V<�p߼/�{=�=������<}�O<#d�<�#;�ͼ�1A��
�;���;��k��]�՜߼���9(����V=��\=~�T�i(��t��<|D=hbW= N����K<)^(=�a=XG��װ�U�<��z=;q����.�-�;.�*=T�*=�XF=�-o<х�<sѫ<U|C=��B=_����?����<�G���L=�/)<(��<=�U�K ;��=��G��ټǉ�<� R<.�<)ō���<=�<�(}=�.�<���<�R<<�����a>=]�=<��$=�aC�� N�!OJ=��<��<��T�>3�&=$��;9���|PB=Y	�è<yt(:��#�`x�<��]�h���}`=��=���<� '=< �������=g��0=Ugʼ�ـ=#2�:��'��o��j�����˚�<煆�Hy���b6=*��T�2=k/�p�ֻ�Q�U
v=�_==}y����;��Լ���:����K�� v<P�ϼ���<��\:�9W=�N$�`�;��r<�̼1S�<��H���0=�M_���n����<~�����=U����ٌ=�E=�O=�.�ld���������Gμ���B<<��ټ���2"��F��=���sl<��ü��x=v�d=m>���^����<-�j<+�=�9)=_E�;���<zp=(��;$��.�<��I���J=�
:��M���L=ﰼ���"����=�����^kl<�0=��:�W:�
��<��ͫ���x#=��:=x=��μv�>=Dl�<喟;��=���<�:�<lo����!���;lY=�Ï<�����\�)�^� ����8)=.q=��=Jg<��Q=!^˼v-�.<=�T&�a�<w˓�l ���W���Y���l�<�GO�lZ[��
%���ؼ�q�<��)<�먼�A��{���{�"�jy��Z��̽��[/��AƻJ�=a<�$=�%O�u�=��;=e�X������ݧ<���|"=[����\��/�p��<ߥ[�j�;�Z><��9��;l�<A$N=t$=�P=r�4��u%��}�<Y��;����x�d�N�;��=kBR�(���\����<E�=k��<�<aC=E�����S��4'=������g<���	��g��</=/�"<}#�<��\�"k%�6PؼҏK=ȉc=0�#��^S=*s������6,<D㉽���<���-Ʈ�(�C=�X
=�cV��
ϼ���<#I����=d��_�9��@F=Uha=����4��<��V��Zм1��<F��y�<��7��<"��]��a��f�a="$=lQ#=�9<�H1=�B!=Jm��P���_<�{<�a��E=6�f<wn=�yG�9��<�� = �<�@��?I;<��Z=�l�8�;�\�a=j��<u��G���j��-5=��~���Z=�u4=ه������J�h;����;��J==�U=�X�}8c��1��dw���>��i�.ϼ@���wλ)��<� �-�r=���<=:0��"<���<e��<ʦZ=�/=�/��^�R	^�ZH�<�]�;����*�"��;<�2<}�=��z�z$=C'<$R=>�x��ō�4J�<4J=s,��a�[<(#=6HQ=��=�?�;�=ʪ⼧�=��h<���<񾑼��2;剎�Vۅ�t��<���Nq�(:)<�!U=g���1;:��<�@̻n�3=#Nf���,�f-/�����0�(�L]=�%���C�5�<~r����;�%�j,=�-��k�^=L^+���X=bDv�ŭk=�uF��Z����x�>�k��$����9;���<[g)=��<�B~��
��r<�rj�	J��B,=�Ia=՟:<RCX=&TH�� S<�R=�_�<y+�<�h6=U��<ȼ�%ʻ�x�=��=��� ���n=�=}��V<�(�x�`�I��<'����H���g�<��\=%��;�ް��4�;A���w�G���D�·�<w��<��:��q�;({�;���;$�Z=�<t��<5����F=��4M:�������G=l���� �K���l=%sq�.f%=:J=,��$k3=���<�+���=K�G=<���!���;�J�\�B�R{5���;f6�}lM��a#=Ё���=0<��&��)��;3�U<[`p�Ѻ ��*�:[wh=g`���޻�Za=�M2<O|�<��g= �r���r<�ׅ�����D�;S�d=j��<���f����H<�y��lA=n�<�;[�=�v;��=���*��<{�M=t���
���#<�uH��� =����*=�-���<��ͼ��ϻ���;I$r�(����.MH=u��<m/,=�K�9W60�}7=߱<>�x<�_�a&=���=Y
c=9a����ɨ��Qrݼ�6���!�� 3=��!=�S=�w<eR=ԇj���I�����P=C? �����;\<V���ռ��Y=�������LNy=�>�;�9�q��������z<�`c<��?��:��<1�Ey��<c�;��t�C���)�<�B�0�ջxu�;��`�sL=����Qܨ�+�-�A���=�b�Ns7�l�_;�F�`��T��!?�x� =��,�,PA<��K=���?g�� @��p�<oΒ;0�4�I�Y��<��L=x���}=�����B��(�<-�|�[==Ixo=��h=o��e
������}��3M2<��[�#��T=]i�~x�<�>�*==�; <:�]<7=��<��k��Q5�CL�<�S�<n�2���<ۅ�<q���&D� |4����������&=Զ=�'�;="�<߆;ߙ9�.i=ם�;�&�<
�(=ײP<<56�:�;G�O=��j�a�	��^��9��)�=6= w'��^d=[ґ���,��8	<-I�[v;�z�0�W=48;l�e=5�c��;.�)��l�<��<����N�^��9S?i=s�S��4=w2=�,� ع��Am�~uk����=T�)��l==&�����Լ�Ƽ��]<_�<=Q\d=ͽd=qz���������R�+�]7<��<gk=uÖ<yS���<��B��_�<2�;�=N��p�O:�B=���=�	ּ��>���9<am�ψ�;��="��r�<��]=�%t<6Y<�&^;��8�E>C�i�>�n�!��WI<Sy��2е�A3��Ȃ<�x0��ь�ԗn�r�"��]�<N�V=�Q��HJ�k��Y ����Z=�sW=��r���*<ށ��ByE�bܺ�kU��i�\:6�t�<�D����=��;��<=�Dl���1={�<�j=%�%�H�����.=�,L=��뼯�e<�<==��Ѽb�<2��=t�=�j�9�<q�"<ل0<�2v�ĥ�]Zм�%�;7��;�o�5� ������:E�'�?���^&<)ɼ���cf�Q�D=�o.��a�<��X��p��2ct:���<E1N�:3=��o����J=��=�a=,���s>����9,�x����:y.��>��<�r%�8����\�;��P��$-�G�,��+=�=s��<�9=�q=��]=7
���8:�U�<��K�)�%��fN�ck�<���`�%;�={�2�6��=�Y��c<n]��(���iü�3�9�#.=/�<y�;jO�<�	=}%=f����j+=����A%g<'>�<�X=�����e�G�������?�V�彼C�N�B:���٥�Z��<Y{:x�9=0밺D׼3lX��������}=ɳ�<�<n I��lj=k�t��%�\TL���7<���w�M=?q��ɿ�*/�<��)=�𝼚v��؜5���A=T�D��?=���ֹm�C�A���f�ZX��I;��c<
c="pS��һE[P��?�e@o<�_�|�D�3[a��=�|0=�$��%��ڼ�*:;�4��<I�m�T�=�,��|�=۱Y���K=_�Q�=!f<�I=���v�<���
�����Q(����R���G�<��7�7��T� ?����^j;]�x=+{.�!	�;¸c<Pġ<�͂<W�=φ��/��<)J��<�Ik�wjk:W��d=<=o��7ڄ�nz���%=?><�?=�X�xo������!.r��,=�;W�RX��:Q=�����d��7b=��'[;�����&�c�<ւҼ_U��J:<���<e�Ph=�*�P�=+�Q=!�=��<��]�z����iYq����%;E=����9=�-=��B={/�9�O=C�<%����=�y��}�M8�th��Ko��٥���<�xr=ky�<C;6�3R=EX=RT�<$�O=\���i=ʙ8=:K��A�צF;���;�D|�!1�<�$Ѽ'�0��G�;�	�\z�� R�;o>|���i��n{��i<�q|=]�A����;MU��/{��`<����į3=c�p��'_�3Ū���B����<k�M=xw)� 7j<�f��@��t�=�Cj�+�@<ޢ]=hV="�ަr��N=J�<I<�-i��̼ܛ�<P�<d�/=�'#���<���<�9�<��=��U�±�<�1,=ͺ�+4�<��<�'ͼ�=���V���#,x�8�K<�Ɠ<�D,��݌;�P�<1kG=�sH<�=��=�JP�����5b=BrM�'�z<����8=G�DD6��.=2�0=��<5�+�qu�;O�.=��.=75<�B��q���[��<�Ԕ�Z�������&��<����*�:�0h����<ޱ-;�M��GkR=�B=��0�m�D�����('��?=��S:GP&�.����D��5�,�� �<i�d�s��<*�6=�#���8�;�X�<̴>���{<	C�m��<�Xӻ��ܼAe	<��E0�&9�;��1=C�<��=�̭߼��}�+��<i�����=^�;��<��=��<�>=1�<�쎻	�9=I�]��T�<�s��s>=2t���sż����b��<�N7���%=>�~=:Nb=�(5=%繼�	=v�<��ռupռ�fV<J�I�����I�<�V<�E>��l�<�:=��=�%�M��:L};@�ü�
���l=|y�=��2=\;+�˼�T��:���z�n��ª�=y�p��X����+< �~�����<�m*�V����=!*�Z=ܘ��M��p�#��(��D�<�=�����<_��IL=��t�nI.=-�=H�=m^%��7
��Pi�q �;�֭<R ;�S
Z= \C�/�Żȱ�;��<�x���<K�#���6�+��;�+B=��?=V\<��<�ּ��<�x<�p�;8;	Ϋ<|f���\��4��w =��;=H)=)�<>�>�s���D켿�M=�C
=#O�]:�C<���-��/:=���:K�)��U<��W=1)u��;��Lb���s��1��5�\=+&C���,=���<s�ۼs�����:�%'��/M����<��Q=Q��=���}�=����OM����<�x�<A�λ�!Q=R`��<�l;1����
���ἪU���s;o�p<��=�~�<����@=4���?d$�*b�5�M;i�'<�2���B=G�ּ��<D{#�j��<���;3aR=���<ձ;=�'Ƽ�s=��Q��%=B� ��9���E� �.=����=Y8�<��&�%$�;��=zށ�;�7�D�<����$;E�q���=Vnf<<k;���ּ
�N�i�]="�;�h=�FL���ּ�)=վw��w=�����6=��=	�<�T׼6���V����k:�(<k�̼��=�T�=��<�E��z�<$�;J<�6<�I;2��hcۼqs�<�߮�
:�)]@=�<u|=7��<�
=[�6�zn�<�i=����<��߼t�J<tO�<�e�4��<P���Rռ#�������F;�v;��=\@�;?�k<�0����<#�/=��==I�=���<4ƻ���<� <ʒ��)H�<@)�� ��@�l���+�4��;�XJ�<|�M=��ټ�7;�� �<b=p���:��8(���F�$=>1@����<�j��A��<ǎ�;��!����8�)��:�ȇX=��s=���<��F���=��e��m��C;�	7<����H�c=�X�I�X����:4݈�p�!��B�1�Q=�	<%s.=�5��TS<�N�<l�L=���<ĴQ�W퍼"
��b��N5�bx�<g�M=��K�گI�8� =���<��W�#</�[�ͳ/=/;=1	�;��v�=Y
<�=�iP��E�;x;�� �TmI<�H�N�Ab=��<C=�0O�wu1���=�= ��;�<Gv���fA=r�=�9`=��`<*��<��m=�cI�����
,<&��<���<�ܬ;==L<^I|���=���;Zټwہ=/��[<�-�K��!E��9��� <	�Y�9�=�ļ��+�ڐ�<�X����<QP
������<�����B=A�D���<i&�<�2=���:Z�;,]�?@c=L@�<��	=bܺ�J�ۺ��ӻLDW�h�㼾��l�S=6q��H�����<	G�<t�����Ol =A�<.t����@=��<��<)��<���r�>B�-����,�K�F�x�#�ߗ =sD����)=�q�$�޻��=~(���������<Pm�<)�9�W��<}m#�<ķ;������=��f��Dj=t/�<ޓ=�d<���!�j�FԜ8�7��2pƼ��4=+��<�9�<(Z�H�c=�=�l;����<*�5��`<^�o;��y�r��z�R�F<N4=��"=���<0/�|g��)���0[u;�9d���f� x?��@L�����ųe;�����<ѓ
����f���_�����'Z6�w9=��<�0+=_r3;��;������f=Oc=s=�;���`�=Z�1<"=��<�JѼ�����<KBD=��:����<��<�=*Z=%2J�3{�<�[���z<��g=���;�-<(�N��v�<T�=!8=�>U<64��{<'6�c�ż"����a*=��ļ��=1_r;�o1�CӪ:��6��P=3L�<�=��)���E����<���*4����<tI�<����uN���%�R��<:᛼�=]CL��u;<Ǡ����u��N�W��c�S� �<��"=m,!�Q�Zd��O��r=}�,=~^ϻ���<�����&<�gD=J���u���E<��X=@��<.G�/��\��<}�*=�'#���<=�a�#�4=�Ӻ�'E;\R��k=g��<�Z�<{O*="\v�ѨJ<�N���D�v��8&��
�,<%bƻ�'=>J�<��o<A9=�g�/����i�<gO0=ن-=�RS� }=%��<���:��<L�<��c�=��;]�J=BkH<x�5=�=��;=ڂ{��<��<=���;*��<vM�<�6���7;=h��<h�
�3[�;��)��k��Hu�&X=Z[ۼ�_w<�hۼ���%��<��'=��<���T���U=�VK=n�K�0����:�)a���0<��<�^= �5<J�|=��[���i=����d��Ӣ�*䱼$(K�^\�0(=��;kp=ƸX=|ؼd��;�8���ټv�D��l���!��Ҥo;�ٳ�Ζ��@8�<�+u�	�Q��h����k�����<����M
#���a��\*�1&���
���j�� =��n�3=B�.==�i�+�j2�<x8�<�=O�B=%I�7
��G"���b����<nD�X�<BȞ���<(Y�VMP=-�������<�,m<`=�DJ��΢;���<M�ܼ'�<Ȓ�;�!�*�[=n=��*����<�ق��j=�1�<�%�<�&,=�ka��W�򏆺{�5��P3�r�伸��<�U���<����@�8�F�=X�O=j˙:��W=�<��K0�<c�;��=��;'�]��XX=XM���/=K���g�Z��!:�\=��;�@=��p<�0���>=m�L���"=¦o����w�%�����7�d=�IT�v�`=P��uQ=;c=�����mu<��~��gz<�R�;����Æf=a��;�w���<��=x0/=��<��x<G��<��><��<�X���6p3=t�	=@f(='H�����4��6�=�eO��ix�<�L�<��0�io=��<]<<�X�S=;�n=jq3=d��R| ��<��O�&=R�J�΢ܼZ�U�/�=�＜,���)�����(H<�S�<=eb;-\=��4<�O=�1=t-��Y�<R@�;�=����,X�;��"��)�����<&r<�� �$�D�6��]B6=Z�U�WZa��u�<�I�;#�M=��>=�۵<����u�ڼ_M=��~ӼT�O�C7�<�N=6d5������S=d^ ��5~<}S+=Ӌr�M�h=�?�<�+��N =�]���s=Т�<��cky=���*����6u<K�a=�(=W�`:Wμɡ0=�;����Q�a�P��GP�3{F=)�#=��=@=������A�==ĺ�<ٷJ�g��~Y����=\�꼍$3�¤�o�}�B9:�����J;���0��<;��5Z=7=W�ͼ*9=|� ;��<(����rX�<�|�<�)d=�w�<�-��򻢼K�=����M=7�;��#���	�!�<�<�=��U�j̋<Z|��.�
�����=݃���= �S��A$O=@�<�8W=�)D�ZX�:ӲG�Jͱ���5=g̯�l���#8h<�=�|!�$%���8f���4��z�{[\����<nP=0�;���<k�Y=VCM=�G�qB�<��=8 =F�0<�+�<��#=���J=Y�={Ư<��<���<� =j\��8��<8Bz��c6=��'��O����<���:�)9=�E�2�D=e��<ys:=�M�ץS=}z�:W+=��=B�%=u�0���=���u=�?:�$y�<���< �S����<)�����<&[���<NM�V�S=ƣ��&��(˼I�U<h�T=wbn�zܼ����8�<�=I�`�=D1�;k��;��
=��`=:��<��F���*=L�T<���<v�ռ���,=L���Tf�? <�>=��=R�Z;�h�
�O=��z��x��K�<����YM�9L���|l=X�=h�v<�\0�XN=9D��º��]��ko=F0%�gPW=��;�p=�c�<	���a�*=y,��)J=���<!� ��><�����f=F� �iW�up�<jE�վ
���b<)I󼮊F���7�	�^�$�ػ�z=mG�<g*A��/�Ql�<��H��ln=4e2=VE�^Q�Vrl�>la���T���;�<a#��=K�<��	��^=)8�;Y�=g����/�<��g�P�<�->�<��%���<��%=t3�xI�<ڒt�o�}=�[<1�<Q₼e=��g=�6G�-?��#t<��f���r<��;�}ļJ=��=?Q��O����<̡,<���R�`�f��D=^y7=��<s�ἇx$=��%���[��1���=���n���Rf��lT= ǀ<��R�@=<��=c���b�G���=�<a!�=	�=X�=L�T=9<�v=s?F����<�?�F�<�o�<}3�0�+<S�<,�{��ϕ;�Η;X��SB=����e��/��o��9<Iq=�~�N��<{i��{�#��3=�c=J�
=�F=u���d�m�&�����"=�p߼J{���9.����9��9��o�<���q��Em�<8Bc�<�������4�j�6 ��J=�h�0q|;9��;�=���sa=��?�F�<3�<�i�;�C�s6<���;�1��a"�(�<��=!6�=�B����G�;a���-=�_�1����M�h�	�����`Pt<�2=����/p�<h̨�'�*��<�<z�(���X=�c���M�d���休�g<R*'�<b���<=���;������&�N����<<�τ�e�<�e��,��0�;=��8��ǼH	�O�+�K��<�=�#^��yk�ʟp���H��}�<�z��a�<�cJ������`J�ADx=U^�����"��?�u�<�˥�� �޼o>�;�� B��L��<�	=;��DGb��=(��u=N<��m<��M���=���˂(���%r��<�=��+=��,�d�1�;��۹�l3<�7�;@,A���a�=��<*�{�=�DA�!Ye;�V=�i)=�~E�8�G��K��=D����=�r㻔Dj�<�=x?%���*=�l���<�(!���2=�0=R'	=��<L�̼l��5��<ﻌ<��W=���%�2=�%;�*���<L7K��᩼��d�[�<�M��k%R=U�>9�=��,=c�:��>K����/=��+�KG:=m��<��𼻦W���<S�"<6@�<�'$=�=G�RD=��tvM;�?X�6�|���<�;x=`�4�4�<��RMu;�t��;u`<��=�'��e!=S.@�e�<�����c���;��ɺ�&�
4��wb<3�E�̌�<�-)=��<*�,<�DD���=x=�8/=��= tG���s��^�;!L�S
�;..
=�J.�x�K=d�.=��=a<��p6=M>$=c���Z�n�čмhh<��ؼr�:R�
��յ;q�ü�N9�p<J��ɼK [=���9�S�N�H<�� ����u�曫< ���Q�c��7���;�[�L�����A���{x��\��&V��@�'^�<L==�F�x��@N=d%^=���<��_<�B��uK˼ و���=����M,<�#C�U��<
����N=IU�|�T=��s=�<�ǂ<�`��W�=�q!��R�;+Q�=c�P��ļN��<����-2$�߷�<�Z#=��I��̼M������T,��8�������ٹ�D�<! <#�I=��ʼ^�D=�=�<)"
=9^�F6b��h;��<a=�����J�v����<��H�_�==�k)= j=MX1����=I�;x�(��5=�;��W=��v����/=5�=C��<�o����)=e7%=.F&=M	�`����`��(<JÐ�G�<�S=��.�}��<< �
=��*=Zi���Am��|	=���<薢<���<�<�n=� J�]kC<��8���::�����U����;��<��`�=����;�e�,V)�׫�<[u�<�#B�|�ɼ>!���m��n��G=a���p�D�A<<���<3:�<l9=<��v��<�.a�� =hI�<�$=��s��I�$�U��U=?H=�Fc;�m����ռ^�9}��N�)<�-N;M���Z<!�;Wx�h\=��:��뉻A�E��5=`��<v��<P�!�=����ü�=|��;�D=�WM�,4=h�g��8�%%���|�<����`�98;;��i=����t�9�0=TC�<�6F=�UռN�;�a�qbƼh�e=������<��R=dW*=nP"<�F=8�R����%=�A��>=0�2��2�#J��
Z=U;�<�g��4��!�|`��x?��  =N=5q=�	�<uIs=ob<
{��g:�b���_B���;� =����2\=u!�;XǼ��S��z���$=���<-�;��@���C=0IC� �=	��<�ݏ<��t=�t;-��;NԤ���"���^�A t=y��;��#=�'g�<�B=�����kv�"��<CNh��=��C��ߘ<�2�;$�	�*�<�}.��
6����<mNŻ�t;��W��5�����l�<�,��
�<*�<�Ļ�<$� ��'=j�u=G"W<H�*=s
 �
�y=�UD���R�c��BM�y\y=\�6���i;` ��Ez�<�=�E��~, =3�;�[߻���<���bk�A�9�!8��!y=64��������l�<*F=mE
�A6�tZ�<1�F=�'U=����s)�<��1���V=#�U=��"�$2=��]=.Dj���1=W@*�;t�<���<"v����4=�Uo�j�n=N�\<���]�<*[�<I!�<k�<�
e;��Q��¼Y�A����s���
�<�J�<�6�K�*=L�:=�i)=ik;4t��C�	=�A�<�$l��Ъ:�]1�2��儽�`�8%���<�b9�1���4��*2���G=��=7�．aټ3�X=��|=�=�T=a�8�&3=D�.<��%=H<=��̻��z���d�Y�;DK�<�!�< �8��#H=]�1��<MNC�����μM2��:�{l�:��L��}����<�<�<@Z��IK�%֙<8�~=p�N	=�7�=�'��!�[��!�;�Bb=Ÿ����C�=��1=���"�<����x��R+e��.�<�=���V=*	=%��;5�=_5(��id�e�b=�"<��<6�V=��;U*h� g���GN�=��&��;�7u=T�)���<�"ünI=A�A=b�O<��¼z�O�Ɔ<������Լ�C3��X<�H=@3�<2�^=���'�}<�η�I�<��V<��</=12@<��j<����?�< �;=Ұ#=�u�<N�<�%��t�d�:9V<�k�����;3:�\3<�=
��f�`�ۮ�<�v.�!f�����E=�~d<��Q�$�h����l�A��A�����<�<���<�a�<�=P>����eq��&[=-r�
�d=���<��=��L�o�ļ�Y�%z`<��T_�<Wb����<#&�	<��Ҽ������(#T=���:���l��Hw�t�_=S?��5�$=7m<=ہ�<��==}n=VIc=2���>��T=fb���D�t�1=`y~=y�0=̊���=9�<tL:�{�	=Ee���Vl=�3켄��<<�)��؂<3�^����_��;���z$^�be=�7�ߢ;�;j!<.<lz�<B�G;0�+���'�
q!��u(��g��nAZ��, ��z�<���<n��;0L1=t�!;��� �<y��_�̲�<0k�=�jμẖ�6�0<η$���?���<<o��R�=t�P=�{�n擼iT��O<N�������C=)�C=��*=ZB=�t���]r<�+g<�1"�3\�<u�ɼ�EH=:G<v�o��(v<q�ܼ��P=��R��t#=�D{��|�<���1&��80=�k`��'=o=�`���1U=��<zVb=_P�<^N*=�>����5��ѓ:�V=�\��Z���XuG�-��g�;�__����<���W��w�������փ�癸:t�q=�3<�ox<�j=�x�<�^�<�R�����<$�D=�	��h"< y��9B=G_�z���\=�qP<�?7=@�ŭ=4��2����<���;�;��U���=n\�<6Q;�І�|�<E�J������J��VTp=�H<Śd<���"����4����<d `�=�G�w|��$&��/Q=��ּ�E=�w=�L`=�/&�Y�L=ʻK��I=��=��y�<�S=�����h=nj�;�=�i^=�� �\�1=f��p���⦼�-8=)�<?���߼��
��HtY<uUD=�Y�<�<���=���<-��z�;= �k<Ҽ%�n�_��8�0`�<	�_�3x�<a�;�<�\���l�)���-.�����x��<���<�DJ='�%=(�%=�X=I�~=��F����Ν;�}= L>=��ﻛ�5=}�$�4J6�fr<W�ۼ�j���U<�&C=8��; zP=�N��gv���;�=r�I�����&�;K;%�=�<�'�;��=�=��;o�!=�4��	@����<�;ü�)��*c"=��7=vNؼ[��C��<���lUa=�KV��U8<'�A=�T���<���,��=(�����;��&�c9=`�<;�[C=ʍG�{�8�"K�<h����.\��a�S ��e-�� ��0ã��H$�r��0}�=��<?�ziH<��<Wap�ACt=�O�< )�݃ <6��ni��	�Hk�����������<�J���P=�8'��VW=�f=�V���<Nݼ��(��|G=#�=�[5�/�<=B\�<�%=c�����<�4�s=���<TH�7h2<�=�N񼦓(�m<ټ:`C��^H�8�X=�+N=W> =m9�W=0�<��M=�ǆ�׊ļ�5D=>>9=���=�7�<(�;D�J;�Y=Eo�<��;�e=��7=/�W=���VY�������B=~�'<�l�ck�_�}��ܣ� ��<��=�L=�E=cXA=s�j<j��=d`h�å�(���������=�� ��5�i�.=���<P|0��F]�|Q��S��o
<�T�<�Ӻ~�伢�$:�d���$d=�sI=;i�YϢ�F��Qe=F6=w��9J����;��M�+�=�� -���L:��ߺ�kC;��:<��<�Z���B���h=Gfw�Z�h��]z=-��=R��� C���d=Sw=2��=���:a"M���e�	���6ju��,=���=��Ӽ�O�����;z�#�J��<�/�fn�H� =��#��W9=[$�<�.�:��m�W=^Jf�v)(=j���8�=� �<i��<x���<��(<�g�<��<��ϻ�)Q=l�D���1=窕<YWO�M2�Ӄ�:#�\;�I���뒂<��W<���1C��B>����+��\V=���-=�	���=�^=�Լ§a��HY=$Z�:�=�_A=�� ��ؼ2B�G?)���=y1�;���;%��J��ڻ�d�<,==y���&=��*�Tʼ!&˼$�+�|�=-rE��Q���j=(�o�x==�T�<����y�D�E���1��<LZ<�=�e��	�<�K=��<m1=�ܻ�������;�1����)�2t���<<ι���Mf�#J�o��;�1�𼴼���5�߼F��;3�ѼK��d^�; �==��/�F׵<[��;��.=N�H;���:H�=f�!�ko�O:]=�9V=� !=�$�<p�=��K�^��?�<I��<��b<�E�S��w�l��>�=�]�w�<�fa<�&Q<��<�WL=6��9��3<4��]�ٺ���:ȴ��q=�q�<�S=�C(=�@=v��=\��)yj�q��;���f=��A�m�h��#@�v��QS��h9�~-=<������L=��R�R����c���0��#7���q=@��R����W= l:�t�<���=m�B=�O��d�<�o�(S<�����0=2�P=�e<w�d=��#�Z�V<��ں����6���V�=,IU=
6�<jr��m�<Du�C�V=(�<=�R<�]�<0Ļ�'�����:��r=3߹�j=ӹ5)7���R�5�d<\W���<���<q����<%�3�P�<�ٱ��2F��Y�;7բ��^=�w2�<�
߼m�c=�7��.=4	ɺ�B;˅=��,=O-=�Żk�2��i��)�:�<���<�9=��7=5��fY=�ؕ��G=5����	μz;��}=�9=��(�y�5<�V���f=G�<@ <}�;�=㌓;��)��%���!=�ռ��g=\Ap=��<��]=+9%=�0O=��<����H[U�5�<�伤,�Ӱ�<X-����$���D��;����a:w�O���qڻ�5�l�=�1����qL<dߋ�V|e=���;ojh�m��;�I��$g�C�d<��6��ˁ��W�;��<ݭ��|Ce���<�Ih�ow<ZQP<�� �B=����������?��;��:0��<�{=z=�C�<G�,��G�ٙ�S	.=���<��p��n<��h=^���@Z5=��=�+2�Z�<�Y˺e�e�!I��/=}��?��+.;�'�<�!=��<���M=�_G�����]=�i˼�]�kכ<��r��OV<1cּ���:�<���0��<g��<��+��*�<��s��&�S�= ���X9/y����%�hh=֑C�M��<U*��n�<�jg=X�(=SR�Q���~9e�R�R�Լ[{;iX�<#��<c|%=Z�=Ժ�<Qi=`]�3\|=#/=�"=�JE��XI�i9<[=���<���r�:�?�B=�I?�Ͻ!����<���d=�P�iΞ;��2�o�<�����<P���c���>=x;=2U���\�y>=Ncм1O=��<Ӝ<�8�a����Y	=��)=kw=�O�L�9���5=l#=�g�;-"���<"qz<mB=!�S=������<�mF�rKU=����Zlڼ���:顃���n=^�=��"=�� ���ͻa=�F=��<&�,=c"=gI�ZsF=%����=�bt=_�:��W�;ZR�<��#=(��<��=y�b����<��<&��<��-��5=E�M�;�d��z�<64�=�z�;T|ؼ���<ޔ'�����x��<NKA<a|����$Q:�<�=� ��B�H'�
(���)=�[-�p��*ԼR����<�����À<:��/��0�KZ���
=�O�<G���D#;�>>���F=�^f=�a�7����nH=��D<c�,=�ы�$�hh�Ze��25μ��F�M'=�;6�=���<�8�cA�c��</Do���q��>л&�<ۭ=�z�44U=�0-=S���;Z<;xü��2�@��;���	V�&ze��KC<�=��w=�r:;�c=�@���@=��q�.	�<T�:�ך,<$w�<�,d;��P���\=�j=A�X�;�\�DkU=�_���P=jA#=�e���������%=���a;=;P� h��&�+=��=FVo��`��ˀ=RK̼��=r)V��6�����<�}�;�Y�5ڼ�0�7<��� �Q���=n�5<]=	�)</@?==��<p��H�W=,2;�g9o:������<^�=ń:��p5=ۚ;q��=��<o��;�^ ��M�g�%;���Jp;WT3<����\��;Y=O=��;��Ʋ:�!kB<2Ǥ<��i��ΏͻH����;a<�=��89����/�=��.=�4����<`9U����<�=��8���;9��=��q�oɞ<�;7>#��?��ټ�jO��)���'�� ��D���RlN����#���=�x��1V=�e=��^=�\�<�{�<*;��9;	�=���g=��C�����v�4w}<r*=,���o:�<��<�� �ʗ-<	��<ː�<	�=/S=�W-�_Dm��@Y=y�~=�[�<�(a�wT=�����J�<c�<Q@c=�ˠ<&�ƺYK"���<(Ѭ<�G;�k�<2�S���A<P]�<�l=ޥ	= �滜�̼�k�o����V<Y�=�F�<_�+�R�;���5�H��
=s)z��H���/�<O��<�[�z�u�G#�-�;�_�<��W;�8�q�%=���[<��Ǽl��S���ܺ�TG]�s]$�n��9M��<�e���<���=8+���F��<�=ؼsR*��B�<����H�CA��b��~�:�s���<�.���j����<�=�S�����'��ZB�PK��H��׻6=\hZ��*�;�<�5�;���<���;�.<[�1=���UU=�<,q���}���:=�<��<��7���t�Xv=����qY�h�S=0k�<Y �;jԼ��8���=���<[��t�W=�N	����<Ug%�XyV=h��1@E�jVW�cV�;Fc=�c=�:���S�<�=�׼�:=���0=<L�L�0=2��;3=q٣��8�<n���<��<�m��"�ۻ�2�/RY=Aj��6�9=��< �L=�\=x�A�K��#�?���;�~�"�n=r�<OX�<QH�<�V�<�A�<��t��F=yzg<��O=��=<\=Iˊ<��=$��\�n<-<��? K<�[=Z!��IX
�K��<]%�<��<N{
=im=$b!����<��M�DCi<D�e�r��=4$��U���_��!�<�g��oC��1߼��~��P���m<�_(<�=����jf���ޒ���C�gT<�+=<d���<�Z<Mb"��;�47=�O�<V@�Qh�<AyO��m-��Q��U����L���=��+������>����<��<0��ӽ��;�<&I����<��U=��v����b�ĺ =_Zq<�a�;��=R���C�;_6Q�+�<�<p)
=���wS=�zi=�Sf=d��<J�+���<�	�,";�[q�(b�S=�,=�Qm��}��TR����/=��t=� �
�<�%�<�E�<�*���bU�����Q	=��t<@� ��+
<�U9=	qh<�����=z�E�������L&���<<��A��Ɇ=o�/�1Z�N���F+=�n���U��~Ǽ�wt=�y��>P[��s��<7cټ��=��R�N=;!ǣ��I�8�����<��}��w�O=~+��_xL���3=�4�:������}�r<Ў��N=*�@�tT?�.Qn=�r)����<���<�gj��j��2I=�F�?I����9\A�h��<�̹n9�<h��`��;:F^=XμXݺ$33<氆�˶9=��E�k��%W��v�<WC��j=$W�M�����"�"��<��<�,=U������Z��4�:�=�ڻ��;<�pV;xܥ��m|:3¼ijw;�Qk�l�g;(ʃ�cN_=�rC;j�Ƽ=;8�J�< ���)=� R�pI=|��%Ϗ� K����N=�N(�-���R�衼������/��q�<�X��ί�ۄG=w]���Sl<���չ׼=�?=p*+�=�<��Z�y-��z=TD=YT���m<�z��N��j=��G�V�>=��]��<R�=�q���4�Q��f�X���=o�]����<�,=W	=��V=R��<�����绤k+��b��<���<M�{<=�;M����l=T1��ң<�Y�!a=A�m�^	l=u��LV=G<������Y�:�-d�N�A=>�=8y�<8���D=<�p�Ok<�&�K���؁�/'%=��UB= 5#�p{����$������=����+GW<o<Ҏ������;Q꼬�޼@l��v���O=�9�<b��[N=�A^��=�=;R�<��7<+l<V�g��;���2�;s>Y���p=��<����`;���-���S��?��ã2=)�/���<2>2�0P=�3=��<��#=V�l�<���<�l<7��&=�&l<}5�C��<f_j�I��<X���<�v���J��5�*l�)^=�&ټ,
o=WR�<�|�<x>=����ļ�&㼍��<��z��m�<�1�ҵ.;m���Lȼ��=Ph=K��;���Ā���,���?;�@���=��7=%CF�o\@=�<R�<�㕼�%�<k����+==ܴ�<��$=x�<��0�g:�π�<��H�pU =�s=�8���=�f����x=�K�<="<;l���<X|0=D,t�C�L=�7D=�e��!��XfA=��u���=��?��J�a�A�S����P��*Z�h�=�m�&8��NQ޼1r�H���m`ؼ{�<��;�<o����=�0���;`��v�:��8;��<'K=M�b@�I��<rL�F-�;ߨ���-/=�N���5���߶�|%H��:�z.�<��/=b:7<OV��ڝ<�=+&�!�;�=X=�=�C�/;kM��6r�:G��<k�'r�<�7O=�%A=~J�:�����+w��R:�Y��@�<ԁR=�!��l���Z�<1'D=dYG<ʼ����N;4?=U3�<6�a���<���9`�s<��	<�;D"�<�c	;=����2�G�N� �<���<����<͠��O��~Ż�p��)�m=��G=N����w�AX,�j���A3(���!=�N=w�G=�==$=OG��>r�.R��
/��&<x�(�ʓ�*<�į,����E�v=i^~��jl<iH=�L=�#ٻX[�xj=!i̼�5>=^
�<��4=���<�l�<�t	�^�s<�&Q��nP<�)@���C=꧅����<�
��$�=�L=�jq��V߼��<\߄���m=�%ȼ�V�����\���K�?�a��(�k��=P!ּ�@Z� �<�e�=�ٛ�D�<'�@�vDh=\�=u��<�˻�{􀼛������<��<�ۼY�><<��� �����[����
;����<F��<�J=6��=��+��w=k�_=}w�<z�����<f|@=Ln�a��<�2=MW�<
?�+�ּ��\=�g=`t%=8:=-\���$=`Sؼ��J��ˁ<�ʇ���;���<��R�k�J��k>�j'h�*��q8�<jf�?=P^=��Ѽʦ ��_=4��<-��e�D=�F=����a�<[<�<e*=1!y;.��<
6n�M��<�R��\�ռ[��:r�-=+.�<�n�<ԕ=.��PE�<*�,=��[���<�M=c�<tY=~B=59żč�;��<�b�<�6��X����I=�`�$��`%��,�8�~-D;T<�����>&=�u���j=�� �jv�;t�==��1=pO=���<{}#��t���2=���<|�&��0�]1���b��.=���<�A�(�-����<��<N���D!=��j�/ ���3=�<O��T�4���<�w� �t�z;=�=٢;��7;�&����<#�m�R�����<߹��"����<�P=4+=͸��:<�<���<�� =M�<-�!=yP�A=��=Y�K�"=.$�<
>���=AH��}T=�E��C����=H"=3��<�Z=�7=���<�x=�]W=�Y��0؇��r�i�����P<�:9�^;��=z�o==X�-A�<���Y���c=�����$=aBi;'�<�/>�W=��C�9=l�<����Xۼ�����K�<q����i=�zJ���#���<��4��q9�ǵ�= ��X�G��i"����#v]�$ 5<�A�
�]�5��<�:{��7<�<�<���7b���p=�+x<���;���<i���7�K9W��~@=�R�gτ;bļ��T=@�<v�<t!=�r6=�_�Z���V���E=Zl�+����/<���Ka�A��<rm��;�p�<I]=hS�<d��<��T��LQ=.aO��	̼V�<�9�<�%��U��Z�<^������Ʉ2��C���<��4='�b=�.�\ K���:���Q=u��A�h<`��������<CvG=�ci=84|�-.=� =�?B��Ko��M��P �O=�@L=3����P��Y�<>" �,LJ�NJ+�y����d:]�߼]�<|\��Y;��<fo"=�\_<'r�J�<���Y��<�X[=�V�<=�ń��w=Tc���ɀ���1=�M=�=���\&�<5m�<�do;�+��/�r�)�<�<�s"=�I��Ż;|�)�+j��R����l_���A=�x=���<% 1=�P��Լ�*у��B �+��>0=�a�<���8�&=� =L��<U��;2<�;޼��3�*xＰ#�9?=�'=��M:�����F�n�<�&,=B�!=�.�<#^=ϡ?=_�=�N�XN-��<(�2=�t�<��m=������JGr�����D�<M����|=�=!O<t$��f�-=obT�{WW����;o�μ��<>)�q��<�=���<��:�+��'6<%7�<���<N	{<*:�H��	}=՟7�}y=ʱ�7���{���`=8O��.�{^ ���5�9B�=ix����q��a=\ej=�~ռ)�/=�����>7��3��`�<=�?8=�~�;=�㼈�<�h�<��=q6
��=��q=F�k=Ń2=	3<�;�<��=����<�&0���#�Sf�<� �Z+=��=I�=��&��}R=wB���(;���<z�:�� �d��<��<�v�<ĽD��q�<���;"�<?2=�
:+e"=LW�1�ۼ�����|��q��6�P�t�'=�O���2N=�yA<W��;@l�����݉�:�sV=w�=�Y`=�f��b����+�j�=)x>=�Y=���<'�a��b(���0�ҽ
����<�<��=N;b;44�<�S���}N="�2=�o<n`��/%��.�;��=�@�Z�}�=���1�;��=��Ǽ�_�ݟ4��Il=Q��<��<\�}�Xσ��P"=X�f��+���弞�==��.+;��<��(=�d�<Hp�A��<K�O�-a �;h��<�<����` <n���yd���cI�'� <�8��5=�HX={�ķ�9����%=IS<�e$<F=���&���[<�Tw��T�&�j<���;��ü�*=s�;�-��.<h堼ȇz<�6�+=T�;��4=[ެ<h �<�ؼ�9=^�#��3 ���z:��E�S=�o��9�=-3��y��<�+=�U�o��<�Oc�h��;��<qT5�b��~�g���i�L��rkr=� G�|�<����<��U<���<�=�<�xzw<-��<��0=L�v=N���n�_=��<U<���}���W=�U<=q5��#�<OK���<�����|L�j*d�^Ƌ�%��<�	���0=�2��E%��� ���t=�_H<T�R��(/=�==�E>�!Xe��bR<!t��#�<���Xx�;�D<E (<�n�/�<2==����[}��xI�<nr�=]�<":�^�o�R����<��<w�̼���=��ڻĈ���1�X�_�Z�x'-=��L;��������4�P�=HTĻJ�<=+p�<β���<�2*=�2F��KT�C��I�'"]=�����Mw<��|�,�]=\WD���#=��U=����(ջ��R�ۯ���?><�Wk���X=��f=:W�<�N��=6�Q�=������kh������C8�����,�(�ϻ�U�;!e=�[�9���=߼�Ci�K5��;WZ<�d8<ʉ[=g�/= Z<,z=��6=+:,���*<,X=���d=���=7�>=-.���Ѽs�.=Z�B�N�6=$�
�MQ!��7,�" =��=s�1��� =w�9=
�7��C��/<c� �U~<���;����K!��r1�>F*��n�����/=��W��_�4��&�� �Z=�7v;O�<�j��	�=7�L=��t�1Jg�v�=��<�J$=I�ɼp> <�4==���<�%=�((=Qؠ<�Ji=o�;N����U<�=.D<�	P=�"g=���;y)�����������\/�;�.1�=:�<#��=Bv�<�����&=��ü\�)�@G��b�<��:��K��i)�����I��p�<�C�<�F_��`��<1���;��W<�6/=��K=io =�R{<6ڋ<��<G!t<>0�{��;P�=�,��,� X����󛿼�"8=z�<V�`�i<g��9#��<Ϗ&�7����<��4��W��⃔< K��SH�ż_�<�jH�hI�^2���=�㝼�df=�}9���}=a��<B��ąӼ��м�]T���C�H��;r#=�+>��j����<Ŏ=�}< $<�k�;�<9��J����=�!�O�#=��M��{��H��<��a=|�=)�'�-l1=��m�0���z�5�4=8p#���м�|�<���<�ӊ�"n�e��<�� =�!��8�?X�;:;>���w�2t���t<܉G�b9�����8�<~X=V�G=�!=�=��^o�va\��0�<E�4:[F=ww ���<P�=oP�Qʥ<��=��@=�?�<��R=X%<�S�3�\=��r=@#);��;��2=�����	�͹�<����]Z�<R�]�����7�<ؖS=Ϣ==��a<��<�b|���C�;��f=w���]�w;j�;��zB���Y�M=R=���.Z��N�<��<�ڽ<{���f�;�X2�Q)u<�T!=O���>C���ZV�p�m�ܻ6w<�7�� �I��&E��� _��<�Aq =��;4r5<&r�<�t<��-=��:<�ھ�8)}<�ʼ��<>u��>y��T��pq�<�(�<\�R<� V�r�����μ�bt���L<a����~C���z<�x=ˡ.=��<�;<������3�<�A��y��<EI�;ݪ�<�,���y=�	2=Mi��E�=�<=l����m�&�F=`Ac����:�G�;&�Ǽu�����S�<_=�RZ��U����"�f<!�I=�����w=����M��c��;�I-<-�1<W�<=�c�^�P��F�D[=|�K����ydX�>�ڻ{k���� =�a=��=}/T���c�Y�;�Y�\��;�Oe=s�<�s=hr�<8v�<V���E� �ۻ���]m�{ƼM6��+���:*�֭��8�U�p>�;{��<�^��X	=a<��4=p1
�?<[~0<�����r;^+�� ;�,���M�<@:{���{��缲q�<�#]�7�ü@��m���@�<����ɼMN�:f$<��%�4;_��;�N��A��<�ּ�);)
�<�PW=��N�"�%=���<�i+<-.�==C>�"
@=u���5�<d�����;0��;����Z^����?D�d=M�F= L���|�](=m�"��V ��j;@��;�V<+�u=#�?=
��_�<��F=>�(�
�3��Y(�֤��|��@;��L=;�=����x4=�L6���k���=�����U$=Q5C=nP�`�<�gʻ[<=�(=jT�a6�<Y�<ƅ�e��;�-9�	�7<|Q=wʃ;3	"=J-6=NQ��	q=텮���*���<<��"�_��<��<Y���oF�<-0��cZ=�./�N�X<���r���^ux<Ho=qMP<��N��-C��d�<\	N<ra^��)����'���L��֓:�dF����;��hg9<��+�+�S���K<��=e-����6=�=�<�\=�^7=�oS���=�L����=��{<Q6"=�	�a=��H����~�^���3�ۚ���˻_7������U�$��Z�l <c�<��f=��2�����^dV=��%�$�)�s�{=�'�s��
��:�	�<��-=�h�;v��;�5�`[�}��;9�*��l)��O��=���qW�=�g��v�C���===��X�X��Ļ(��`�;��l��Z=��=:غ��E�<�<jn$=6G�bGK=j ,���H��[�6���c�����K��=4=�yj=���<\�f=e�+;ɴ�����C��<���h�Q�8Q�<
���n�=���4��<=xl1�(�<w�9<� �����:;'%=�P=�)o��d���_=cU����)�<�ټ� ����H�d�G�݄���3�OAz=^�*=��;?%�tU�<����e�D=-�!=*6��^F��z<�K�<��c�����mP=��<�><���=-?�L����x�Ցy�v�=â<�lk=5�#<R�<B�<��;l =�`��\����Ic%�G	F=�t���<�r<���;��=��;�<��<��<P��<��6<&rǼ�/���:b;P�g�_�Լf'=� ��V��ڐ�<���R
=!�l=��6=�0V=�
;��D=��<�ª<�-�<Q�=��,=�.�<�s#�׺�<�n�<�}<�{X=R���訌���=��k=;0�<�c=)��< ��;���F��xFt=|�;��;ŀM��5��=��+�2i=VQ���[�<�W��W	T=_�;I�m=D����;�Q<�6��]�<��0��^�?ju=a��������d����3=�8U;e�<y��<��5���=3ߞ�ܹ̼b�'=� ��T� ��mǼ��v=�Oy:&E���^��M�DIͼ�r
��m_�1����q|�i80���<��g�����<�=R�,=К�<%�������Y�0=�iȼC�2=jA=��F��O2<�3�<^~��6:�wh���.<r��;X�2�E-=�:=�o�u�=�m�;��s<�,�3:�r��E����9�<�=9=�r< gk=5A�<V~=j��;�Y�a6�<S�=�P�۹��9=�B��bp�^!2�?B�5��<8�C���ؼ?��<�<bl�<�"��k��s�3ٰ<L�Ἡ=ϼ�]8���G�A0=1��<P���~T= *%=��Q�3�޻��,=��/=�W��V=�)��e��w��}��ĮI;�4ѼЏZ�mdd=G�Q�UX=���-:���=�C�K ��wм�ܧ<�=Y.���N�<��#�$L#=^M�<Xs��)�<&��P[�;�nG��<Z��=#�<��`���2�,��߿��8����8� �<������=hX;���O��x�<P�<��ﻼ[==A8=8"���/���*��6��,�:����~ȼb���a�y�Q=R&/�R�0=��O=�L;L'=0�=�)�<���<����� �O�&=�C��o������R�讦���D��j=�ʹ<����d�<�̼�㍻��;���;���`��<��Q=��-<5�<�=<bC��l�GN:��T=�V"�!ڦ�/�;>L1=w70��B�T�@=%�ͻ��v��Aܻ8`=�8��U�}�ȷ+=��=F�C[D=>���fg�5-;=��=�T���L<��=��.<:Q1��  =��μ��U�+�S<i���;1B=l�U=MJC=���̼==xeL���H��i/=BQ��@�;�l�<��<s�[���$��;�e��6��G���M� =��>����=�RS�)�;�<�	�@p��r��<q@<c?���
���<�W��R=����:f=H���
�`=	5c<Cc�Vk��F)�zs3={�<�:��ɼ�h�X�2<\4=�<d����Z'=�N1���<�ؼB,h<�<���}�I=�Ş�n-#�U��<Z�<&he<��0�(v�;�ּx��;�W�;<=�֐�-I
����<�)����<:bU��V�<�O��n�\�|�=Z���6iK=Rw��;|�ټ{��j�����R=���i�I��U����Ч���:���$=��<ON���N��}P=����!=�D=��	=G 4�j*=�J�<{ �,�� �������;�cF������?<O�=W}���Y��<�á<��%=р�Gis��+߼��?�Vm#�̭'�n����J=�<��J�;���ɯ�<YO=[Jk<�
= �9=2v츩�";����n�Xm���9�mD=eͼ��*=_p��c=OV�<���rR�`d	�9*��Z�T(����]
�L�¼ ����J<���j=�G���;=!�U<�*�J�j���-=����D������<�O=�ǰ<���<jc��6e˺��=횗<�.G<�==GZ�<������;�*�TA/=SŻ��=��t<��&���@=UD=�0I����:G��Le]��)�;�Z*�Ȭ%���<,0����6��?;��$=��k=�B׼����u���N�A��<�,
�lL��h�t��<�Q=�5�HCռ\x=a���^"z�BJ����<���N���}�%<N�:��=<<x�j�,�;��L���D������<=�߉<(�����;���<'Mu�F�;ƺJ��2�IN$�[ȼ������&=~�D��4c=�1��gY)���=v>�<�GZ=$�9<�ŉ<��==��
�Ow=��=�y;�e����t���<j�S=�F�ߵ2;6=�1=ٝ2���<���[�׹Q�S<�Ek=a�f=t;=-������<39=���S5�<��<�KN�<����T�<tӝ���0��<�����r����Ɠ��S=�[=��»�f��춼�`n=J�<��<��<���<��><{�<�Me=�N���B�<'HP=
�=���;�ɻ�����z9 =����a�<
Y=h=�����,ѼG�e;.���ּ�x�]��;��Y=�4$�5F�@P%=$<&�Ӌؼ�P&=w�u�O��;��U���<�R,<�C�<OZ=d�T<��0�� <lwa=�����
;��<=�O��>�Q�w=I%P�vA<Om��mB�<w��;��<i�W���<����W��.��'�)=�P���#0����<�%]��P�"���3(;�t���<��w=R�S���?����%@=$�_<�Q=E��	���-=��#=���<���;r;������N��3�<6�,=���H
o<&�,�rY����<,��X=��빾E4;�*=%�M�;�J�H�=�(��z�<$%=g'*=r�e�=���#����΃��i��6��>=�0�`�H=X�:���r��k���żzP8�+��<O�%=�:�Z�9��*=m[��쳻?H�>�� ����ּ�"4�X���W|�� ��YB����:��f��<�Wf=��'j�<fDc<;�<U��<{M��m8����;s#<_��l<���3���8]=��C���9�/�����D���1�x���wڤ�1oC<̱`={�<ThF��t<鏽<�E=O��<>��;C�<�m�ݍI=�h�=�(<9R= J=&i,��zq�ز�<���<�G=�3=_�%���="~»O=� ���p� Ѩ<�l'���}�����=��CF�=�M�r됺TA���Nr<Rhc��f�)�뻳.n<�<f�/=�VQ�c�3�������=��:LJ�6��}[�<�s���J=�<�iA=b�W��(Y=�3�f�-��6B=?o�<�;L�<,=`��(�����6$=RE��q��<&����ɒ�P6��S����{<��=U�:Uj=7Q=�~h=s5;��G;�ˇ<ב��9�8�n�>�<n=(zJ�v.n�[C,<�}E��SD�Q��|��}�<$�W=����޼�qL=w#�<�
;r8��KK��C�<��D���2�7�<��<?��^7>=@�ռ%yB=d�i��;�9CG�쿔�=o�b�'����U��|���<�yn<���<%=sʶ���?=�02=S�V= �<��<�-;�"=���< W8<�V?=�~!������v<h����8�<a?�<�~���^=��F��5,�o07�R�<�!<Jr^=�X'���t������ˉ`����<��<�m�<}=�h�<�\r=��=@�8�>�L t�.ݍ<��p=ø.=K��!UZ=�M����<2廃)<K:�o���=���<�v�U�5�Ř?;]���!׼����ӱ<3,N=	&��ʡ���t=��;=�
����Լ�<!V�;m�<=�4@�v��<]�=2)�;D�|=�>�;�U:v���,��q8�:{�W��g�;��Ȼ+ϒ={=�;QP=��ͻGU�:U#�<a���n���CR�/�<��3=z�,=4�^<���<�cμT�/=����`����v��;�s���oM=76=�6���=��������	=*#��_�;�,=��U=�h�<�tr<ơ�������<@�k�lx����o?�<�z ���=Pk�Ї��P���G<"]�I坻�-�%ng�&	;���^<j��nX<�&&=�ԛ���M=?��;�3�=��8�`X�<��Ƽ�:d��<�u�=�P=e���`s<�?�<.{�;V����N�_yF=�=B�l=L���Z+<q.��?/=\��<`Z<vUM���9��w=�Q.���2��լ<"�ǻa+��4�s���Gۼ��|=�4=�7��k���<6�<9�E=/=L�e��g�Q�<<�gi4=��,�j��!#�{�=�m�=�r��Ҿ���#�>i=�£����:�=�a���l_�N#�<F�=����S&=O�N;�&�<� *=�&�����"=h�<�8=.z���S�'�[��j��S'�K?�-f���څ���<ܩ�=���`=���< y���IM=�=eY`��G=o�=0�3�ǅ���� �ϼ}
=���]Y5����<��=U'�<�<J�-���<̾�<w=��<)�< ּo~<YS�<�n�ND�;�6�<[�X�&r�����;����"<Yk�+E
�Mz*=��s���Q�35��\���2�����k�;i�:4��F;�s���d!��OF:��$=���f�hM�<��H�4y�:>�Y=8��N;�<t<J�p"��=�<4Tͼ�޻2�4=�tN��d$����\v���=.���E<�-<2�T=��!��n�<�G=��<�߼,��=�|������<�.{;-P)�
i;�<�<J�
��:��ڼV[��͑�I6����$�ޖ<�A=������m=��=r�<��M:�B*�r��<ZT�<�4�<�\�<ӳ�<^�<mYt;ee=o�<���*r =Բ�<mA=ʏ-=�`B�KK_����=S�P�=5==F=)|<c�B=��v<"��4�6�e|���!<�n;<,�ϼ��⼈>�<|5��H<�7���[E��S��%����A=�Z	�#~���B3=�9=$�ͻns=XHF=� �<n��V�u:뼌�*=�h=��l=f�'=��O������2�9@���w&=�g�+�����=�E���B^�<%>x;��b��+ӼpC���;%Ȏ��Z2<$.�=��;�t���<=K��3"^=4�<�}j=H�=�����g��hH;�
I�J<��.<��=c=�c=���<fR����b=75�%1��R�3����<�vJ=+{��V�<��4�*��<�u���ƫ��o=W�߼^Uk=�EA;M�!=��;dR<��=A��<�U��m�_��fu���9Aq
=�7;p�]�#�n�fF��k9=�C�b��;�(�䰊��=�K޹�@ �K�r=����]����;�	�<��a<��`�S��<)rH<>`=��<	��6<�".��G�l9=�X=`�Ӽ1&�=	�<6�Y���g�YQ=�r=�����O�<��1=i��;���2g�;�`���OZ=�<2a �q)=�q�<��ջ �;]L��竼�/?���	=�!�<
u�;K"<
sY����<��,=xWB�	�*=AP�<ǵJ�Bt�._:jX	��ԯ�D��-�=!�=<$a3���+=�F7;:׻�����zp<^|�<�9!=^�/<�{)�l�&���;�<��J=V��<��>=�)������M��<�X����:�i3j=/�:�2���4<l����+=�����V=�~@=�wN=O�`=F��a�T�o�
�?�Gɇ=� �dۏ����<C.�<���<=�f�$$1�&��EӼL����ŵ�?Ε;��+="�\=.f�:_����K�󐼮�$��`ʻ�Ȩ<j=j�U����X���Kh��˦<sS&�I
8��)=M�<�1Q=J5=�R�<�;�<���%1?�X��<�8��ڪ�<^�����@��<6:=�K=)̺;Λ :Q5"=���<�o���*<�R=�UI��\����<ѨP�MO<��
�|.�վe�c�<�FJ��=�N�����g��i6��9=F�a=�ټ���&5K���;Vx�a�{�d����91<��F�2'=D�K=��+�8�E=k+�y5<v3=<�|�<�҂��5�<�@=���]]=�����<�:��W=��/<5ۮ<C`I;�v�͂�;�m=�.���nw�m!�<7�t��������p&����<�5e<���;$A=i�J=�h<��+=g�;�%!;bYP��<ZIͻ[�ϺJV�<o��<�D;�y==P�<wy'�ΌJ=�2,=t��M�<�=�I="\k=4����μVl����:�uYC���?=\��yt\�]�K=��:۔�L�b��x;;�c�<���;0�;�Y�8\:�:�)�I�P��hW="�G���m��&k��-f�f~A�yw�<��1���U�>#�D�;���r�`���Y=��Ѽr"R�����=KH�=aͼEXb=f�~���<������I�<MX�<(��<i�� ����x,<a�z<$O|=M^Y���`����;��^��e=�w3�~��	^='q<Q�.<ؐ�w+�9�=��==�WP�׎D��>���5=��I���=��=<��Ti=��)��\��<�>��a�?���:�X�ȱI���P�-�y=<oX��9��!�f��n��jv<!�q�ܼ��`��W\<� ��L�6=�=I���<5U�<�^!���8�UU ��[��!�4��#>=t��;`�x;�b�<�[<������0��v=t�λ�q,=\(ĺ�Z=��d��=����t鹇Z��y������\��t�V
<�'2=��<�(�<�=�Y�;��<��/=gs?�9��k_[=�;��k��"� Ё=v˼�)�~V+�`�<���=z�(��.�<S�,=Z�%�"����2=��,7X<M�A�%����<{p�;�w<0M3�?��;���+e�?G=��=��<���;B��10��
�����n���F=7��<m.<�q�H�@����<�=I�%�<�aټy=����<�ȥ<��@��\�<���B�"�l���s8m��T�<ڶ#�"����s��	:=�_�g��v�<��=�p�7�^p��3b<paE�Ą�<�ٮ�5]9�x�K<q��<����=m�=PMh� O$���f�'� =��A�
=�������uZ<�h���";4��<߸< ����A�;&w�<�Y˼�n���0=��<��<����'v^=��)=�~�<�Nf9 �k�&�ҝ
���;JY�;Z����j �\C<W���Re��)s<H�u��a]<f+w=i�H�bq=�&=�b���O=c��<�K��L	�9ɼs =���K���!=R��B��o�<o],��!=�1�:��u�
&(=K��<��<�v$��Ҽ��������v���
&(�u�<C�g��.�Q��:�� =!�<���_n=43@�vE�<�'z=-���=	���=���<�8J��R��g��,b׼-:1=z��;Wp`<�;.�"�=}����:=ɖ	=�Te��<M�8���=��[;�U
�]>���$d�L�`=(�� a^�����.=�׻� O=MV�q�+=S򔼎*��������
��E=i��<i:��m��*}�b_�XL�A>r;�R*���伬�i�%�&�32��`��^9=B:���/5���d�;R�<��h�}\<� ۼt}��}a���=�x�9���<2�;�'|<1�d�=0=l ;=֭;<���U@A=L��<-��4a�;#0��=<�ю�=w�˻�(S<��>=p:$=P,C�w�L:j=��G�MC���c<�^G=��<�i��U�'���V=�:�<4<j�t�G=k�X�9����q�7Kn���:�J7ؼz�ἰ����.=��v�j8Լ\!
���Z� �7�$��}��a5�kJ�<봈�"6=�O$���C=¦����=���c��y����=ĭO��6�<���<��A={��;qk���ٛ;�(Ի���<��S=�?�<#t�<�qE�[��<k#7=4n��v�M#�ى=��=ݽN=�]V�zJ��U�;&G�<C.�<�9�<oz�<�\;�����a�<�yp=%=Rv=*f��?�T��+�;�=��9j�����|?���j�.\*�<b	�? �D V=�A�����+�#�X^t�r=H"X=�)d:W�=X}+��{�:>��Y=h��=M;<C�\<�Pϻ8�(�i�[=��:=x�~=�W�<C-P:p&='�=]��<��D�*i�<��<��9$����<F�B=Z�J<�d=m/5��r<{ؼ$�<�/=+7޼��<�sY��s����k��|Ի'�i��`=|�=	y6<l܄:?C�m�;�ü�D�h|5�f�h=�d̼70<,��<u(�;l��;�1 =�ռ�==�`�<�?=<(�3���߼�'��	�J�1�.=}�%;F)=�X�<.c
��Y���U=���:�߼aV@=���b�>���-�ϗ=4��K!$=��z;U2�<�SG=ZR'=	��<�����J=6�׼���;��I���:8�g=���<�a�;���<�P,=�&�}@�<2�W�s74��t;	[�<)V�<��<�ɼ�&�kfL=�K��N=gyȺ�&p;�K(���:��6;a(;.)��$YH�S<�GM=��
�q�j<[A=���I�$��t��=e8�r0D=�!<5�V�Xӭ<�1&��7D=��*<.�@=~$��� =�(���:�D��I�´�<U>�x�Q���!=�B�sW�<�q��} ��?�<}�=Lw��6r��H�'Q=y�,��|�<��<��Ǽٞ>=�%t=p�/=��<���=̽<cۿ<m{�;w�h<�a=� �<�6=s��<��<���m�"�F/D�}��<����<cvӼ{��2����¼�:=�H�;���<�Y�_��<=��
=Ql��籼<!A�tQ����5=a�Y�,�.=��d=���<M��<���<���<�< ���k��<��<�co�k=������4Ǡ���= �<]��Pk�<1�q< �~�F�q��g�<�h�:��C<��S��=DI���f=�ɼ�0�LǇ�̽<%_=3���b�;k�=1nX��`E�(����ȺH�<x���<~J�<S�����,��W�<����82=��<N��<_����Y�k[K;�%>=�S�<UP�:'���<��3=\f�<�[����O�A����<�(=8�������;�;~�
<�"�<��a���ؼ�B�<3{Ｉ�<=���=DWf=��i<Y7���'��gJ1<zx"=O <<����Z�ռ�����1����7>�nV�o��=����^�<�B=�U,�H�,�#-�;�D�<��.�Y�&<�5�;���-I=��(��
��2��͔9�3Ƽj厼t=�=�wK=��$=H#�<<�w=�$��[��vN̼��{�c�̼�G6�_E=��<�w�<��s����aI�<�4=i:�;1���n7��5i=YԻ��=
2���a�!�ʼi�
=zC;D>�<��;���<�6=K<5��o=1G�U^�<\�N=�w�<�-�b�Ժr� =q�J��*<<�k9<�Q=P�M�w�==��;���*��[�q�Y�� i=�xW�j�g���6�-�=K�<�������<��!�|t=w����j'< �<+�����\Z�<�"�<�C�8t��x�k�����O6�=.F;>���,��-���S����Iu�<�Z��!�ܼ~[�ѱf=��=�+�<G6����;��;���<�M=�rO�o*�:����ZMe<W o<x�H=��~<�ᐼm��|G6<��=��<=
8� �\=��:<>�=}�m��:O���<؊< �������=�D�����<&R�:�=��,���<X󴻫ϵ�1"�� ��;8��ls=����{�<o�T=�7�TPk=ȧ=Z�<��$�%�����(S�^����-1�@t�J��%_N�7Z=����d{Ҽp�f�l��Ѩ9��#��U<JwE=��K<��\�5=�/<�&=p*W�,�0��{�ftE���=��U=�<bK�<��B=�%�<^Tu���������K�\,��,0:���<��d=��=��-���w�<ŕ�</��<��h��VC=ӫ���F<�弈ח���ټ}�Y�mDd��y6<��.=��84ܺ���[b�ԑH���q=Fw��X$�V�|<�;�x9��[L���#���;��z;��7<_#���^�Z�6��_��ㆼ�����1=�	ӺeQ�<��<1l+��f=�޼�9;�i����:���=FE=e=S�������ȏ'��G3<��X��v&�bԳ�����=U�;>~o=;�;R�<�"�
�<��=ų=��H��u���-�	^H�LLA=x(ּ��0���=��<>f�<H����<-�����5;zF�<�pR��k=zr�=\3=S�%=>O<��R��주�<W�e��%��һ��Z�<�;>�f�\<�F��ˁ�*^�;8�j;L�<a	>=tQX�QS���h=��>�Z�1�鑽��j�W�#=R5Q�����;w�<=��s��=ܺ-�j��<Y���`�<��=`��<h)�Zz<���lU���缌�&=��<f8�<Z�=x]*�@�<���<�W��Nd�����u9�<O =�sR=�NF=m ̼w�l��5���=��=��<�IJ�����ˡ"=��T<��s<�;<����Y� ��	%=5��]�X=>�M��q�s��;M�;p;7=C��;���j�D<�(2���$=B�|=��Y=hv�<=�A���<�uO�0p>�������uھ��`
��a�<ѣ�<z0=9��>��<��,���I=T��#S	��-=LZ=�+��@G$<��f=R�;�ۄ�G�:=���<7w|;�=Uͼf�!='�6�p���#&<���R�K={����
=.�;���<�x��?��:%�'=BC\�z�j=˝���~c���Y<�\*='��<�(ڼ��C�?k<�d��Y�>�(�;��;�<8=�j������r��.;d"j�q����=}�=�lS�yu�<[h=p�z}H=RZ=o�P=�<�1q<��"���V����9�%lL=��8���X��kJ<͞�_ڒ�or�;j��<��\=m*=��~�%;K��<vd���d�=:h�h��<j="~�<����n$ܼ	ȋ;�Q/w�N��<%���,�<iX1����<�@���==��I=&�m<'��<�CJ�҂��Wo��><=� �T�T;U�m=����6=�p =U���F]:6��<+�bI^=AB��,`���̼#�x;8""=D+����dY<DI)�?$�<gr�;¢żS�;<'
���d���x<=���> #�i+���*�����r"�<�#��"�C��=M�a=�Ŋ�Adڻ3!��8<�ʹ;V �<EE<)�<�D3=?��<��=���\
=x�E��&O<��L�Y�%�sz=�U�=O��<�=wz�:A��fP��/п�}��y�k=����U���!꺶�(��P=b4=>�=Ly�<[��<�YM=/���k=|�=l�5=�F*���<�8;�#2Ӽ�<'��z�<rT=��8�l�C���<��<qM���/;�z6�][<�a<���E'@���-/0��_{��p<� <��1����;7�{��p�[ᐽS��~�<���ct�Wh»fn$=���=t|F���<J|W=ab���ѓ;zG=���3�F����<S��=�4ϼ��L���<P�B���E=�tC�¿��,f�C昻K����C=X�b.��o =�M=�9[<�;V=�	Y���<3T]�m��<u��;d���ϼ<ɍ�zZ,�Qip�q��'K�+�S=��Y9U���R�<�X�<c(<�ac=%O`���߼�� ;rμ,B����e��(�h���==T%�6K�<�U��;�(�Q=��r<��<��3��/��<y;I=��=��M�_�%=��ʺ�e�yX��\�cA�k5^�G��<��ʼ���;?��V�Y=�X��_=lE�<Ym1=�1�:W��<�1\;�v�v���F^=�6���=��l��eU��9,=� �<
�n��=�F"��8�D-=�.j�(�4=��:}.�96�<��E= ����1�<�u<�A�mI�<�-�:�F=9tH=-����M��uO7�zE�<�Z%=�+=�튺�<c?�� �A=�:M�ò7=��<H��<�,�X��<��<r���oC��ּ  = ��hQa=]8=�]��ک<^,�i6�2)j���i=X�"�?Y��KEy��Y�D��ļ��/<��<ZA<e�-=�m��\Dd<`7=�d���$�O�=O/=+!J�D=paF�����7�h=
��'�=��<���;�U�;��u��\���4��:�:"y=�+.���=��<��M=i{'<�<R�ؼfA���疋�s|;+$<�B�5=�5�����<��<!=���;ԙӼ)�-�Huz;'�M=��'�u���s��<X;ɼMM���<
D0���S�d�}�t�G<U~x<��K�/�B=k�=m5�C�h�����X
=�R��<�d=5=�)=;>�=��Ӽ�}ȼ��<�f-=]�U=�� =B���6���.^�Inŷuл���W�����:΄�˶P=�k��vM��G�<�$8=^�#�]�)�^�C<���;��_< ��$L�<,�;�`T=��6<�.=��U��P�<n�;�ZȼV�6�a}<��b��;|� ��!=�`=�<��Ҽ�3&�s�8=95P<��Ƽ�$�<��<I	�=#�;c/�)�޼,�T��es=�7��ꌍ��b�{�=��_R<�</�8�=��r<�X=���:_�:=�c����<,�<�9=�m=�<���=�v���=!4i<�ҫ����<��<� 3=�L�=Y�<��<;�<���;���;�������<�|��0;��*�ּyN=!yV<�I��(��<�LT<D@:��`=��<�=Q]h;o�ļuLD��M ��:=*�@=��0�v0=��v�PK=��=��5=)p2=YT7�PM�;nώ������/:=%Dw<��~��3��k3=#Z�hfg�#<׻M��jP=9�)e��BAf�T�<l���>�7=��=5��;����^��<[١�q܅�8�h=��'���Ѽ��� �|<x��<°T=ߒ:�{ǻ� `=k}=8ٳ��M�����<�i�<��l���}����;���<���<{�<u@=�,<�,�\�Ҽ��<�]h<��=n 4� UP�֕���&<����ȣ�<ZI��蘀=�8=���=U_W����a4=�(;}�Ѽz��n߆��5=u�<��+�����g=�k;ք��K�<����Ҁ�<;����uT�{�/=��9�n����z����ƙ?�H�м��<smh�6)=�I5�h%����O�٘�;R۠</�=�%=���<Z�7=jO<C�<ua����z<hv<=���K�ܻ %N�&�<|�
<�-	��PU�H{8=���<�=�<���<1��<��2�*������ �N��᯼�!��Lg�<CbҼs���~nU�E�����<�l�./7<NM0=���H)N=2��ps;ڪZ�dܺ���<��F�D����߶F����Q=8)�<8݌<y�K=�b}<,��)#�<���<n�N=�F��ɜ���=��<*&=�b�:'g�<4�?<��I=�V�R�)=o���=�<UE�<���A�<~��ب�<�]�=2��7=��$�d��<(\��SM����(=O���
3=�L<]�<Exܼ�߼!��<9�K=�<��='���e��Ga�g.켿����=8�c=�W�nZ=��:_c;K�� �;.�X=���j=�Z(=}����<��ӼϤU;��ϼ��߻Xq3��#=s�=��<NF�fˢ;�G�Mk�;n� =F��<�S��D}=�<{rм�:�:)}¼�G=!?=m��</FI=&�<��><#�<9ǡ!=$���&=�ok<R�9��hN���O�i��w�=b��<kt����=�]��K�ߜ�<N*A�DD�=�& =p�<�\@�`�o<PHI�K)�F��B"ȼ�3<%D=h i���
<��Y=G\x��(��8"�����佼,᩼$��g"=�.;;u_��O=2�y���+<�����<&X��8=�t|�<w0<+�K=i}�;�~�<C&���=��/�`�7=�::F���͂6<ׅ򼄭|�����OZ� .=bs/�n\e������]��͂<~4�'"�O���^=�����#=@'�ǻI��n��0e�<'�L:=s+��"�B'���=�K4����mT�Lt=��p�Q�;�8����I	=�3><E�:"i<����V5��(�<N�L���弰k?��L<�4�<g���L0$��=��b���gJ�<���<%=	�������h��s<��~��	�<H�=d�=~B���K=�qH=�$
��]=�{H=��-=��A:�\<4��Y�ؗJ���=��<-�";*v��S�7��oy�,蚼y����<+�E�]lN=jC�=�ڼ��=7k="ݴ:��c���%���:!�2�qbS=�>�;ƚ;�{��X�%��k9�k97=�,=\S�<�఼�0ݼNL;�A�=g=a�̠,=�v�<'�=��m��P����<w���+��<']8=>[�<z�<x
=7!6=.�PI5<�Ȋ<�\3���,��P=(�;�*=.ڑ����<�= ^=�{W=�2E��YG=��S��!��!�:�c�~����N���<;Q�E<�)������ ��TP���<1�s��O���<��ʻl�:��b=��3�4�<R��;мa��܊���P��<^�)���q�2����=߽�$<�<d5����̝�؄|<	7�<v%8�QA�=����으z�V���{S�<��U=��<�I=�<�9�ŸL=�Ϻ<��+=���;�J���$������x=�^�=2g��ua<�-;N�1�ʏ���P=�2B���>=��+����<��<��Y<���J�g<�\X=7)�;w��;/��<x�Z�t!�����-_*;��d<2� �E&�<<= �s׵<Y�8;�+s�O5]=#.A�Ҡ[��������<�8,=G�[��H;ؘ)=WܼL��~���h=���<ʡ�<�_=������?�6����i��@�<O��B=p�����h��1�Щ�;[�r�A�<��]����<WsY=ZӐ�Ԥ���%=�=�9�<|����cE=Ѧ�<�9	�5�N=�C�=��j�ۼ!�����R�[N�<t�<���;r�:<����]-<�-�,L1�W��<�Xϼ��ż�){�Y�q�e<�
�<��N=�<=ל�;��;�6�A=�dH�[YI<�?b=m鲼\�8<��=C��<�['=��1<Tޡ���1�"�; ���,���i��󖼧J��ǌr��i��� =:=�.�w�1qm����<ݕ߼�?=,0�=�Ml� y2=*�H<]��<��ݼ��1<x9����F<��;Z!��D�ߏ���E%=}FJ��=�<q
��F.`��p<"�*=Z�W=i��<fi!<�[<	�)=A俼5~]�A���:�B��Ą=�
�<8�@;
���.r��W��6(��dT�H�"��,=n�+�C�#��X:=�ἼXX&�Pi:;�^;�,=���0�*��L-=�e"��ө�z:==H6�%Sl<t�=�ʐ�g��C�=�x��Ț;�T4E��OI��j�<=�\�`����+��T=�C8=>���������'��<��C��2\�>�<���y��x<�JW8=a`=J�{<t��<~�U�O�M���<����<s�<֟^=C�z=�&=��*<�S=���ۜ���#�<�"�PZ":S;<Zr�<��b;E��<�r��ټ繐<i��=tcO=���,=JX;���Q��ݏ���<��Q���u<��}<��<2��<��<���Ḫ����<�
=mއ��lA�A��<��D=b���;�=u���ȇ;m�h=I=��<<��_��/��v�<H!a=���<M��<@��<���_�͏Q��}t�#�=�-�0�A���Q=(\�;�R:<�p8=PлU�Ƽ��);q�]<�/=n?/�����=��^=/4l=a#s=�]�<hs���{��>2<"�<�ڻ�j��@=uDc�|hk=��j<`���	��O=����<:7=�#�<X�m<�;�Y�=><��Ƽ�\=]�@=�&�0�Z�\�=��=q�w��;Z�B=��ۼr�)=�6����M߅�k�0�2�@=�H��#�k��<N�s=w&�<.Q���<l�=W'=� ���C�&U<V�:��&=z�4=u�"=�:N��Q< 0=���:++�p�<9*�:|�0�+{Q��Q=6?O��L)�k(d=�#���(�3o��Q�[
_�C�.=[�@=p�<<7F��R�<���9�2��;.*ؼc
��"0�눓�%%�ا<נٻ\6=�U=(�B=��:�(=P	���x��,@'=\s#;Bۚ;c�<"�4=��_�*���?�^�8h�<��K��7=b��J����<��w��\���I�<��="Ff<!;K=�0��ݼ�a�4l�<BB�<6�=�؊�|��<�C�&#�<����N�7�ἇi����j=�#�<u?=L�9=��=�ʼ�~����,K=*��rG�j�<1�o<xi�oE=�Ș��q�є����=F�_=�?<W���Yf�-���;'xJ�Ke=���<E�}�<!u
��&����<�Y��<��$Ѽ^ч���6=^����P�7m�<�.H=�_;�$X=6��;��=�(���-��<A�e��o=-S<���=V���s=�5ܼP���E��⚼�q=��<�[=P69�>��<=�;� �<����e=j�m�?7�<=����+�<Q�<ՊI�1���[*=\=����e\=R�����<=W�<�z@�?3_�o(�:�]?=vҹ<��S=åX=L�=��Q��S=��0=���<ݸ�<x���<�����j;i/'��g<�?��`[q=K=]d�<'�6=]�B=M#�6ݔ;72�<-��<U�=b�<�˦�$Ѯ�h2�u_D��=���� =�Ȉ<
��po��0�)��"=<=м﷚<�4ż�f=+�H��I����<���2�ۼ!����;��;�WG=C/�TIL��]"���(�"y =2�L�	Qu9)�����JF���ys=�9=�I=3��<]�=P�<���%�۩o=h�A���=���<?H=S��<��9��H=�`�<��I��-��! ��U�Y���<���'!�<-⁼!Q����=4�=@A1���I�K�@=N�==��$=�\@��s=��O<��¼��<����y~=ɐ�<Z��_���R=A��f\t�������]=<v�;�E=��:a��<Ju�,�����_=m�ͼ��c�i'��A��k#���<m�G�U��=Kd��j�ee�Q�<�  <<g�;�o,<�.9���<]X\=zv�<��}P!=�U<�n�<g4=/3�=T���0�����;N�<�;���$�����o�W���%���=1E/��j�DS,=K����=�.��11P<uk� q&���;�>�<zx<�R���,�<��ڼ���9 =�=I��<2�=ٴ0�jqQ�W!�<��=��̼�1=��e�v�==Onc: d�<�E�;ա�,�_=��F�g�7�>�=.�';@��<ӵ&��|=���<s��H����<���no���T�)X==&<��t<�-ϼ��%=��:z��=	�<�[�<)+	��_�<���9���Z_;�?e= $=K^�<a�=k(<,$t��(4�8T���T=�`
='N��}�<:0���;�/j<��(=Sd=�M|��%=�}������D=��/��h=�]���Ӏ<Ybx=����мDuŻ��=˶C;�jQ�� ���G~��쬼)�\�l)Q�nM<��=�_�;*>�[�:�M�<��:�y�<�?��A;�	�=dfE���1<$Kb<�|����)! ���պ:��;�%�0��<>0켼�ļ��<��<���<�����Yo<?�3<a��<�?A= ����IJ��g=��x�5�`���=	�	<,F������GJ=&$S�1�j���"=� ����<�o
�,��<�E̼S�K=4�}��&�<����'�+;,�'��m�8�R2�f�;�6�I����j� �B��l=43)�E_=8�$��r=@��<�v���>�]����+<j�<W�h=���<"���i'�
�.���D���d��
=맆��L�<��U;BZؼ`	��ov_=���<�� <*kO<�
�R�1=/�W�����<�D`<�5=�`K=�m$=M9)�� ��=�#|C<:&�<,�[�+=�=`�żz�a=@�<��S<�� :���<6�6�\��<�_Z�˘<�|K=d��&��;��N=I��<�������<� h=��̼'�p<2}u��v=�$�)��IT;�^.���@;�cL=��<=���<�l%=h�?��b
�VfT�ɾ=�<Ҽf�<��<�-��?���Ǽ���<m�|=Y=�l;{q;=��"�@����,�==�}T=�����<O�5��ɢ;�� <�m<�%��yU;�W%�3�(�ݸM����<".6=$�
�4tR=A�=�,�;L�=p:�H=ʋ�;N=���<v��f�M���=��Ի��?���;�qb=ў�<�6T�g��<��4��eb<�G�=5��<M�>=*R���"�����=f����<���}c;<���?�<�U�<�4ӻ�S�<t^�<�?=��߼ft)<�;f��<�
=u�*=���)/=�=�С��	�f&<��8=#UO=`��=�Q5=�M��71<\w �Ei==W�L=��k9~=�k&=�Z=WVd�\�><�aV=�rz="B8���<�����=�
P<��>�E� u�Է���Ɓ��D��HM=�>��w&q=�HX�(�=]b!�ס�;�;V<��z<�a��^���������<=H�<b��<�DD=���齆=؈��0:��X=�^���E=��0=��<f�R�K<X��C��� \��<�P�`��;��{�o�=}��<S�?<��9=��b������24�-Lv<k�=ޘ?��_9��/�;��<3}�%���;�y�;�S˺uV��h�Ճ��Ƚ:�09C<�mX;��Q=���<U��<��{��t�y�;<Q=��.=<H���t=ċ1���<����N
��/&��<��
`�</u;�9a��ޤ<7@<��'<Z�<��<a�߼Sn��ߌK=���<Y�j:6�4=��=���<�f]<I��<-���&�'Lp�]`=W٧<�fy=�=/��<��2�j��<��Y�M�9����m =K=��"�0@����<��K���=�"��A�i�r=g�<
q]=�0��:��<����ǚ1������8==u<���<�N=E୼��D��Rʼ٨�<���qB<K�=ۭw�֗<̢C��A!�z��ʢ?��;!��<��K�d=��'<�����4L�ĉ�a�
=�����Nͼ��7�w��<�6=���<�xͼɪ�����R=�j���=v����g�l��F�:o^�:�Y�=^4���A�o�a��F����<o������7S�.t�nD;=s`�<̻�vZR��H0��+=�N�i�N��cg�,x=�{���g,����:J��X~
=�-1�g��UT�<UD7;�[=�	ۻ�f`�U��"�R=R¼s)5��/��ٷ�;)��;
�ܼ��/�T��#���ZI"�E� :{o�b���G�^=툽��]����lk�<�<J� �M�8=7�j���*��ן���*�p�)��"@=ג <p��\�ػ:�4<b]˼���;����Lk����2�%�AB	�C�J=�T�Ŋ��"=�=E�I=yB=)Kr�����6�/j4=�%=��=G�B�Ih0�E�P���M��H�;��|;�QJ=���o�Q;�@[��<�GJC��(=��I��']=1�[�u*��F�<�k:�x��;y<�8T���[<�7)����<�ы�J�J�S�\=���<�4t<@�<,��;� ����壂���k�"�4���=0�4<�<M=�j��D�<]��<�`�<�8�<~�,�(��!�ỉ9=W��<��'=4�缨�B����<*�Y�=�X=G
S=V�<�9�xn�-�:=X�<=\��S�k<L:�<2�༔ٛ<R%G=�ͭ�\��<CT$��#=�7�<_�ļ�<��<�$c=�y�08W=z�<?R��U�=u�绵�i<!aϼh�<4��<G���ջ��
=�ِ<���<J=��L=����&A��|=�n�<.�<�[�獩<'�\�Cn2<@�]<�O�;ݘx=7&d<E?���g=H�i�{�x=˗`� �����<��=`��:s���Г�<�
<�蔼4=�U<�B���ɼMܼ�[�~��JB�6W�<U�=Z@=����2��G���W�<�K�;A�޼�?���<��#=��6�4�.=u#=�Q)�U��K��׫<\���v��C�S�0h���= �j�.�<m��-8=�pC=��,�̿k�S�v����=��5=Op�<�"Ƽ(���Ō<-�|��T�����<������;��\=u�S<�#;�.p<�-=��<�ݼ_�L���ռ�ʀ�o?���b�gff=p��<�
<L�<��<�3z=�����4!�<x�<0l)=�����?=h�+<��=�K<[G��F�S<��B;_�׼.��h;������ñ<���<�86��@J�����-<w=��=�������Y�;����H;�1<�"=)�Q�ʒ!���p<�R=�������̥��s��ѳ|����7�
�L=� ��\�� ���<�ɼʣ8=G<D�/�Et��,h$=E(W<��;>1��窻+=Z,W=�;�<^tn�CQ�<�)5=�'�%�E��W<�ˑ��pa�*܎�d==��:$NƼ�k#<�l;��=��w<G�<P5o<��)���<�Т�'�J=Xa=�}=��"<�O�����U�M=�&$=��W=��f��tm=�}���J#�Q��<Z;�"�;���<�%�<PP9L�]���*=�	��~J�WC���=����@=] /�φ4���<�V������ ��h�*=V�<�x��s<�<�[�<��r<�jM=ѳ��=���l���|_=�I=�w�<Ĭ#�� �9�:�<F�g=]����g��J�x���=):�4�м`<�G =�<0�D<���<4j�;� =��=�\�����_:���=ӝ��u=���;�+r��K�����<��<��T=� 	=I<=��hh�<8�1���F��1=�?ɼ$�"9Y��<KI=��K=r}="Y,=�3�<�<����<��:Y�<��+=������]M<�/�[�h��;��� �<X}<��y�G.��-�/<?)=�]��Mݨ<{]ٺ΋}�o��H�<�Ӡ<��
=��%�� ���<=ի>=�����7� �S�Dr�<�Yw=�{<�}����߼�tN�-g=H�3=�w�d=�=v�$=�:=4^��MY�R��<��3=P�=��4=3L�F-=����h<=y���`)=�m=��<��5=��+��7�FIX=��=�Mu=}�v<8ȼ�z�<��N�r��;e�,=��=��ɼT�	������
�eCN=�c<_�0���)�.$��-��T�;�y��43��/x2<�3.��h���fȻ�b]<���<���� X���&����<��W;�𬼀ɟ:�l9���6=�V�;6��<�t
��轼��T����5�<Vg���l���$=��[�I=2���Ҽ�L����b��'��#-=���2�5=k=�^B��[:=A�켇�q�./=�}=�g6��������,����#=��;��y<��=��Q�|�D��=�����k�=ضP=h˄<�=��;;.g=_����j<�m�<%�7<�5�<+=*��<1==_�;�/	=�b���˼�`�<RDO��8=���:Z1����e�7����ʔ�qR�:�O��๼�[�;*_;+	=d���pE ��?=�	��{=)��<G��<�옼f���"�<�:z�p�$�F���j�I��=m����m=	�=�#��8���Co���#�)-@�XEI<�>����<V���=ۦ9;�t;��L=-l����g=*�=D�B=	�5�p����3d:T� �����Md��2���K=i7�
�=�V�<����fN=��0�D�l�X�?�T��f����3<�ay�P^�;�m��k��7��D���v�<��g�Yg�`�<�Y�:2'<�6���<gR�t�S=��h=��ٺ��<ѥ׼6�[�[��;1S���2=�����?=��5<]��<<��9L��<Kg�[�X=�/=c'	�kp���B�<��6=�n&=��<��B=��<�'��w�R7=?u5<̇=E�P<O��Tn��(+���<�m1<s��;k�E=��h#_�B1=�&�����<�s+��9<=��5�+ü�kӻ�U=+RK=�G����e����:j�K��k��z���=��A���
��f=l�%������
^�<5=U�=�ϼHm= 9=�.�X$j��c��v�;�`�<�`Ի���H�<G=�v����;�������>�G*�u0�U��񹼻���~p�?�c<��.=�^c=�/q=l�:w�$������5��;��<dk�^q4�L7;�}=��0=]��;�'�;#�=�K��v�9�ZM=2�`��|\�7A�<9k����!�nർ��P꼴�D=�3-��i;󼶠c=�aQ����<��d:��
=�D��&�C����������s�=�ĭ<�<��t=5瓼�� �`Cw�'d
�8 < ����=E}|=.�u=��`=�=EV��:��<��Ļ�t}<,��;#Yi���<��<��]:�(��Y=f������=g+�;#j= �`<NrѼ�\<A�y=����!P��F�:�3�<�~���#�W�`���~=�=�*=&=\���N��9J=��=e�5=<��<K���S-�"ۭ�� �;� ��s�;�_
�1t[=��#�h�ռ���:��i��3=�W��>�W=��<�*g=%�*�7_滟1��5?��P���*Ǡ�b6��sk<���<���<$����w�<v%��m���:�_7I=���v�λ��D��o=�R꼥7 �Y�<I�.�	�#;)�==f\��0P�<�<�;��!��g-=���<g��<���V�|;��<�᩼����5&=C���m�<���C��R8��c���<�8S<n`!����4Ku�c<5���.�;�[P��]7=��*=T�b��<�?=v}��>�a��[=c�ټD����@�(��������<L�=�Wt�2D<�Ge���`7���޻`�����<y,= Ӽ���=�;=8
]���<9�y=X=.=���������i�<}�4�V<�mU=Ő�����R<
Po=�޺^f5���	=��ü��<,{��W2<�<"1=?킽/��Nz)=�8<؜.=�r3��C�<j�Y���<"�<}��<�<<��<i���r�(���1�C=��47��1��Wc�-:=>�;�	��}=�`4�#D��ì��#N�v���i��obҼ�+�<���(	��5����_��v#���=�P��4=3�v=�]q��N�;��<��{=)Ƈ<�#7�9�F��j������c,�������<j�U=\��<e(������<Dd������x��-
�-�M���X���Z�Jn���<����ɯ<��J=�ͻ1�\Q<	�
=o�=��g���3=��w���=O3='�ҼZ~��'��t҄=V�7=7Mi<�G���������9=��J��=��e<�m�=_��<8*=�T�N��(��<Y�����:��<1BW<SS���?^�Ͼ%�a�m��%�<A&�����;LOQ=]�t<0z�<M��:�>���	=��=�i���ʹ�B�!��k>=��*=+���s=�>=�C=��a=�Yt� u�yg=��_9/��<���}:��`&=�˛<iU�:�;=
U%���I<��U=��`;yF߻z�=S�<�M�~�#��cK�B��*wd�dK�����<VS.�"�;�C��*=�Na=�-=I<��3=�N&<R�<ϭ�<۔�<fs�<����S@�Ή�<����<>��<�<m(=O6��Y�ŀy=��L=���l<�<4���j���W"�2�=�W�!.����;�p;���J�U������<k?�<
�K=pv=\%�;}��=S8=������<�.)=Vz���r� 2�{k�<�޼A`�<�=6�	�>+�g�x=ׯ���s)���< ����	=�<�.�<����,�Y���}�ŊI��	�	=&���u���Qм.$�=K#� ;S����|:=3ʻ.��<p���9@��9�;z�'=��`=��6��&a=]s��إ=[{=i�>=������<�耽�5 �D�b:>h!=z0-�p2[=��=�ڧ��m�Y��<4�����4�¸��I	=܋�<[I�<6&L��dd=����x`�j<�t�%�>�6�q=>;�?=\-�<���8��<\0�1��<��!���.=5��}ļ��`��4���N�<��<R�<%�<B.F�'���/=�H�<�*=�����8���#�ؼ0���<=�I=�^-=�KQ=+���a�<<��<a��^�ռ�N'���`=��=�=k"=2f;o�;�6�<��=pؐ��xN=n�]�p軷�Ϻ7#�p��&=vĠ<Le �[e�`�ȼ��S=�+E��g�%7��$���!=S:S�1�U���=%��O�Ἰ>��Ic�J�=xqu��3 ��mL��P���1l�VP���<�� �����S�� b<�S=}�8=q �����8��L�u�=�AL=��<<�d=�u�<Z�"��}���M'=�}�:&;�/ϼ�}�<��8=�3�<Ő��%C=[�s��mT=b�v=N]�;��]<^0=E���M�:�	.�I������<�۲;�S�<��$���<2@�n��<��<�4��f+�=����*=�t̼�6�<���<��ּ���������^=p�6;��5=�e6=�#�M_=-&z=H�<w�?��#��la=��=ɝ����s;�
����H�<�֮�.�|;m�/�bp"=�nK��< �Ԣ&=6�<c�+�==÷[�=c�=�U�;NIg<"kѼ;�<i�<��P=��g=4�V<�=��>=��<��<��Ը� �<M�=쫼��W����<=h<��T<3K�&�<��X=�BA<�黼�@�:M=*�����B�.=�;<e���E<JY����<�u
=�_=��f=0zz��+�"��;��<�m�=z�=��o=B9=����FM�<�.;�f<ʯ�<��=N�1;\���1_��=���<��E���T�믰<=^;���;��r��(=D�L=�����Ӽ�����
�ֹX�"I��2a=�@�Lj��t�8=�>z����:VU�<�Q^=��4�1 �<�1=�5='�<fl*��C"=͛A=�k��S�B��鬻d���(�<���i�<`B7�\=?�<�b<e/)=�1��.�;�yy=���<m\�<i�ɼm��'ۺ��H=}8;(X=�}м�vx�m���79=N��<gDӺdVڼ(n��~����X��h=�M"=-6m�����Ǽl��;�C���P�����ʝ~���<���<1Ⱥ�G����<E�Z�d
=�ۻ�jQ;
�伄U=�E)��J;�L�=���<����:��=�$=�0̼�E=ڀD���=-�&�Zӏ�S-<Q��}@8�񒼾�&=�)��
�C�;G,^���;PX�rC4=)��;Zd�<|�M�1��<f.���8�0������<3�<��{�شm��f,=�a"�9=�=�򭻽`�<�R׼�S<�o�<ƈ��(�<D[)=�&�<X�輟'G=&����G�<̏<���<��<N*��3E=>��<d�����P='l�9��5=�&ἕd�s��� �D�C]��1�=! ��6x=�4=y��<�=���9�,��ڼ�)����� ��JF�<i��}I�:&
=_��u�:t��<���;�;D�;�Nټ�v@��w��YO/��u��A��-�o;F�ּt^�<��w;$�g���>��<V����V=��ؼ�'�=�|��F��<���<��ۼ���!������\�v=��w�B�t��w_�\�Լ�7=2K?=�aM<�:<������G�<hT`��0��.T=>7޻��'�7;�=G��<DL�<?�0=5"��V��=�:L=TO<��F���������<} <�"&=C�=H��<D�<�dJB<�b=�3���s�c5��Nf���3����i<��X<Y���r~�<[�/���)���(�3Gj�ԑ�<:Q5�"�h�(<M=���ׯ3� �s�w��=]x��s��6��J�����<~�<�D=��=�U=�+�:�<�D;�?r��	�1d=#�V=�E[�Y�3=w�=a�p=y:�~ ��6��=#3�<Ғ<
�<�k���T=�49ջ� �<�f�<��<yOn����<l��;�r�_�<�=VkQ�Kͻs�<��=�3@�`=�<sMd=
�;�e�<C�
=[�漧={l�=2�r=�"�U��8�=W�<�\<�N<��Ѻ,���b5��Cѻ:�=X�:��mp<.�6���k�c=/�[�R�ͼ�"=��<Hl4=-=4(�<�h��{�<E5���˛����\t�;��=:;�<��"���b=�r�<1Y=rd^��b3=X4��lh<),<��={�5;�0I=�f���=y
����Ի~^��{?��މ��[|����9G��Gº��"�����<_3#=R|�;-?a=���<���A��<ܔ�;?kH���n=|;������<���?9`<i�=^��^{��:����������;��T0=Sl< =�*<a��<W/��A��<�*���4�<q�&�,�{<�{�<�����Q�W����t=Θe�
��k�<$F=A驻@e=���<<~�<�Z�����<-@���O�-!�<=�3="'L�͑��2=�n4=��u;j������1�<�n=��<����/K�i�.��'!��V��wk=��E=h��������D;�H+��s$<�c^�H�Y�u�Żf�<���@/Y�@��	��;���讼܊��q�<�~=
X=q!�=��}��NQ=����e&=�A�;���9=r(�9q�O!<�=qk�~�,=HO=ِ��o�^�r i��&=#����/߻��ټ����p��T���g����J$���ּZ�>���W<ܕ���0=˝g�e,b��� =,�J=�����8�.=(=��9��63���G=c,=sN+=k�Ǽ"3t=�=N���< _ =�d=�U��*nx����:��^=��=Yٍ<r�$���-�����|����$����:p���=��<	{>=�Q��0�A��Mk<�G�*=�<'��=��<��<��{=Tq�<0�<��k=�l ��L����;�0b=�N����S�\;w���^�;�䰼�>�=<i7�a�^��H*=m�_;4��2��*�<~
�
�&=�dм���<�il��<n�)����<����=9*�&�<m�=0��<��C=x��<Yv�MT=�n��i-<Y�B���;=ю�1�D=u�"�)�#=y�<�W=�D.=Jl�;&���n\�m�-=�添b״���Y���n��8FS<Hڦ<�=Y�ZH���QI��5i;�u��f��xM�&Qb��-;�R=����P�!=�->��O��w7�wݼf�M��ڵ<��(��gq=6�?�����t&�^��<ҳ�[!B��G#��se��z�<Ӌ��\�����Ѝ�C�j��Q=�eV=�+=7� ��(.=`��`�=X3Z<gu4=�\��I<Ϻu~����<�_D=b~N���?=ʱm����<�����h'<N�E�&�X� �K�sY�,���� �1_�<�" =�>���o=�o���K�<ݤ=���O;��G<ʯ �y����/=-��<��3�גͼ	=H�'�FT,=	t��j^���(��A{<��Q=9{�<r߻<>��:��ͺ7�<s�;�g��j��<��-���F�@��=?�=|Q�<��;��A�G��OH�X=R�d���������<s��;�s	��6=�^=0�2=���s�L��:TY<�h=?�=�_�<���:����I�)�b�X�v�=��'=�=���<�� =�v=%̵<͚��N=c&�;3ڞ�+��;~��<f=�$<�J����\<��<��5�'��<�Rw<Zi=�:x=��˼���< �{����)6�=n�8�_�<�+;��<|�t�HT=�\ϼ	�^���Z�����
M���I=Q�
�o�s��ȟ<�����E=�R=_�%���<p�#=X�6=ੁ�o�ʼ�uI��Ʊ�5("����<��<�(N=ۆR�aL=1�9=�==��
�W�m=�=�<WDX=�=��6:qr=p�[=^ɟ��%��{$9��<�Ǝ����<�=�<���<��B=Ie<'���<�Y��)���]y<%=��P[�8�Z�ځ{��2=�L�<��R�����eh��#[=�$�����;��;_�=�u����=~J�;q?�;�H;Z���U}=f���F��Z���<�Ǽ����`m����c���A�˼y=���;8�<��F=��l��*;��g�l�<���h�);Q���Ua���;�V;4���
��ջ��n��@T=��1=��k=�Ġ<4o�<��j<���+77<,�}��;�p(=�Fs=�z�;K-�����<�2ؼ6�_�h���X�<��;Jk�<ʜ<=� ۺ�!�;x�=nnx:T�J=d��9?�?�F#��?k=zi��GM��(/=jｼ6G:=Cx���`=�-��;����B?=�M5�����!<���<o��<�/��>*=":@<��H=}�q�[��<�<失�jkx=E5L=��/=�% ����<��+��}<�&/=<4D�Jڤ�@�)���<6����D���O=>Fv=�:=��p�����hK��7=�ei=9���c�;p�U����<�o6=U�{�����	Ƽz�"<1c��(�_���OE���<UQ�<���{�<�C=�O���6>=���4�O��T/<�r�<�&Y=9�E�\=�G<��[�I��<��i<�r�;#�K��Z=�qO���r�VY�����
=dI[<�8����O=Chb=n�J�b<;�Ƽ��Ҽ�7��8��<��ټ�T��d�<x|ʼy	-=^H8=gn,:$*�!;�:_ߪ<E�V��+��q��:ݰ�<���<8F�=�r��'w��g�{��=���;������O��"�<�W1=���aV�p�f<�Vj��ݢ<�����<��<��L��¼Wxb��N���;4�׼x�(��̗�&�u=��3=��Y=��Ի��F=,�i�΀��N���|=2�J�=��<0�+�5���,���s[=��<�F��<���7�;/k�<g�F��Nd=A	��'�<�W�<�/�;?Gw�Fy�<�s�<��l=u�P��+=�8��㧼OeS=3&λ�i#;s�������9=&����85=兞<���<�,���j!�ȝ=�y!=:�A���պ��)�*P�����@�=�N��{�k��<���<��d��ü;�%=���;EI=v�-<�;�?=�=><�)h�W����)��Z��W�x�L^����D=����S��;�m����A��$S��#�<�m���`�<�#�O�_<|���W�=�Q����Z�@�=�fZ=i�<���:�Q;�.���˺Eu=��f�m�����<��&������G��=l=��l�V�?���S�s�8�KK|:�>=����Q����t����<ub������|�˼ڜ<=$w\=vA�<�q=:��<�P�;d��<�8~�k5=�2L��W;��ϼ��»,�Q=�Ӂ�]�z=S�O=�m��r=��a����<����ӻ#I�⻼ɐ"����;�%/=��{<@�w=g<�+��ˍ��59=�=�T=�H�8+FA=�滼{- =F6�<� ��bt=��8�z<
e<��;�=���<A��X�B:��
���2�����-�<�=@pI=]�b���ɼ�9&=��=wp
�+�;��ռ��1<R^����H=QEC=@��l`��贼Tۻ�>=� y=A
����ں̯<4�$=��=�)�<�<�Q�c{����*SO�q�[ӆ9�U:=�j8=?�o�h3=��P���\;",k��fL�P�-.=���<������P<F�Լ,�#=���<����X�l��c�<31R=�7=d��nB=�?�<U�<��b9�¤%=	1����޼��N�&g"��`�<������<&�=3���?<C��,/ <�R�(=��@���n��{����1	�0�= 
��C,��ۧ�����<A漃���i@=_9�.��<�2f��\=�܈<��=����ś=�l =`�����:�P�"d��
C5=]�%=�fG=�U=4#?��c8=W<�v�$=��1��3������3,=��{�i�=�F=�˖�{�G�����nb=��E�0F#=q^�<����"o�����a#=h�A=!~w���==(|�L~��S��<Q,�<�wr=*z�<uP=JT�6R;�p<A�i<�s�<@��_�:���;Иj;~h���l����-=���<�����\�g�;v��:�D=��<��;W��;[V�<HA#�_� ��L�!]�<�t�<��k�hm�q�Լ�+����;F�����=�F�j�Ҽ�D��O0I=�-5��>]�{��'� ���=����]Z�Y����A=W
���
P�$��N�s��������R�b�z�w�� ��#�5���v#f=V:6=,�^<��x<0���w-=�
&=#=�L=8�<�4�������Y�מA;��=9�F���r�>��߼�ռYD?=)S��'=��x��0=���<�`�;1�1�U�+;~>�q��</�(;U(h�S��<n\Ѽ,�a<<e<�9�=�����C=�[����<Ol7=����,=���<�+һlI��j��U>]���"��� =�w���Q�M=+=�t�<KU0=�U=��< ~a��,=/d�=�;�<u*i=x��V<���;�K:�Ϋ	�qh=�K	��U���<9k��=�=��Z���Z���ɻ�u>=��]�}�<nZ.�Y=�<��3=������;��v��1h=#�k��yȻG^d����<lU=gra=��j=��.=�|��61<t9��&O=�k�<�X��È�G�F��.=}i����<��=�N=D���� �<u�=�ٻ<D ����7;��=�Q�;y�缒�Ƽ�d: ('=�#���q�eռ7&�u��R���y�����<��c��p�;~�=���;��=��=K�_�����|<�<=$=��=|�<�H�1u>�}��l���5��O��-`��=��E����s��;V}ɼ8�S��=�=�$@=<�9<���9q��w:]=�Xe�SM=��ؗ&�dw=A:�QJ</%v��i�a)�<I��;�	B�O�ۼ��G��X�C<x˙�έ�<HZ=������j��(<Bz�<�Bj�;�<�����0=��<�#H =���<�@��0=R�ϼ����/A<)�l=��ݼy�=4�׼��=>#�<b�	=�[C��#�=��0=�M$=�[�<.�v=oj��	��϶5<@Lh����8�N�;H�\[=���<#�+=��;;�V�=]ݼ O=�@��=��F�[=bh]�noV=�\L���G=��+="��<�����A���;�Г���Q��r�<Dyr;'O��Iv��_����~<�EP� H�������:w�������<�΅��l���ż��i=�X�<�RL=W"J=�}�i.6=QL@�hJƼJ���
��0
����D=]�c;�P�|�x<��s��.Y��� <�v��B��%ºS��z�����<z��r�1<��/����<M1�<'����G��['� n�
�=�,�W�=�Ǻ<Ѽ��|���r<��2[�<C:ռd+��7,&�A�ڻ��=���=x2��C	�<�4��ހ����96�<� ?=�0����;l$�5��ǆp�<g=0�2==��<%T=U9�<�(	���]�E��<R�����ٻ\�=� ����;�|�<,���K=��.=�9�<{��&.O��ǻjח<��9=~���&=z�#<�3мPX��V���ĺ��3���6�m��{����ù���<���=�7�&�.���� �ܣn=0|>�Yk�<�<O�o����<]�l=�4���:�w��<ӼG�:鲼�̼?<<������żY�<G�l���<�����<d89<��=J[�<<;���<�P7=��<8���6����s�Hc=�W<� �;�="WԼ�A�𽄽S�f<�FV�d�.�NG��r�=sv�<8S��P�=�&Ụ{<�4s�ې��|�/����%����k��+d='<�:�;w�~<�����7���>�J��<�h���<&()=����ˆ<����fR�<t�'M\=��G<U<�;ȓ<7l������J<�yP=.�=�V���*��h=�0-�����b%=/#=TPϺ�g(=��E; Ò<�������<�Y�<<b�vm�<О���yܼ����E���	5�8C*�H/B��"�{01�2%��w!м��a�I�@=y,��tA�<AMZ�L��:Hf���?
=9����a ���?=�h�<��.��Ո<�p����<�/�=����ڤ�b��;_c=�7��N���;.���)$�4��;��?�++=��;c�1<�<ăe��z.�أ��s3��ķ��.z1=�4=˚�����<��<�4=� < ���Z��b�8],<�m0=M�`�؊>=��<�ZE=d!K=��6=�O߼i�2�,& =�|�T0�z�='@Q<�	=����'�4�W�A=~���Ƌ��n����м�L=(�:=)����<��<��5==�����W�&��<b�<ԃ��<�%<$,�<�߼����G`<lW��8p+���
=��;;)�<������9�?��x�B��)<����L�c�<3£<��(=��=���o=�s�rlw���ѻ|�@��"�<�C�<=���s�`=�;l=t�=�=��/�9<��ɼ�}�<��T�li
=�值`Ȗ��;]�:��0��*��_ڻ�xk=��=����0�����<)V���=1b�����<]6=�lO<��ϻu�������M�[�.nM��͊=�K�6���z�WM�;����3�f���Ǥ��Fs�����E�"�[�u:7=Y��Z����<�ؒ�Ʋ뻪
�<�I_=g��<Q�<���U��
<:�&�0���d=��<�4=Bgy<��.;�o0=F�<)���;J=�9P�ch6<��2<����`껪s�<�9{�p�K�DW�xH�<��<^ۼ�)��+^=��u�FY���oI���<��-=�w��W=�̫��z=��%<�fZ<T΀<|�|�lm�����@�<my�;fQ@�}[�q�K�P�t�<),�t׎:ڜW=���Dx��)�ƻG�=o);=�G��Ce=a�=��X<�<�]^=�u�;B���,��I<�V�"n�<(���P��－3�j�r=0W<�[�<�3)<�0�<���<������<����v�6N>���=���a���c$�s�4<t�P��;��<�NX=�c�<��G��<�<�81=��M��JR��J��z=�!;�	u=#� �蓞���=6=K+=U�>:rR �Q;��pX���T=�u�<���<W��;`�!���8=ԯ=�'��W�y=+;D=.�<�T���a�(�b��FE��8�;:�E��*\�[]<�{ ���f<�#��?��h'���=����K���n�<��-<О�m@Ǽ�Ｕ�?��LJ�<��<�uK<L<t*��<�H=��R<.� =�Pټ��=�Fk�0e=��=$�9=}B �d�1<4��*<=X^!=��M=�ܤ<��O=dQ�B�y<��Y�3d��j7=�><� '��|��?g=p�/�v�U���#�o���~�<;\d;��= ��e�=�D=�6%=p�R�b�=�c�<<4a�O�<���<&�T�0Po�*w!��c�<l>0={�P<<{I=�1����90�<�MC��8=�"�������d��<��"�<:xA=��=C.��Ϩ�<N~>=h�`�R��Ԋ9=Z!0���$��;)���<]�=;T��x�S<U�=h��ε�R�v�`��C+�;�К:ۚ��?�=�e�9�8T</�<��-=X�;7��H�,=s��S^���_��릻w��j:����<^��<.�+F-��ȷ<�LT=��!���Ǩ�;.�5<��\?J=�/==��=P��d�@�}< �@�k��5c���<C�V:nM\���<�Aq���n=�\=nO�>�����<r���n�]<�T�<]�@�cy=)z����U��<We,�FC��#��՟�E�9=e��҃�<�Mn=#Y�
�<'��<=e�b�B�'S�;̔���=oʼ��?<�}�<g���z�`�L��%=<vd�<����~<��z��k���F��+�����"�p�B��z9����+�U<�˼�ϵ�7Ea��B1=z�8<�r����y=�a+<1�d=�,�<A)���=c>�����n:�� �|���fh�<�����b���;�?������['=!Z�;�'�z�<��<-��<�-�;ى=*>��y�0m-���h�R�c��m|=�v�<Jx�N3=��¼�5A���<�pz��j�|�2<��������0t��W��ّ<@V��M���MY=���&{�������8<�H=��B<&1r=�)��o��ٽE�DP���b��9�>�8�ۦ��p��fbS�ݕ�<`.�;��<(��<�>3=*���M�;ENC=uXc���;��;�$=�d�zn=(��<�x�<��輍�i=�����ϻ��3=�l� &��tI��GB�s9�<�B$����Av*�V�ȼ�6,�l4Z<).=�9r=p�(=�T;�A=y��H��<��B=�4=DR���9�<����0��<����)��B�<=��&ż��c���6=})��7=�й<����w��5 ���1=;���s=k��;I��;K��\(�Ѵ$;�ɿ�1�<�?B�t��QS��ý;N��^?.�nv�λ�=�9E=�����Ƽn{D=Y��<c{X<�ȇ���?=��{;�*����@����-<o�&=�����ڻ'�<8�nW¼(�?��Zr��	=��=�S��$�;��
<*��9$�j�N;/����L=JB_=��K�l��<AbZ=��S�籒<*6f<- =��N=��2;D�(�r�
jD=n�n�aڏ����<u�<�����\��-)��=����nļ�e<܊=�R�;U�*>��,�E��<LY�oԜ<#<���<C��:"�`�3��< ���X���q=���NT=�D�<�P�ݞ:=H,E=�<�셽D�=w�=�`r=��<�{p��_�;��l=?���jf�qc����<|�;��Fu:	��<�Ya= �:���;�*=W|�<��5=�`��4<IH�<���mh=7���¼o��8x;e:�sm�5�<V\�ߞ)<y�!�6�%�M[f<7�m����<���<��<��<[�#��Gk=Qߡ<W�E=Z�=� ˼�I=Fր�iU7=���� ��|�@<+�ż���ѥ.�;���;JT�<) <�y�������N��té�@�<�M'�XМ<J#���!=t��/�k;f�<+�G=	p�<�m <�8K=�z滹� ����=x�c;Z�o<5H�<Uw�.6<+ϣ<�z<{�u</�j����<R_H=���B����F=�8P=N�y=mf<�)�<k��WL�<������
9�X�<�6<�R �5�=���t0ռ�*<��3��+μP��<��3=l_�f��&W<<��O=��@����=o���='�=t$
�H��<��<}ѣ�M�ϼ-���Y���\<���<���:2 =øG�R3<!�<�I���m�&���H��<������9#A�b��ue<��_=|�R� ��<��ʼK?�"\s�~X�<��<p���?K��iz��	=�%X����"��б&=��0=�Y
��9;x�b����
=��7�k�i�b]y=`±��=0����I�<��E=��0= �F=f�=��*�F=�;��[��gb��N=�cQ=G M<���)ބ<v=�-z=��;��H��ʮ;���<�M<
#=�&=)[����,=&
���<�Oj�饂<\a�=��:�d�=�,̻S�����<���<�M=�p�<7;�<Y�:� =f?=���[�{<%�8=@��,�a��	%=A<�$�=��<�.�:�V�<�x���z;yɪ<nW�՝[�l����rb���2�Cc���5���J���]=V�i=A3���b;��<<���<u�]<�C =ҷm<��=W/�9���i%�<�|{=�ڎ��=��@=B;�;�=�Z�=�B&��P$=.�X=	���ZE=��=�x�:Ee�<���;�u ��	����(���<�t=��ӻ:�������O�;�ƙl�_д�4q弈|�<[�����+=O <��"�^�����
|+�T�[�л�<�A==��;˭;Я�=�=�k?�Pʻ��=4u^�{R$=�"r�X�<���:+=����W!�<�V���[=����m���q<��<�	#<
=:=��<��=���o��<���<��<h��<�`�<�&��#L<�D�ޙ=�n<�f-;����>=���K��,Q=�c���<A��;s_��i⼽�^=l�=6����Ǽ6#Ի��j�L���<�����x�����>Z=�f<��x=G�@=��(�����@�N~���dJ=e�3�=i�$I;L弑g"=A@6=V�t=l7���=`�=Z�˼��h=f>�<_購?N<�Z��y��<�P�<��<;��<A�D��gC=1��"L�j)=L���6�_�o=�=l!=~)<���1�>=�T��FK=�?=�D�V�{<Vw��IRH<h����3O<?�=Fn��>d5=nk=�	���s<���;��N=��<��+��;Y=�0<]Y��_q�<�=�<3�6<�X�-�D=�c#��WO�#!ݼ���+����V�wa5=��>=F�;=wd=XTF<>-2<S�����:ŏ�
�7������c!=�/�1"U=-|�D�=�riX=�=*RN=�_E�Qu�ՐM���O=<V�ʒ?<=,	�;n�6<��=���;l�:�aR���<R@=��`=��<����0=��}�+Ȇ<�7:��{��M4<M ���R���?;��<��=<ϼ2주zμ�&=��<�"���+3=T��<�A�<ˢ�=��:��㑼#�C��U����=w��C�E��<[��:_{u��*���J����<�~-���)<f�h<!�O=|��;o���+vr�|�U��x<�\=!bnR������=��<��	=�;@����; ����3�KD=��C�=�.=�1�S�B�7��M/=R�R<*μk�g)��c�;0!S�oY��`B�ϕ������=��a=M��@�;�Ea=<ښ�̖ۼA��E]�q⤼<=��N<�ud=u�.��M�������]=�6h���V��<�j|��e1��\�?���`�<&�t<��"=7�=b�!� pN=ɉ������/<�	=�;e]�<�5�<�aI;W��ʋ>=k<��t��!r�<���_U< &==��<��K���=.��<cb�<�P�>7J=�/=�ٔ��ܼp=�<�?���4v<�=Hs-�Q�=]�����9&J�+�˻�=�|a��켩Pļ��
=#�V���k=+H=B��<C��=1���WL�iA<<$����+��2K����,=Ƭ=;y!��T��l=��b=��=@zM��LX��ȼ��ռ^)�<�WK�[|=�8���K=�^=]H=s}_��:;�?<N�f���
=�T=4:=0|�;?=M�E���<=�f�;���<����S�<���<jڼ'7�I2)=��<��t=!.��$Ӽ�A'�>���a@��!D��������9�,���;=30�� �� %�1������<�6����K��;�)=�Z=3vμ��<�C4<Z�=���9����<��'���a=�h�	�"��T��B�%���?='U��Z%����9��]�K��i���3
!<���H2=p�j�m=�v1<��;o�<��)�/Ļ��d=W�<�=L�X�O7=�"�s�
~�%­��^�Ae��몵<�X���<����z,�yLl=]Ļmc���5;f�)=�=t�������2�Y����<
�<X+�V�ȼ�JF=Ѣ�a�%����<v�¼^N�=�}�<5Y=D���<���;�Xt=�b	==���<!s���^�;�Ž�&��}E�;ܼ|e�<�l�<)�f<�`�<ʫ��\��\�<�=?���<�/ͼ��7��<nGo�[���8�<D�<�q�2<�kļp?=1�ͼ=� =�6\���<�R��<e=Hd�<r�C�<
�=~)L���.��,J<���<���&�M��e��*�0��/�<O?ռnA��ᅽ��(��s�ޞ�<��޼J��iF=����n<�2�<)zc��;'C=�=�cH��}=DV�=�as<�1�<�#V=��<��j=:w`���ng��/�q�G���N=.	���������2~��$��a�Y=*e <�/j�`�=E7C�-\�<�H�d�W����+=m2�l#Һ����Y�M<�=j;��!=Z�j�W0���y���F=LWF=��)<�iV��"�=�;�:����=��;=@�ּ8���a�A�_��ױ���:�,�)����<9Qs<�0=
E�����n�f=w#4=�Dm�{�O<�U��KJ�������f@;��*=}�Ӽ��û�L�	��<'�=h� ��=�W�<�9=�<=�3/;i<�d��<����<��<�?��yx�\�S�}th= 9�<W�Z����el= I������9� �޼ХQ�s/<�M���-���H�w��yo==cټ�q=2{��ч<�V=�R^=�g��B5=����+`����;6D����<ǲ�����0p|=�������S0=�N/=�*=&���RX�Y�Q��Q6��dA=�e���`����N��:#<=�h��AļL.�<�¼^!<7��p�:<b\�<g3��w�<���<?�	�/����Iu=ou�;�� ��k=8}�:Jq=ԅ�<~��ڱ�;�T<	0�`��@�={�<x1@;���<m\f=�AT=/��<��-=��(�aD�<���\��<��C�N^
�,��<}�<�N���6=��<&,=<���u=�؊=�l=���<�t"�W�V=���i�c<��{<s�<�Yc=:'.<�<=���<��E=��ż��J�� ���Q���y= �=����7"���=�0<�,�"�=��coe=;`2=PV �I���e�?��-U�� �U�y<�1��1O�"Z�x]g=M�=b2�<�G��ң
��	<Y�d=�l:��j=���;]?ʻG��}=]�A=�i,�?2=�1�\�;��4=�%B=}C�<x©<W;�ӂe��$�<��j;14=xӃ��g�<l�4=��<T�&���Ӽ��c=4��;4���90��!^e��=<e�;�R8��|a�X�K�eK<w2 <��D��#ܼ[o���0V`�찼���<��P�x�;�lm=]j=[؂���*�a=^��WZ��xC���<�}K���;9{g=���S�<>C"���J�e ׼�#�^ǈ=��=+N]��屮LՎ<�"<ؿ�<?Q<�mk<v��;�(λ	Z-<r�I�R�}}���`�-���O=Vj=�Jh<���=�ͼ��Z���=/B��<�$����Db����<��X=uF���&�}�;��d=���4�9;�����缑�`�o]�bϙ�e�:�,���Y=@vI�GM�;G�E����<K����3=nD<9�����=WO�;Z/<���<��}=Вe=xo,=���=b4<���9�y����:�x�<@j=�3��x-=W���#�n�}=��P<L�#�~�(=�Ļ`�,�*uF=��<n!_=��=e�=�I�� �X=(�+�|=��~�;��<SN��|6�<�׹<N���˻��ļ!�:u�.=9��OWJ=h���<�<W��<��+=�M=1C=���Q|�(�m�ͷ_<�|=�V?����*�T<�K=(5k����;o�!����@'���<�|7�r%��{E=�cʼ�w&=QJ��� r���d�����	=h�= -=NK�iS=M]@<��U�U�;a'`���=�Q=��C�F��������:Y0t<�G�<�<��\=Vm��i�=D�X����<X���D,�F��wu=_Y�<��@��,����<R�<z��P�B=#,d� 1����j=\��}��HiJ�U\$��:	=?]=�./��i!��F� �9���A=g�=�=C=j�m<e.#���w=��s�O+���1=�����=tT�<8�*�|�<=�B�<'��=BBb=�w�<��=�(����z=��x�V�
�G=~]H;�Q��토<	���/�f=i����@��5�<l%���
=<u������<��<��=���;��5=�bA=�y׻��;��c=�A=7�<h�=kZ�<~��=>�=1�<VN��7M#=����Mb(=�%�g�E=Ǧ;�V���N29;��S:26�<]����Dc<�i=�tX�]N�I>��a:<r��Ȧt=��_<j��:O �3�=Wyu��
Y=�s�<��=!����<-.�<?rZ<��<��<�.�C=�;(=���;��;���<V��;Nj�<������0�<Ӌ�<!L=��<2@�K�2�O:J=s}"���D<祺��Pg�����}���;=;�P�<6$�<�٤�6�<��<�/=&�v� =>�9��'���^�o��;�|7<]����<*�;��=&'=��Y�wm��lY�<:uZ��A
��fּ�?S�2����j3<Vz�<~�9����ؼ��˻2�:�2ͼ��<P�������;��])v�����+P=7���28=�l�9u�|9W��<[�K�7ގ=њ�<I~]=��=Z<��<�lr�?�D�¨P����3$b;p�n��<�=�6��л�<_��,E��rA���u�:N\<0k�<��R=?7ռ?�=�=kX��h�<��b��<�==$a�<:\�?�?<q>� ���<g<!���	�J(�<��V��'���l��3�`M=�����=@�N�gʌ��9��o����&�
W�<P�G�ͤY�q�7�O�&�m=p/.��=,�=9��<1}����<s��Q���u����| =-8��č�6���uF:s�=�~=M�J�0ټ����Q8�<�C5��9oIv;bbo<��=B����R�0<��^�}�E=��)�:�c�m|<O�k=wV\���ۼÿ�<Q\8;5�;�T<�d˼��ۼ�gż��������o=K	$=��2<��Y<���jх�-f�<�U='�;=�2���.=݉�JJ==ى���ٹ<��{<�	K���J��u�<���=�=J2b=�䬼b���[�<;c`���z����̵4=��R���|���=H�<�=sZ1=� ;����;��O=>v�����.�<�C=dzǼ|��`u��MY=�w���=�1j���:q?�([=���j֒<��=4����eQ����<yJ�@2�<Q�>=��E<�1���t�<��$�H�	;�\����<�5>��}�Ȉc=%1=�=-��<��ռ��.�?�?�	���a=��DCT��6r<{t���Ny����$3ͻ�=�8?=��1=�=�?�<
ll�"T��r~=k.�<7g^�>�Q�$zY;Jŉ;�^�<�X����<�Q���'T�`羼6a�9��=���-�=$g����&�Įͼ[y�<�=h<���������<��<�~�<� ���r���E=�]�<��=9q뺦e�<����0Ż��μ���<g�V=�����+=��- C�ǒT=�VҼ%*n�� �;�-缯\>�	Kؼ3>;�"�;��<}��<9UI<\[^<�	���<уb����<\c����[=6��=Bм��<=w�5<�EC��c=9�R5<���>�_B�=1;l=��=�?K�Ӟy�+���ݾ'=�-2=4/G�h/7=��Gޯ�	$�<���;�=S�~=�m1=�=���<1O�W�:=]���N����<�2=�k���u<ᣤ���B������<��(��I+=�r��3>=�Ξ�өz��@g�m�3=�:=�^�<J�9If�ya��_ό;6?�¿'��_D<�;G�A��(l=3�a=�0=�1�T�j;ߨ��Á뼎��.6�<��l<�e=�&=j<_=yv<?"�<,0;�=��<�hj=O�@�=��R ='��<F<�V<lg�k�=���<q��d�9��߼�S<�U�����<~1�<��q��F=#�m<)����hP<��H=��<�^u��@[=9=i�K����<j<ػx�=;4����yh<\ñ:N�K=r)��l�5=Q�+<W1<y��nۼöb��;���Z-=k7���*A���Y=G�= ��RU+=���;l`��~S�c���3=>F�Sp=0	b��ᏹ!�=i#=ѳ�<�,!�qJ#=����<�N�2���_�Z�;��=��G���<A�G�G5��B0�n�V<%e;�Kp���˺Jk-��M.=�  ��v�<׼j$E�Rm�}G:�V8=��<H5`�c,���7=Z�/��0-=��<0.�����;D����b¼U�u�[7=�&:�YR���#=��1�� ;��f���*<פ���a��)�;��=�u;1�<Ɔ���-9ך�F��<��W=�+=q�?�|:X=��=���<1���Nny<�2]=�bR=�5= �z;T����A��;�-�<[\��?q<ʫq=�79��c��
]��f!=�h��3=���=◧�~�[�X?�h(N������_�dn�eQͺ��]��+�<z<�gڼ׸�J�=W�9=_�%��>�,��v^��4��qC=#�;�b=k[�<-K=o��;=}P<� �fz�<�J��[��<
'�;�<��D�_6ٻ����	=֔=~���4|5=Ż�$�=���<]M��A�<0JM�#RI=#��M�һ��<R�a�[Ɔ<?$=��J�,䀼'�h=��<`tK�xTM=�Q=_�<��@�����a�.=�l�4?=�PP=�}�;F[%<�W=�=[x1���<,T=����ӹl�G����m���<�ف;(�C����<"⵼ ��<FM;=���.�tM���,���U*=�!;��2�<8�S��a�<��<m����a;��5<��=i�&��Լ&�@��$����c�����:�<�Ke�]u�<+�0���ϼ��=��q��31=KP=4 \���*=��"�r^��B=�m<�P���~⼄Q'���Ǽ+/r=��)=+
2��-8<5�.<��Լ��;<�bڹ�����cK����vQ��L�<��¼�=�t����2���L�='�2�Ę<��V<t���-G'=�E=S�'<�� =u7����7�[��^�f<��:���<wP9=���;Ny/=�v8<}2f=Ӆ�=aQT��=i*�wƐ=v+=N%l����gG���輺�i=�%=ۮ�:L:��wE�<>��4.1<�W�����O����<P����rV���A���<�$ͻlo=eH�;�Չ��-˼js�<5$�<0�:^w�<zO��!�</�ϼ�aż�A�<��z;M�<
���ٻ��=ŴB����� 	=�0���@=�O~��Y<%�C�0d�ܓ��=�P�G]�<O0Ӽ��`��jy<�@E�;���G<��:��i�<I��L�p=�e=�����U=��^=�_%=}�-=
0)=�J�<;�*=�N�d�<��;��=�w��8$=V��;��l�B4D=�ah�<����ϲ�<!���,��<{MF=��=�5�<�݊<�^'=˙p=r�*�T�<F꼎�I<R�b=��q���L=���l@Ҽ]Kg�qL�<[����*���X;�d�;;[~<�����;��-ȼ$���Z��<��7�Sr�<S?=���<��;t�"=WG3=���!{��w<��$=��<ê1=,�C=��ɻ<���ń-=7.�<���#� ��o���-�ީ���<�����f=�IE�����Z���Z��٫��#Q�/x=��<6��<���qaJ=���<�<24�� =����:	<M7=ؼZ=��<�/�<Vʛ<�;=H˼������ފ�O�<؃=��3=�ja<ӊ�<��,=W�<�sv=����&�>�<F�0��y�:�⼈�L�~eY�2�<G��<&/.�Jf=ܘ��J"�E/�52=4b�<��T������.S<z��t�+��Z��8�)u=<���#=��a���ؼ2�=�
=}/�HT:�*δ�~i���d����h=k؍<��<�ڂ�g����}��6M����<�<��<=^�Ǥ�Ъ<�k�=ˈ��~�T=��4�g���/�<��D��^�<��=�{@=�Κ<���&qC��C��,�� H����<�b����<����C�<
��<$�=ψB����<n�I��P�<{-���1$=y���@|<$� �A[�<'k�<c��<-%�Le�<�]Żu�l=~mM�%od=�TF�Xvػ�r.<�q�<�15���e=�k�<1��t��'e=BE��|��a���=#1�<[�m;U��/?=�T��H/<7~�>�;�»�a3=�Du<:X��ގ�G��t@F<�;��.�k7=��D��rf� �m���[=�5�wp�<��'��=�P�"&������<��I��Mr<�W:=�@L=�nż��U�E.j=�����=�1Լk΂<��?=����b�A�Uȇ��.���L:�~q��6�b�=��K-<�j������.��������F���=�b�<� �̮��m	9=�S�U�|=>�y=�8�;]C���ϻ�	H��}��S,����/-�<�f.=�W�<�1&<� �g��<�3#��'_=l4���Z<�Q �߲y�>-��ӌ<�,=��e=�>�<��8���
=�浻૘<��=g�<a{�����;�=��Y�س
=<oX<��p=w�=4�V��1r���+=�zܼ:�s�*� <R;����a=[?R=������^=XIS<��<�l��?d�������E�S����=8[r�R�
=���<;=�M�<�G=Y> ��x!�nDD�����"=kQ[�H�k�dw����w<*J<z����9��x�p��ͅ�珁=�GD<��ǼG�_��;�=*L�IO8��V�!�=j�m;N�H<VQ��/4�;� =�DV=�p)=���(D=G':=ܷ@��(`=b��<n����=b��A�M=V���g���=��|;, ; &^=��<$h=�Kj�_1N�d�ᚻkD2=l�7��W4=T۷�=<< �<I�m<�=�����*���I=κ�A����<��F��&0�>���L�;�A����<,s;=��$��f	<ӷA<�D��;g3=��"Ի�o�� P=ÏH=�8�<:E= ��<�3���<Ϗv�X���d�%�����Q����9�P�i��X��x�ԼI�<�5{=�}t=����7��:�ؼx�H�d�#��2�<�� =bU�<I����<�A��<=�ܼ���:B�+�<Z���}��ۊJ=�;b�'=�U';�a.�y�A=̮����뼜�_=��C��3
��K�;�
e�m�#=� =8/׼7"@��<��F���O��Z��<r���{�<(ü������:6�ʼ�׏�/@; ��<���<�'�M=�9��?�<�rD�^]���6�����o�+=�~ =r(4�����#�a[;k��<��=�<�̔b=��S�:p���8=[�::Q.=_��<��<"Y+����<pNn���j��ui=NB��4�x�c=�%�<J�J�|(n<�X=�C�
YK�I11��{$�Eb�<�����b�<��=�J6=�W�<0�M�9=�ӼU?��F�Iz�v}(��1��k���=1H<P�>��XZ��63=o� ���<@ÿ<Fo+=%����}���S�c�f<�/i<�= ��{�<+���vE=���<�A�<ݟ<`3/�2��<��z=��м�f*<�e�<2}�<��a��c����ۼzz�<!-J=@F�;�dj=(�]=��3�:����!�@���K�*�==�O��a��<��G<�k=c�I�aԫ;\`=�낻Ѿ˼�c�<�����i���T�n�J��F�<��+�I'=�8=о+;�L����y�M^=Z1�"�<�!U=�[��n���2��缢(��kU<7G=�=�=[0=��<X�1�p{��.=�;}���b�!=�4u�/�=��Ba��B;��=��������S��i�*U=��=B_><�q���M��� =��<E;����$=����Z�<>�'�eoD�ޝY=R�B=6�q�ڻ�g���z�<B�P=��<��=��?�܆⼊��<j�;�F=b(V=8|��l�.��hӼ��G=�$6��>K�b	<�l��{��1���<����?�=Z����=�G=:'�<f;żpa���U=TR���m�<FN!=b�<:<ǻ2�L<Ɍ��^2�+N��\߼r��<��E8RF�<���2\��;�¼���T�Qǻ5����
=���;U <�P��X�<=m�߼�;�����=%���5�E;��e�A�׼p�-��&���+�:=؀=�O\���/i�=2��<�=7����<`ݫ<v�J���R�ć<L�	��/�<$�X�uI����K;=(��ʷ:-TK=G<���<fV�<RaN���<}�9�R=��7���Y�Vw0�[	s=(1����<�G���r��K׼Hh��L���AN��p���<�����.c=EE�H ����<�)=�K�<�[=r���|Bp�{�]=;�;==�9�'V$:Hz&�ll	�^�(=��<���;ʚ"���f=��,�֧�<.Ԣ�:i� y����޼���<�o�<� c��G�\�=Jpc���!9�Hx<T�ͼk+�f^E=2�ż[�<��k<�%��i�P+=���'~=f"�;n�=|�C=ɴ���;�<�oP<�� =:<n)�>n;�]���o����$=��;��1���<9ɼ�3�<o*=d�c���D=
^��qJ����<����E���༆tm�H�]� �5=�j7=�Mμy�V=��<{�<�hS����<Bpȼݠ��������X<ǗZ=C��<�ӹ���ּ��:�P����<`4�����'=�c˼R�2="�5��k==�^{=��;�=(߼�C=e�.=�t�<�����
=a�D=����|���Z=� �<�k`�����r����^�6@�ND�nz��w�u6�;�Є���f��u�<�#�;���<o+e=�wy��am=�T=��<��-=cG5<7�G=K`0=��ͼP#/�4�`=�~:=x[l=�n��4���[�=.�^�= �e=��D=/��;b�<hgQ��=�<gi�R=�A8=��6ī<{)<� E==��8��Ԇ<Z�<J �<'�]<h	�<z�G=t)��ѩ�.8]���T�2�j�Q=`!���!�_6=�m�:I¼ߔ��!�.�s10=#���'=X�W�Sh�;��n=�3D�����"���fQ;��C�X��<j{f�Ͽ(�Ⱦ�'/=�2��\�<U_�<�QK�e?="+��k��-��<6k����&=�Bo��������d<=|X�8y3�}��<�b<� ��b<�(N==�`=��:���I=
�#�*W=��$��5+=�G�<of_�i����[M�N�=I�� *��o:���3��|�<�==���6#��B�<��!����cD�8RN�(�ڹ���;�9=����+[��"�h�4����6�u;Gj�<e{�<�Z=q3�ٝ@�}�-=��%�*=P�컈�F��/��P#=��!���=�.=��l<O�#��k��|�=��Ҽ-�|<�P�<�L{��+�<��
=V`�}==kvI=F҂��8�<��<m.�<�0=P�#=t3=���<�<3�%�,"�o?
=mx�� �<�Ld<���<�\=:�A<㙣<��7��c,�A��Ϛ<0z�����p=�����<zW_<�n<��=Yv�<Y�$ߍ���<�C�<��E=�o�<�+���=�6�p�����c=�m��`��㣼c�<�.�|��;����*M=Pa�;:���-P��CR��r�<zļ�q��C�;0��<]�_=���y�<���<!E=��@�(�_=�Ɩ��KX�� �<��<c��<k��m����Q=T�~<�1C��+�<�慼�k:��*=�e�re���T=O��Z�2<%a:H_��/t���=R�S=��<�œ<�<ۭ�;�vQ=������]��GD�B�K=�f��:<�|<鄊<^?<�w��=�sׁ<	��j�ػܗ7=s@6=��9�(7d�=f����<=R@�5�=9�<f�,�~y;�u�<����8<:T'��S�$��<&�G=�G;�)3��'�k<dN��<o�'=N#V�NS(=����!�=n��:�D=bJ==;������8-��d�؎4���9�7A=k<(��2��Ȟ�_"=媿�\9˼�I�KU�<yj�=��|=�s[<��:�,�cGD��:=z_�͊�<6!ؼ�-_���V<K�ݼ5FƼ�`>��+�y�z����<`v�v�/�7p$=�g<���	�<rR�=���<I�C�{k;�^d<��a��jV<�,=�s<{US��������)
=A���t�;�i���1=TZ<Ռۼ��'=�\���M�Y����;=��;�:i�D��<֤<��<�vg�>�&�m�3������<rH�� e2�	��<��z=�Ra=�79�wO=Q�ȼ��_=�"	=�B?<�Ќ�L��<ص������]�#�i�x�|4w��H���~�<�
=�+��.Td<M�ݺ�g=�c�\�ϻ��\�έ	=��*=�V߼47�<�v�<:$�I�8��Ls<�X=JQ�<A��<�,�������<!a�0�];>S3==�~=�X,�L����%��	o���<�� =j�+���]=��?�gpP=2�;hv<��F=Ui��Sv�����x=��l=.�-a;�DƺM�׼�F�d�<I�b�Z�����A=�a���J̼�]/��~:=�i:=�3�<�W�<�sA=�@>����8P��L�<eO =��Ἳ�v<��3����<I�j=�\���=�a
<J�<�-=��	=�=
�m;S�6��[7�!ӹ�W�<Ǉ	=o4G<���t�<s�<cd������ =��<�<�@�cB,�⛹<o�����<��+�j�#�����-޼�p~=-�=�2�%>�@����과�����������<��m���r��������K=�?��~�U�#�;0M=�qR�1ɾ���˻C���qs=b;��2=��ͼ4	w<?{5���~�ゝ<]�M���R=���:��I=��j�us�u.�^k�<?��:Y��;қ�<&�����<��<)߂��ޢ<��5=:n���԰;$>_=hm��e_���;���<���:��<bk��B;#Q��9�����<����e-'=���<ߪ~��*w=h��<\�>=wp��r�μ���꡻�NU��ܹ%�8�*=��P�<+o�����;=��<�0*=�޻.#=�Ѽ�$'���<-�<{0=�k<G`��ɧ2�]F|=��`��E�[� =L��<�&�<i�c= �?��_=�<"�]Ѐ��8=�$���Ƽ�ک�1�;۷&�f�>����q���B��|�����;�a�(��`�ټ�UE=Q�{<=�m=���<j=v�=ީ�����<�<�!8=M����1�<*�:=��#��<��[=y�C���C��e�׹�~g˼j����e�z��;|��/�)�
�~<l���
5<����<�li�}�=Mߊ;(�ֻ���<T*(���F=G���3��<�j*��  ��i��!.�\�A�0�Ģ�<)�D3�;�R�����<�^=DC2��O<�"=w)L=ӻ�I=M��<�W'=4 ��$���V�-n�e�e�"�!=%�"�Hf�q]L�m�<,��^�1���<�r�
�"�=m�	=_?=�H$=6��;��=ӞY=���<-0Q�7�s�q�S����TX9~b�<t�n�kH�����0�V&��e�vv[�S2Q=��H=�=Y<�<)�"����<���a�c���L>q=S1�<?���Y< %�������<34;��T���]�m�=��=�64=7���+h;H>�g��<3�;=����U����  �C(�;��x<#�
�R1<A� =��P=�kD�E�<�C����crU��^1�ʎ�o{����;��"���5����V���#�/=������A���	��/J��T-=� ;<v��<���<4�Y����f�"��=K�ꮚ�MD=p�5�;V=U��;�N^����<�u;�E��;���p�;���C�C�4�mk���N��[�9̓�<�� ����(��;���8����?���T� g��/�<�F-=z�d=+aԼa�K��;�j0�g|� R���k�:��<=0L��8=9��;�=�Q�<9p�<wP�<ّY=t  ==�,���u=�Q9=�.2�7�H=��.=� �U";�> =��<��4=z*�2�̼����
�ʺ�<g6=ѭ|������J<ąG=^�Y;qe=hD��^�?=���YA$<�A���k,=c(������6;�6��ow_=��;�)�<"�ؼ���<#�B���T�Z�̼E.J=��]��j�<����f�<<B㻆Q=	"3�X��<wX��5�_�59�Z�Ƽ��=c�=;�+;=^S�A+�XAC�V�C�@���g���>����<Y�c�I�5i뼔�;=I�żF��<�K=��>�n�=L�#=���9h�������@�Te8=y���P]�<���<�1<��]���B���o<&��;<g("=����?v=7�=�[�����36g�דt� ��a��<,�h�b��n�<~���;��2ȼ�H����<�!��S@��T�;	ż\S�<��<�+0���<��<@�<�D��h�N="�=������<�U4���¼�c�< ��}���n���*�P��<$�2�µ,=
,8���=�k��גb��Cy���Y=�I��fY�=��#�H�I=�+���Ż�<�2~=؈d���E�p4�'�$��%�g�/���]�G`����d�H��[�f�v��e�Q�D����l;=�!K�U�3;8�<=P�����<+w�� 9;�I<{&=��i��{��G'i=���Q}Q=We�<���-E�<uo��/k[=���<549=$#i=�x����<8�k;� c=S���U����[=���>�<��"=��J=d	w��	�q:�<��<`�f���<h�N=#���U�~?~=q�Լ�=<��;Kk�œ�<5�T<v"n=��c=��~��A.�\�<_�<�����e�Z�����`��H�<F�<Л⼊�n�ؤ�<z��.��;�I=zo ��)=���<���=�D�wq߻W��K�T�����5�<�{ �خ(<�~Y<L��<x=�	�ռ�����(f=�B%=x?�#�T���w���<c=)(ؼr�Y<F�<m*��rw�=��w�d�?���<��<�ͧ��[<�WP����<y ��^��#a=# �	�뷣�S=�Tx<��i���м'i����<�N<Jr�<�q�`:$�i=ԉ�wQ=h7,=/'��i��2�{�F=�=�_�<�I�@{o��h�<z�;=On�<,m�<���<��˻�
=��<<+;�<,=��<+�<n��^=�Q�<�n�<[W�l�?=�컻�^�h:�$�����l-#��NY;W{�Q �<�VH=�3T�`'�F�<�)��D��s����l#=���}��z���e.=�c=�H�;f��&�Ժ��7�B�\�_�a=0�=��;��9=��g�<:�<6�
=�:¼5R
�{���H=T�<*R�lU��d�������{���r�Y�0<�6=>4���ķ<i��<���`xT�l�����蒼���6	O=�xм��f�~����k�=Tr�;\?�<]�L�m	u<�s�;.�6��[���=چE=�[�<��n=��+<A�Q<���;j������}=��]���d�.��8�<zT��������d���<1��r J�l+=��;��D=��M=�F���C�;T<�<'��<�A=/�=��b=��w=���� 1���Ȼ�3�<�`�:0��P�<����O]����ټ�>����=ef�<����2�ɼ�x򼈫�<�G=�,����<�����X�,�<���<9:=�!=#�]�Y���)=�:=�����<I�-�pf>=HŁ<v����\1=��0�s]�<�R=��;�(=Q���<�
�$R���K�%�	=��=K�����:�Ok=Q�)=`f=6a���!�=#��J_;��<!�m��&�<i&޼����D�<N����<Z�����<흨�����ʞ�<�ǻX�s=�r�G�=�i=�FX�2�@���t=�u���r=�d=C�4�ݝ�;��μ�d���<n��g�Ļ6Ď����9m�<�o.=i8�Q��n�<��U='������Zw=�IG=��~���=\AD��I(<@G�=����!�;&|_��s�<��ü���<��y���b<�f�mw���J=�����<�-�<�Hϼ6���L��<��U��ǒ;F�Q=�H�<[d=gŉ<�+��]<%|<�T)��I�\���E���/���N�r�@�|�k�ĝ=l^t��jZ���r�A��<�V|�{�<gB����<i�<�OD�?�u=�����4�Cƙ:BS]���J�	*<Ń{�"!�<���{�D=�Me���]=���<(�<��<�2��E�����O�fʱ;X\��V��`�"�/ �;�κ�"�<KK���5�Ñ�<M��<��=�i<3p�<�=U=�#�;_�D;�S�w������Ho�A.K������Y=8����<r2;�9�}p��G*<)_�=>z��/����M�%�=�q=��T=�dm<V�3�圣�O���=�T=��<J�=zIM��X<-z�<�$����&<�qW=���<'\=(B�k	L=KJ��\=�d���<s�C�#Q=KLĻ�=�jn�9�J=G_�;�rR����<Ɲ=8����6��!;y�O�+=��{Ǡ�v�=��<�;!��UK�t�1�_澼g��<=-�<�v�<��<5U#=G{�<_�V=e`=W-����[��/޻xf#�,�%=a})=������}�<�H='�0����<^2���g����=)�C�+�� =�w�Ss����X=� /<q�%=�P=CR��� �9i�������,���=Jn���J��P=�ͼ���.��:m �)[(<���<}���;q�j=m-=�=߻��\I"�Ra@=Gț;� S��;�<9:����q(=�|ͻH%�<D�<Y��b.<?��=�z�;�8��|	=���<NH�v�Z���<U��<c�=d��2�d�x8u��6S���I�+t���� =�<^�Լa}*=�+=g&�<N��<�� �(ǐ��n�h�^C=}���F ���9���꺶J� �;�n<���ѧ8�훶;��D<؊��:%�<��7-<�1=��=�h<Pnh=��R�@��<���<�H,�j��:���]� =��=� ��$[=ȧ=�`�;iw�<�˘<��;�	�n5��5���_�;)'=��b�g�S<Itͼ���H=�W=�"S=9�S=?�<�dc=o���+@2�C�ռ�o'=ª��CѼ�S�'Z�>�=�X�MY�<�@�<�5f���;<�<�;�<��Q=�Ae��ܻ�,�d=Mگ�a�V��p=0,�7"]�w�/= =��_�DL;��= D;}ݼI9��O����;�����<��;�O��;kBM�C�W�(c�� ��;=���<��$���;����"˩�C��;p3��hGB=�V�����<T(d�a�1<�!^��=aI��\�==h���ڼ���MK=�@9���F=��7�ƃ�<�ga<��b<A�V�6C��;����C�O=v�:4I=Ӗ<<����o�;�����p/=6q���Sڼ0T<�xd�/���`%�<������P��;�;"Hȼ)�T;��˼�&0�]΅�Q'���t���g�
�2�Vk=c��G��t�;%�h��g����=K�g�i �;>����H���<Ŵ����.=���
�&��T���z<�&Z=�Ph<~�|�i����cm=]�G�ml�;쀚���e���2=�߼�1�" ��pF��vu:xCA:����c=ы�<��^=�ɀ;�i�� ���Q\��м-X@����<�9�=��< ���U�%�$�<D/<�P��'@I;�8H=�ػ;�>=y$<��h�ᤖ<6�N<e�n<����ъ5=����)��Uu�<lu�J�[Ǽ*I=�u��Dj�<�A��s�g����͗�g��9��H=���8��>���;`殼�~�Ҵv����<N� <�;��	=�N;f�q�f�<��� =�伡��<8��<Ӳt=4y�<�" �SX={�� �q<WL�v�z��}W=�&@<���Z�<�t=C�*=�7¼.���cK�����K�<uxc�V�`�G�(=�<Ӧ�<��;��<���:�,E<���:��O=�fP�{GQ=J�ռf=��������C�q�3�h���O=y�;�Pa<�^X�6_պ5�<#��<��J��~ٻ��L<=�)5�Z�D��D4��qG��﹯�
��9Ϛ�<=Mĺh�<�𿼅gl<��#�����<�<�/1���!=�6뻕��(�P;��Q�|ͼ.�]��vl=��<Ɂ�<޳�;��Ǽrc�;S`��U��;6����<�<��>�<�p������=� =�N(<�U<�%,�4�R=o�<
x<�'�<X
��w���i��{D=SE��p#=.U�Q��M��<�S
="	��P�r<c@�<i�A�\�L=�"<�b�S
�;��=V��!�;�˂=��==�����=�@���x�������<»�<^�o<:=q��}���')�xD�;}i�N<ڭ���c<�P7=?g=s� =K|���e�fm���<�V�;Ny�[=��k Ҽ@�w<,lw=��D=>�!�OU=i��;
�;�v�1=��;냐�Sf ���=��<�c������ľ�H�����{*�p���T&��X�E=�d���m�<��t<��m�1�}�M�<�+=�y���N���(�M'��j�<oB���V8=���p=mm�;�ɼL�<II���DC=���<F�ļV!弌�<���<5�M��� =�6ʼnd�<��D�>��7=�df=�52��}=����=N:<&�P=�cм�^3=�~��H���<V���%����ᤳ�z�.<Pc�<��f=�$���Y\=2;@�3�==Q�=N� =V�h�$���<=�B�0���\���m����U�?	��hB�|��<�7<�!=/�0=<�1S���i��gw�h��;2�)��u�<�G�:�J=b#�<+=r^¼�^="(��t����ڳC=����A�K��<}�_�o=J��<�ش�ڟ=.8�R�J�k<���=Ll5���N���E���Ǽ��)�i�A���<LSS�~G=�]�<�T=au"=��L���;�]l<M�<���<�Q�<��efy=�rۼ��;���<��ς�<:�P=v8X����<�F=>��:X�=[�G=kֻ`S=w�N��lc=ߜ-�֡<��L<��$�˪����꼇+�<S꼶�����;)�Q<W�7����=��ٻ����6r���<<Q���a=����bՁ�x=Իц-=��0=��'=����S=.X���<V=.�ؼ����c��(�<�4?=��o��G"= ����O�ų�<���/���<os��������t�<ƣ���;=� =,�1��.�CXH<��h=x�;=�{`�1%<@��<H.h�rL=�|'=��];��p=�Ɨ;W�T���<{���|}�8�q��L��C�W f����<9v�;��<è�<װs��n���5=��M=Q{�Y�=��e��X�Zw�<��n�&=��G��v��Ͷ�<d!��C�<��$�[5�=�_<o��<�c�L�k=P�[��� =�a:�=ՠ<�s�"y���<ز==�<y�B<�9�g��!����=�r�5�C=�?�;�6=��};.�<vi漑�9:�(�<621=���;z�=�I"���Z�v�c�?=ÿ@<-9}��m�3�)����<w$=-x =ݗ��~#����<I����M==#�=��.<���<���<U���L�;�Q=�:Sն���W=�EC�~k>=@�;������ѕ�࿈��~90���ż��y$<Ġ����I��Jl��7�;Iє�o�<�>=/<b�Y='K�CE"�AM��W��:0E�0��<�,Q�\I4�4p�<�#��q �N寮�m��<YM��(<��Ž�NZ�<��<}W=N�"=b,<x���2����;!�;hZ�<��=��<�8�<��;�Я<�<�<��ּ�D-����� ��<��'=9ԯ<� =<���;xf�<I4=g*<{��<!c�9�-�ێ�<u�\�o?9�/�[=�H=5g����<�N!=��Y<��f���<�KH���;��ʼb�1=��i���	
=KhA=��X;ynM=\9T�e=*<��/=n�z��E�G�<}�<��'���x=���FƎ�/r�������,Ԟ<��V<��@�֙����;�(�o��>��<)�
;ea<N�<G_m=� �3��Z#M��{�=��P���E������"�=<�����<=`= ��9H�����5A=R�=���]�<�NR�<�3���,=�,�W��<־p=���w[b;�s\=��.=!=�i&�'ef��׋�C_=�{��59����M���鼋	B���R�y�ɼ�N=w`��7=����t<�k��>j��ͼ.w�=����C���=Ә+=��V;�9�=S�����?=��$�y6�P��<�Gi<�2�V+=8��{�<�F����eE+���<���<9?�<���;e���E-�`�/�ul=�7	4��Q(��6=��%=�o��a���m<um<=�%G=�Ȟ<p��/���D�:�z=�;ςX��	���,*=1m^��x>�X�/<��\<��$=�g�Rǽ�01���/6�����e��q4�<p�]��[G���7=by<~�<In3=Q�c�ؓ�<g>8���y<�~�K<c�O��;{EK=�Xm=.@t���&�ya\��RD=�[�9Qy�
�ּ�h=��e�=R!7���
£���_�=k~�62O�$-}�z#=�\=�}�;jou�Y(�2�=S|=��i=�Q0=	Mû}.��ہ`�|�.�S�c��{���|�;��������!=�p-��X@�63��Ʋ;g�=��<�$�<sP�<�,
��l��o�>��T>=O�<.�F��me�[�<ZNҼo�� +���z=�f1�e=�pf=�^ �F���m�����</�<|0<Yfͼ5�c��<��;=6R=�~!�CQ��P8�<R�=x7�<��4=���<�*W=Ja<�$i�.-�G��;�{�&UP=��<���<^�=�.=��)���7q���p�>KE�+e&�=���1=+��<&�|�/��<ȰG=�����;T�==�ņ<i�&=��<N��<�«<�Y��u�=��	 =1,�<�F=�	==�"=�#�<�a���7=�M�;��f��}3<�)��N!(=i�m=��=��Ӟ= .I�E����5ؼ|C��{��nY=H�,꒼��b=0�=���;���\&&=?�<���[�Z����<���<*�	�.<���^�<u��f���e����<���ŝ���}��쐼��=�:���-�7GE<N�7=�/<��:�m}��V�<���:�;:=�z<=Z��<FG�����h�nI$�O�v��<��F��&�;hm�<�R���U<�r�"SI=o?�E���<��f=����T%=���<-�=!L�;���p���ߝ<��@</�<�{7�h�:<-�ּ:=Gy�<l�����}�ݭ@��3F�%= �=C
e��;�zJ��{м$�i��.=��~�<�c�<�@:���j�K=ص?=�V��E=��{���`��%����<(�<"�Q=��\����;�䶼R[�<�x�P��<�}����=��<`	6�;�����;���ۄf=V�|��j�;I�E�C$��^o��5)��3=���"�\=P�f<�`�;Ҙ=j��<�@=E^X�� �<����y��5 =����4�z���˼���$L=5�H���@���<1�=�*�:���x��𽱼?� =BI������%�A>Q�{�2=��r�Dլ�̒=�E�<ixV�1=���m^5���`;Q=�	�:j�:-��}�	������;nSN<�>�<{H=j��<��E��K^���=63�<_1<� =��S��P��J�<�5�<��M=^�=��o���;��g'���T���=�=�ejٻ��=2�D�~P=MdO<�^Z���9��P=�l�d�k��B=:���Uc=���Z
��K�?D�� 7�PO��i\��F�B=u�ؼ��i�<�;<�
�<�=fq<3N%��v��T
=��;#�=��m�{|
�����VX<5�B�T��<�^�<�RY=�V/=u�a�
�����u.��\�=ҷ�{#�=m�@�'S�:�̺\����<y�t)=�o<jtD���ɼ����c��y�s|�<m�<O�E�<�+E=C��<%Js=GI9�N���X�w��Q��q�:Z'<%�S=�3M�h�Z=.��,�B�v��<Z��� ��;TB�-;
n��V=;ɠ��/<<.d=�#W�Ӻ�<��W�uH=�V���<�	N=�.�!���&s���׼.k)�����b	)��A:<�嶼N�&���B.<,M���>��}-���)=մ���^:�������޼����Fb;��=�X=�=�<�5�d��<N�[���������D����=|M�<�=�^�����;'�/=%�:�k���U<���K�j<���<��[=���;��"�޺�;l�=�G?1���;��E��(�}��z��������]�K��;x��D�?�a�@���x<I_=�4�=����Z�꼗o���&��PY=C��<4ȧ�����{�ͼS}V�!#=̀=��J=ba��i�
�S�+(u=�k��T��G�<�G=]�h�/>�Zf��-�<!�"=��/���F=��F=P	O��*��d&n���;f��<Hs��o�𼃴=j/=�N[<�
켵������<N�5��wC���&�v�Իn�<�;=�핺'?�<.����4�<tH�<�ۼ�K=�>�<.m=�T=�W�:Og�<&
�W��<�H!��D	��Ý<�܃��QH��G�;��n�Z��(�;�>=H�W=~V�8��;	K�;�L˼�=<�ȼ�gZ;މ-���:��:=��Z=[*���=�6=�b9�x��<��%=�P=y������@R�<Y���I��6=G�==�A�;�P<�u�p���ON���;ι躗[�<�w�<��ܺy-�2Ц����4�ٳ_=��=��f=��;<q�����B<[o׼<# =�M�����6�'��<��ۺ�=r�+<o0�;D�;�H�;I�����<ٶ���f�#^9=���<��i� �<�e�����LV,��^={��@c=%b^=T	=?��;oBd�?�=�}��_Ɗ�����˅�<�����;=]^Q=��<	p���|q<��<��B<�C�>�<�r�x������H�<@���=<�;;���&�<*�ϻͫ�h3w;M�R=�p��$=q�*���$�wz;=ttK<��r�Pۚ<-�0��˕N=��G�u��}pS�73��l=��=���;�)�<�����=�=��%�}=����,�=��ܼɣ�<��(�<^l����;�K=�����s-=�h*=�%��<n�̼Un�����3�"={M=A���/�<t�;b��c&M<m�K��gd�N``��Q_�g�]<IL��f=w�F=E��<��e�{��;Y⼻���=�,*�R���3��3'��V����/�"b4=�=�X=����l���&�6#,���;=�+=��=<�~;�;Z��=)�`����_z<�`:�X�><�e$�T2��� ���<��W<��=�<�I�\�@��[���V=����(��8�˻
��� =�f�=�M�9�!���Va�I.=�w����8��#&<u=�#����a=?���+N9=S��;@+P��9m�e�=i�ۻ{Rk�d�<Rr:��;��	=Y#<.!�����e_==�:�<�g��=��>=�D�|<�i�\=�e��9U��q\�,�����<%�	=y?�a�n<�"�<=H|a����<6Y<g�P���I=�s=�oj=��-���ӝ`�^�'`9�R.l=��h��W��TK�Qܔ=�z<,�`��̈́�����G�<�|K=Q���u,����)�E�<�� ���i��)��4�����~:��O��.=�,�,EѼx {=�ٍ�?<�%�h=q+O;K�;3��<I��+=f���Y/=�R,�)m�|T<�Å����< �J<ta�'��<x�<��O��<&= h�>sԼO�;?���[ꩼ�O��=i"=3V=��<�1H�0������<���<��<�z�����B$Z����� ~��I�ȼ���|`��ZF=�0=7����h=MV'=f���[ ���a���C����l*`=bj������o�<{_=�a`�f�C=�gQ�V[���
�=kSK=�C���<��=�U�<}�;0K�]�=�]<Nl��l���R�<���w)�0�+:�/=+�e=7=uv[<j�A=��=�
==�
=��ü��?��{��㷼��� �0;�&���=��?��4.=2=#�ܺF��Q�ͼ��Ӽ5w7���=�b¼��0<q7��;�<�j;>��<��={��<��;�(��_�7!^<l�ļ��*<��]<�<��!���<-&����
�3�\=u����.�R�o;eP=x������P��u»)|�;�l��Ib:dL=�v�<~/<�<D=�������=��8��Y��N<�W�����]=�7w�L�E��*;=YZ	���ļȯV=���<��<<1�a=�J�fܰ9d�<�f�I< )��)=^��ti<8m�<�E<�h=u���+�<ʓ4<�]_���/�<d�O=,
�k�a=v�F={��<�gl��"��(=�]=��<@a���)�<3:�+��K;:��c����<��c}=��P=�sQ��/3��S���<��:=+ ��)��;;^�;G2��B�%'�V;(;do���f��$e�lP!��a=\>�<�����U�ك�;}y<���<?i=v�E���v���i=o$���w�7=��E�{<-��r�&=en=|=���b�E��46�m�	;*]�;�=��Q��=��=��$�tj���@H�6V��}}7�،:=�����>��<~��<���P��<�jO=~�<Q'�<r
ȼI�<c��O./�7�\<,�<y<� e;q���R}K=��T�R�0��-ۼ��
�(�=���|̼v�ؼ��M�~�X<cAҼm� �R%�K<�<�>����;%3<��W=O�=fQ<�\=�#R��=����^����<j�*���,=HFa�����U.*=6��<!�ļ�N�<J|<<9gj��\=y��$�q<b��<
�m< =����q^�;���<��I=��.;nQ2�KO=�_�=t�k=~�	����<��Y��m����%=ì��O75=�+\;z�ϼ�p����;��=;e� =��U�ں��� =����<c]�<�b���ȅ�H�F�y�j��]�<ֈ�=-���"��ℌ�Yu��;=R���n�������a��<��3��,i�2v���=k��<�7�gu;���Ǽ_%<�&<�*=���;6@<7;=)J���%ۼv[Ҽ�������;����-�>�c��<�oF=���;��=V���"+	=�@X�0k8=Zs9=� =����fk/�4�<�3\=���<�S%=�<@b;<G��<	װ�����y�����<<
G=�LN=��@��'O�R�0��ȩ�	s�<�d<�+�::�r=vJ�<ds�d��;��7=T���<��`=����<��<zW
<!0_=�_��+G=}�=B`F<�h=u,�_�2<m�Y��4l��;0<|�W�1���;�}���F�<�k��␇���P�͇�UH=[3ϼ*�3����<�W�Xɼ:`&��7�1oU�ɦ��o����o=1�i��F���l)��<.�<7}�l����[�<���<IM$��g8=%D�<����<T�x=7�E���J�P֖��������<U^j���=�9����<��=08��Ma��q<���;z�p�C�<��żPo:��pj=+Ě<Zd�<������
=���<A1���=2d�<�9P���V�\T<�*=TO�<)w0��=���x"��@a=X��<[/��%5==�<^hZ<�(�<�&U�b������= $U<T���3�È�L��<f\��o������ 컻���>d��� ��Z=V��B%:=P�,�D��T<�<���:��d�o��_}=��"�;�"�!����!<�=w=�Kn<(����u ��2@=:�M=���:��<�=����<I�f��Q�<�|
�5�<�=��.�߼"�%��)$�%��<���%#*=e!��4�<�0�<(�ļՒ�l��S<K$���k�;#�j��bK�����^C^�|o�z뼬0�<HT=S��<�ϻ�c�<y,��@b=<�"=�ּij�9/��<�Zv��=��Q=���9+^=��?=5S==֏V�.o�D�=c�
�͛+<�==��;k;L=�]���2^=��4���ͻX�<
˃=O-=gG=}��Pd=������iP=&����l#��ZJ"��R�2�<x���kT�?rּs_�<]���{=۪=)z���;������<��s�=�Ͷ<W�v</Jo�}�=�"���;U;�������R=��
����	E���[�G�L�h��_� ��,�<��)� |0<q@L�=�׼��c����֙��I=3�'�#��<X��<��6=L�L�&�E����
r���+:u�g=�b<u�2=+6 ��u�<���;���p!<��F=Z;X��oK=�7�1G���j;=��z;�張��$�����9$���	��U4<�9~=y�Ӽ5LI=��8��;إ,=\�=  =,/2�[`I=�� =�h��1�
�`�=r�=�Z=�E<�[ɼ`\�;PMK�����6x�;$�S�j<����T�<(�F;�<�-z���^=T�p9� �ɣ1�4�;?f�<.Z�<�X%��~����r=��+=�~n��&
=�3o��T�<��<t�o<,=<
?<&��[�k�|�ֹ�v(=�%s=�y�;$L�:�;
��=O8�<�:��l�.�<9᡼[�7�5
���<=�`=�O���q<��E��`����T7�����~���'�o:��;V/�k'<�p��<|H?=�!�<f��<�)���w���.�<eѼ��<,��2H��t�:;d=y+�������5=����B�j�(=h�=B=�5�����; �7=�~1<o��<'���e9��/��X-:�<�V��>�<�LT�c�����<��<AId��|�<��˼���ϝ=��?���j��y�<�}���fJ�ͶC�Y���c���'<�r��`�`='��< ���?��?=J[s9!� =^s˼���<�F��9==6?=_�;��<�&��0=�<8[�6�"�����{1=}�ջG#g=��v=�\z=������"��_=�m<l9��=�t<�݄�.D;>���Fd=��A=}�=�3��bټH�w�#�;Pn�="(����T�,�;�'�<��;�z�;	�P�]j)�S�<n�.=��=�>X<4��j�<a +�)T�;���ik���|>��tX��^=�:=���<��<���g���S��:���	�<��Y<Tu:=Ͷ��΃�<�}��{+=\{~=?nb=�7��Ɨ=W$��'Ǽ�N�0������ڻ��=[M�YW�<0K����A,񼩎X�ʝ1=vh�<���ȏ�fk���<�����H=h�=PSp���2=�m�,��<Rޑ�����ȯ�a�k;��=|a=S��<��:<@�
�u�@w�<�V=�����I5=0�G��6�r�=SH��r��%�<*�N=���<�9<��<h���?t�:.�: �<��<��T������x{=����9`�2�=�E4;f4�<���ς-�Vg=�)M���̻���������TA��v�=3=���<�{����=����V=Q'< �e��<����a��Ťh=e���r8�<��g=���<p�I=��:<��'=��'=�B	<��`Iw=P`�;ҡ�;�=��<Y"�
Z���k<�X�:8�;��;�����(=��b��i6=\k�(l:l����_=�x�<+��"��8<fN.�����	�<]�������M=(k=ڧ���y�	66��H��wN���(=r%��,ӻ��W
4�D��m�\�3�<��<��=_sf;��<��Y�_^=U�����9#�<�1̼�d;�o�;�d?=i�1<#��;3��<��F�=�^�/}�<{C�<�2=e��<�w=�݉<a�Ż��A�Fta��0=3;�.�3~;<���<W�;=2������<�K��n����;)?��>	="�b<qQ���!�����J=�B�+aD��;�~)X<�.�;���`S�<��żBSC=J/���*�:24��I9<{s�<{=!�׎<§=j�=���3<�Z:�<f��<�b��W�
<�O�<�=z�e<�H˼\tt���P=�':�w��;��	=Z9�*#�Y����P��!#;�!,����<���<j���5�Xz�<`�_�t��R�������I�&=�LQ<4#9���b=��^=��)=~@�����'���n��ۉ<O���;�wż6�G<�=��9(^7=P�><I�m;G�_=�����r�=�I�g��<���<5���U7���<r��bR/��<���Ҵ���w��[!�M?�<��<U=l�;F`���O=��^=���:K� =���-O=���<��@�6�<L̼ܾ��K|<C8��,��4˼��<�+������������I���E=L�,=�Dɼ!��>�=t�ܼk!�vZ�;�����C��h"��._��W;t}G�( �<m�=��p<�~<�ҥ[�r�s=+��:!�l=(��<��<�2(=�仲j0=��4b=���<�1O<�T�h���仇�<%��4<��kk=�̼��C��[=?��NZ==���<]��r���
>�<�v��Y��sz<��/��~;�X=�� =�|<�[b�ϛ><���<�Թ�<=?���"=�Њ��v=v8�<ܷH=�x��Z=��<�a>=(�=:�3��#�>��<�c���=��=}m=�<���>���\=������t���q�%��<@�=T<
<םe=�9��i�`<�}�<>����\�����j�=P߅<c��](�<�=P=e�=S
D=�z4�CO[�%=JU(�D��<K��I�U2=�x��'=<}�� \=�F��yg=���(�m��ꂼ��<5�)���S����;%t*;�5�\�m��䎼���!>���=��;���<��V=9�I=<zb���2�V��|��xp��>2<��+=��=6tP��Ǽ��k;�"�<d�����2;�Ti��랻4��<�
=�q=Ş�<�<%y=�}�<�R��7S<�X[�����yM�<�P��n4=bf��e<�ֆ�t�F= �=P�8=玵�%�;�7��/��`;�?����o^D��L��&N�b{C��5-�⚞<(=y=�`x=M�+�°0��d_=y���ak=�N<`7�v<9���Y�EC��G��{��C�5D=N�<b =1��<��Ӽ�$=纃�<�<�O���/R=!���:[�˵5=�J=~"L��t4=�I�=��?=�d���g<~@��H;<D�����<FB=t�Y�	Z`=�J���;x��<��<�A�;uҼ�ּ��D��]=�l:8��o:�<� ���ϻm}��@X��^���0|����;�f�tG='�\=I#�Ŭ<: 4�g��<
�*��$�<O�;F�~�ʼ8=��-�Dm=7�+�3Z=�R�<�=��4��7�<�_�ֆ=C��v	�04��~a)��fs=/)����[=Z.c��[%��B��f��^>�x԰<�*:=��&=Mr�<��c�[�<V�;d���KE��N=�/=S-=�컼1j<���;���e/=�G=�)�<Ỳ�^=��p;�j]�ˡ�<�R��<jUλ�=a��%=*������<.�ѻSz*=t��<�h=�OD=;P��#��=b}����)�8�� �<���7$<�K�N���Z�U�P:z�'<���Ԃ<�B?=O%�<�=TЇ=P�`�u� =�
/=�?����;yE?�Cr(=I\B�˔T�J�"�\ޞ���W���t=��=��(=��<�~2;�,A��V����<�Zw;��~=O3�=>�B=�x������M鼔S<=F9�O1�<u�J�0�<G/�<��j=>���f�VFc=�q58�2=�R���<ŗ[=������.��?;d�<=���<��=d@=/=�G=(�
=���<��G�&lX����|v;�����}N���ռ�D.=��=��<T�<W��<�H�2׼H�=s9����<p���H3��8=O�=�>+<�ͼ@E0=d����	����2=�<����Ú�/�8��O�GFF=`�X�_ػ���<�F���<K�2�G��d��۹=3�=ê<V�I<���<Y`3=@��[�2��t��˂"���ṕ�M��B�#�Q=k'L���;�>�?>���<��v�x�N�8�p=�{O=�y�Nh��ؼ� =�����\<=<�F=jzP�ŵ{��={��k�ۼ%��<�l�����1=Pu"��Fc=���ſ��_<����X��V=䴹����<�U���E�+�p����<��'�ѷ�<[�;���3=_w< O������yHR�Dm�<,苽�>a��`l��B;��n;UA0�+�,�up�����G;��X�����Y�;�s���"<vυ���H=��<>�1�p=��*6=>�y<<;�<�ӄ��мA1��F_=���l���_�����Ct.=�P�+�D�^�����<�=���9S)=���ąQ�l�K=�\c<�/=�s$�!e]�G�g�t"��:�/�Ov\���,���=:;�<�
=Ob9��Y��s��P��R=���;ʈ=W���
=	��<T��R����O=]����[=*( �/1=��?�%?_<�L�<�B������rm���Q��e=H��;���9��<���<��p���7=�Dռ��/�f��lY�;�U��[�ٺ]�8=��B���<��P�B &=W��<�&�Ɯ�<,�>��r<Fم=�S;��"v��G���H=�xk��6=`�*��=�w�<~�8=�; o�;���T)�<��S���G=�gK�xO<��p�@�p<����h=
��=nK0=�h#=�g�m#�"f���bb��v��h�<H��4��=��`=��+;3ּ�~�<�Dg<��.<�sļF�켥O�{yv�==���=�0;���<b�ߺ��lh�<��#-�<���<�&�ra�ޥ����f#���,p�;z�<�-f=�e<!Y�a+9�Yk5�	 =�R�o���V<d��(�k�<�û��<=yȯ�?(;�ԩ�g����;��,=����8=�+=r�̼g+=sL=K|Q=u�q����{������<� >�0���=Vf=��������$=�_�<��b=N@��V�F=�AO=�l�@�!=��5�j��<���UK=�i���|=	"f��;��	*B=�t��K*����j��K� �=pv
�p(2��L;h�=�\q����9�����c���0<�s=}8~���
�
<� ����=��n<�:�;�=��d=�c:=g�&�o�:=� <�O==�4D==�+<����v�]�C���L=�d=�<s�
=��G�W�ȹaf=p�<*�<��n;]�����Q=��l�\�4!|;�ڻ~�B�2PZ�Gw=��<��=��O=�����0�/�<
�Ѽrq�\�߻�SK��"�U=;%�<����E����!�)Vt=[����<8��-f�=��<�'�Q�E��o��L�-�<���V�~�%���=h��R8#�|����W<��r=mg�<ڒC��7�;U��<��=:<�<t|�<L����B=�װ�';(L�<�Jļ��=ID�<K��la��#H�<~���\�<�k�<��l{��l�=�PC<�C��'����k�� [���$<���<pӄ��4�L�H=��<�n=!�<���:Ԯ�<�G �f8^=�s���M�O�r����
��BR�8B!�_�<�Ǻ�¨<��v<�!ٻ3k�C\�������F[=�L=��B<.�����<)���5<N�E��Z�+Z�;i�+=(,'=aa��pH�VE��y��;�C����7 =�4�<���:�~<���=6Ļ�}B���=&�g�7E������|�$�<ʕ7��*�����4ļ�����I�T�>=�c<��pK=�?=: L=�߻4>�<�j�n:M� ,���=���~�<>��<q=
����６�ӼF���4M�f�=���$e���D+=����Ɣ97HE��`C;��1��V"����,=���乼���<d*���+�'q=��8<^�<��<�=��ջ�&��!�<�=�o��9�W}���)I=P�={=�)�� ����>=����pY=4U)=�h�<��<�Cs<u��<a��I���C�<�V=B�^��y��:=ſa�H@=��K=�Z�9�)=j�-�-��Dn=���]"l�A�<%|�����|�=F�A<�u��
��<N�l���"�S�6��U��?�;s(��l�<�o���鼘��=�c�帽<B.�<Z^�<g�뼕�4�>�ؼ=��<=dsS<r5�;!<=*8=�!�<�؈9b ��ʼ���dp�:��.c��N��=�<�=��o�Ƀ=7v�:��<Aub=�;񨼒X�;.��V�G�A��9W:=x$$�G�[=@���3�ɼ�s��)�<P׼���<��H=.�w<&O4=hȵ<�����<@�=�4�<��;/=O�==��<n����<���Z�B�^<7�9=T5&<��=g�<S�\��
�4E���O='���z<{�)= +����:� �<Gu��Or���'��=#����L��q�<j��;x��;A�&=�1(=�`=�)=	/<n�_=��<w)=Ѽ���9V�=�a�����<;7����8�4I<��������¹;�D����%���bS<�};<�#��P0���=�c�<� b�׸��Τ�	��u=��T=�KT<^U=��7��D���R�8<�}�<�	;�d��G�꼾��F�;#��QCU;x��:$I"=�3�;xUټz�5��.~;Ed:����� ��`�;(A%<�[ԼeXL����*<mi�;��j<U5K=d��<��t=�n =�X�;,щ;E� �-@O��!�9��Z=Â=�ދ<H1��w�<�;���F�<��<�X�<~�<e[$�G�i=|��� =k���6�<��!��a��z���&�?=��=W�����<J9�R�"=}�p=d��;)==�M�<)L�0�� �=���'��)U���a=�p�:�¼�鼮q�<���<Pa����<XL�<�9�:�<���������=#�<E����!L��}�;����h���*J�<@u�<B�M<Z��<����-=)r��A������<�a<�3=�W0���=l@��,�9&/Ѽ��D<��ؼ�2�.67��]��W��;4����?���S=�1#=�Fɼ��P�D�`����<�#�X\���^t�<��?=���<�����<Qo缢�<��E�;��<��x<D�L;���99�(<8j'��u<~�;�1=ۆ'���7�������3k�kv�<Ԫ<ӏ��"p�i�9=��+�b�F=� ���v��a=�X�j��<:���0�cq=?������|x<v�o<cmX=�7d<1:���=�����<�4P=��.=���<K_[���<%Q*<�)=�~=�?�(�B���	�Ka�<^�b=qYڼ���<��ؼ��\<��!<���;�C)=G�0=Z����}�<R�m��Z9���=7Ｍ�f�R�	���j�=c���.S<S#��V	k=lX��y4=F�N<�ټ<?�9=�7�<&9x<��U=\����(�S.L=��U=~v<	r���hܹ�I�<V��S��2�����\�j$��ѻ<�s���<����'$�<ؙ�����<L���ĝ����q/�=��`���&�d�Y=7�k<�H=fNE<��=> G���`�˯q��Ւ�X�p:��7�=����)��=��l�9�;��T� ��<��y=���<"Bk���uD价��<v�=g�伴Ƣ=�N���,�<�g�I��r�*��dP�G伄��������j����<��;n�:=1'F=j�&=ބ =с3���'9����<�;��G��˖<�U,=�.�ٱ�<�ή<��O=*D =�6�<��B��q�<	w=�]�<,� ���<Ͱ���><)��h�&��[��,��z�Q��F�m�
=@-���R��� <+V�<���;Yv�9�B�&p�39��3R=O�B�4�B=R?]�V�4=jS9���;���Bd�4aF=,���2'=}N�;�s=Ϸ/=�Q=�A���E=�JU�`f�<��+=O�<|ż�R�<x=�	h�ڒ=f����<���<NI0<��;Q���S��;$U����<|?4<�I�=G��<1�������)=͸l���e==�ƻu2ﺇ�N=N�6=�Ö����;*�<_0o=�4R<��e�u��<�I��<�_>=j3=ܕ<=��	��"7=7�<���?=�ƺog�����<�<pAc=,��pX�;��;�^=���'=z=y9�ĩL��F��+��E��$�<Z�6=κ`�g�<MnR���м=����<� ������2�Q=;��<�*o��s�� ��<��!�n@��@Q=��l=��z<��t=W���ѻ,(<G�<���<��Q�S+�\?=�e�;@�F���<�?��E��)Y<ٽ,<,�<�~C�d21��^��TS���N�4��<P=�F+�C���@����缬�3;"��<�a��ƼN<�.���a��,���=�~r����;;4�<;���� =�x
�,��<��<�Nؼ#�V�<��I*<嚅<̢��2U<�U(��	�<bj�S��Y����2���<@G-=;<<=i��� ��h?=or=܇<5D��cl�Ғ=���.����;+�ƼB5�;�=K�=�;���+=n9�<�B+=
i�;;�<	���Yһs��;n�-���I='�=ya,�%T�2����^=�oR;��=��7��{m�7鋽�~�<^S=w^+�K>�:�t<��X<�8��bL]�)�@����< =*6_<��s<�q6�F��<ԭ�<��$��
 =*Ub=I���+~=y�������K=� =ϚD����~�U�b��rz=��<_�@���G��k�<�c�<�]h<��,��GM�QO��O� <7'����PFY=�_ ��,�u�6=�F��;�=�L�<sX�� xo�Zj�<q�=�x"�����h-k�Uλ��B�䎠�	8�<�+%��y=+�<7���gr�=�P��iC����}�<#����B˼�EU=`I��<�=ļqeV=�2��E=��޼�Zp��|W<!~5;fN<�ҵ�j��<�V=���:4"Ӽ�='��<<8��¼>�<�����W;M7�<tC=4�K��9=ule=�]=�G=��<<5ټ��W<�	=6Y#=�Y�/��m���0�\��a�o��<2]=��=2¢;��a<�P =�c7=���<ŇD=�;�πU=U3	����;*@�<�m@�	1�;V��:&m9��-��0�<"!�'F(=��<���<G��>I��R�O�n���o��(��<n�<�M��T=�==�?=����7��FJ<~z߼�0���m��9�<�A��K������f�ݏ�I��`{=����mټ젉��<�+�'���<'n=B�a�$� ;�������v=���5=���;!����|Y��Ƕ����<{�+���5�En�=YI�2�H��S��E��W����f;�s@<ᬠ��@J�P�-���<m��<��=�q�<�o���!����;�E�<���<]<��>=}��.�<M�>��d�$ڼ6�U�}/><�ﹼ .��׌���y�m�"�[-<�R.��k0=q t��/-�y�|<�c�����a�r=�Ic=qwy9m�:�ϼ��<�	��2=�혼N˼�<��K���1���<������;�_c=�x~����ޚ=�`ϼ�	�<)C0=�g�=Zҁ:E�����_��(�<�1.����<�)B<y���,�~�)=HQF��f�<Mtd�D=`��<�%�<
�1�;eq=<�4=H�f=��1���<�	t3���<��=lZٻ)�Y;\nf�d��<o�8=�� ��_G�KnD��k�UO��w�W=_u<nW<��<��5=A]�:B�������E�o"�<t� =�����<��\<��<͹%���޻ch(��r���;)m������%�;f O=G�#�?xQ�W���R�u�%=
��<�{<=2��@�r�F����<�?=5�(�V�<��ûć�e��-����b;k��a��<(U"��e;=�G����w�l��<4w��Ȍ�2$;k�]=\c"��PU=lM�;��<���u�<C�\�c��������L<�G���О�����E;=�>�<"���-�F=�hQ���F�U�8��~u=,m<[*������:��}!<l&=|�Ѽߌ��S|D���Vp=�U�<qFi��� �A�Z<
) �!꼟���˟�=��U<��Z��N��B6=��M=Ԉں�/�=ZF
��nż.%�Uv���v�h,V=+��<F��<��=���<>@���d��%o��y =��O�Y=d�ռR=7�3�pp���?=�<|���=�K=Wq�<U
=�ܖ��+��|>H8����=����=���;S(�}4��׭��l8=��:�M�;�^��<=���� b��I�<$UϼP�F=�R=Ǵ��0I=}�=zd��q��1�<ɍ����Q=vb���M<���<
i�<v�"=k|,=ʅ��4���ɻ�x��k?���B+=�u�Xa��r�;RK�=s'�<�Q��<�������<��/;��<N��p�^�i��2E\�
:�<�<=�.����3�<�Y?=ɝ|��[�<Ԝؼ����O�<�o=���:��S�`�-=��B=L�O��el���-=�q$�m����@=�0<r�����<��=� ��f=6<7��r�<��l�q_=���<j>��<�g�;t�;@ZA<{s!��ɼ<d;�;Z�������=v�yx�<�#=e�<�O��zX=�Ba�)n=����_�2���A=$�(<��</j������j���<*�I�)=T�=�Eg�ޒ^<3�1�F���C��5^K=��=¡��ʜ;[�8=�ŏ;�q=uab;^��;����XBy�bQ�;��<�]B=�<36;^��N�<F�,=��S�0az�^='#�<4��<u[/=��=���f�7�f-$=�^��(��<!��<��@� �<z(�<�0_=[g��hI��-�<��<�CZ=d==�|\=e
�<+�T=D_�<�R�:C�c��p绶�3�D�w<Ye�<��<�FR��K=U��yni��\��?f��e�>�	�`M�<�W޺��y���=nZ.=Rcܻ�|��
[m=��<�)��;Bk�<ZZ�A��;�#�=���1$=��Q�4f�< �ϼ�����8N=/D���N=r�Q��B����K=l@u<��ܼ��=<�<,�z=U�q�u2=����<4I��<7.��q���/��*
���L�
E9� �;���n�S���;��!-<Ue�<f�<,I�<��<?�e=�%��!Z��qg���7��Ca�WQ�<7��<��$������Hf����MUw=�7�<�D��<t�Z|μ:l�<
��<	�S��m��ۓ:�<�#	�<�<��c����d=#=��C�	�8�/�<7w%�n��<��Y�W^�ܢ���<An�I{%����;6k=%�(�e�G;N"=�����E6<8F�<�MW=�F=�/�<�>3=���<�`=��
=�W���S���<=�hH�4M^���<�*,<2kV�v���RV%=��_����#q<t6���%=a.�R���&�*w � ����<@��<
yw��P7=�r=o%>=T�;8�/������%����%�j�=^r��4���&����M=�������Q�<�����8=G_s����<�/�<Ua��b+�L�Ի/v[��(=V(��ui�ƅI�-�q=��4<�"N�bS�/iW=��<�������i�M�d��<�p�W�	�b<`>�����=w4�;�R<�뮁�Ҿ�<5�5�;�y<��F�C�n=
(7�t=��P=��<�m��<�3b=wk;<x��<+��<���N�ڼ�|�<�<<�,=�����F=$�����O�i��ܧ
=�1��3$=Ѕm�����<i=�iO=mYӼ���:��<�1=�I�!�J�j�j�p�s=��/:���< :�<��1<
Nӻ�м>g7=�P��F�SK�j��[߻ Z�?l=f(Q=X��5i��)=�li��|[�8�W���=�Lj�42��_!�;����=�-=d⻞�P<��;:�$=I��<mLE=��+��=�*��}&�;�+��m�;��6=�&��}��<<�ʼ�<Q�'��k��qB�@/g�Kx�< �=�a�<i��|g};ղ]=�= �K���a��o���j=h�i=�-t� `�.==3�;��i
��-��=m�)���$�Ye��̘�9Yz<���<+E?�r=�����N=� мs=B�:9C>���^=�,�<W\|<(���`��v=Sݼ�p<�X��Θ��Ἓ�N=F=łL���;�U<̲����_�$����&.<�H�<�=b[<o�<�VԼ�J=�b3��N=��<�C=0�<s/�<~�<gμ)�^=���1 �Ñ�<�2�<�!�ӑ��F=k=��=:��;�u�{�g��<��4��}�<����-�<�Ze�馠<�`<lR=���:!�h=��[=���`�l<�N�����<�)=Z�(<jݦ<�4>=�-�[��;f�<|�Ѽ^��~f;Zɼ�=9ml=�o�<��� ���K=0sZ��9����<x=bG=Ӑ�<s�;���:/��)5B���8=���>���gໝϼ��6=`��<���������=4�"���"� ������:�:C=��K=	�=pE���#����;��=/�s�}�o�z0��U<���%�!t�<���;5�=�6C=Y?�Y�nN!=r.;<	02�W6�<��{����8\=z��l6=�<���!=����4����yZl;+��ġ�<<3!�;�3<Ȁ:�dS��lj�L�K�uzN=ɒT���3n�AQ�<W�=�Wb�h�>�_�ݼ%�G=��;��	�<I'/=�;�1�<��vt<^�;��(=�Z�<�Ӽ.��<J��<L�=� =�~M����;k��<���:�	źg�R=��лz�<����;8=�=�r��=���<��@�x3c��nܹ�7m��l�<R�!=na�<�F�<���<��B�n�j�Һ��eՎ�=m�
�5�yR�o�}����=0a=��=D ���'�t��)�.���(=$f\=��r=�F=��N� ��=�I����<��Z<�;�cּMW�u�D=���;bl�:�ꝼ
�<�<��4�����y�;���H�i=o,�<,����`(���<6)�<���Β�A�M�z<�bټ�-<�l-=%�(=!W��C�0=��K�'7�ˎ(�U�!=͙@�s˻����9���+��݇=n� =��Ƽ|�!�%?<z�5�gp=;��ݘ	=�1��4 ��T�<���}�=ua��=fY��>��A�=�k=�V�<�
�<��=�*�=qM=��M<bU=�<��<[TJ��x0==�;�p����{=L��:�ܻ��u� Vl=��=lC��I�<�J=(��od=�T)����
x�<���<���<�0�;4���mpd��pz��aG��9�&Uk=5.T��f�<��(��貼J���
�J=9��rF�<H�<{��<V6*=6K#=?R <�?^<O�>ּ��2=��=���|��<6��<����)�O����<�
L�_ܠ��>'��%�<7�Q={9�[�=`6=��=����9�<TQ='��<�V��KF��?\�¼i��֋=��<=�I�O��\t���7=����p�<�0=/�f��Ο�==���;^�v=�KA=3j=H�=�^ <�'��3,<�����<��{=Gag�	}4���	��E�:u��/8���
�ii<����]6���R��<.=j9"=h��<�ݼ��5���<r�/w
�X��a6��#=�EB��=E��<}^H�V���@�<�-U<Xp��W�A=�u1�������; ���m�(:�ܧ<~��S�<7Im=��p���/=�=%����j��|g��e<ϭ�:�F=)�<�3��@?���n����P:,=<��a�����;Bb�<��[<ۙ2�z�ż�ڲ���;�~>=yo��cc�ik¼=��<�="=};�#��=!Q=��3���<=�k;�Aw��<4=��f��9J���z.,��L�:��b=��⻜Xx�I�<�!q���:=j����d]�;��2�g��ԫ=vi�<�����fL�ig:=�.2=d�N��H����)=g�*=E�:=��S=���<4��<L��<Ȑ$=#�<gc�<y�]��<��Z�zb!���A����<��h=�3=��F��=�`s<FF��=Mw0={0=�@��#@D=��j�Q_������;4})�C���3H=�7мm��� �5���<�8>4��O�<+���k�Q=��$���;��=б#�ٌh;/�f��b�<8�=��b���<Z��<��Q���r�?k=Iw���<�G3�+
��J1�m����-=�B&�%2��Jb=�����mo=S5��/��<j�c=���<�����6%��-�<�~�� c���7,���[��[=u�"=�7=��8�cT7=͸=��><��<6$=�U�΍z�1j���:�_P=��l=|�c<}W��{�<Vc�H#j=�2o�g��<W*����.<�tм8�E�ɛ����<��8�
YV���W�K2�<��2���<2A�<��'��jD<��3<�Ew=����W�f=�n�<��+=]j��^Gs=580��G���|ӺSG���KN���F=��7��{=X!L<eS�tt�m��}�H=:�o���H=8SF=�$�;��;V`<�]9<o�E��V�<?��,�,=�m=����{䊼ě7<��#���¼�y�;�Q=�<(�<v�4=�=�<I��<�»�OO�C:;Ж���q�<��o�V��o��<�}��O�=�ĳ��v�	�D<>�b=AW��hc�nVZ� �]<��!�:��uh�<�fżrm�:�３��<=�=8O	��7��؂=��d����.�0<� ���=8g����7�{�=���<�A=6n.=K��<ڪg<��o�بk<��׻�Ml��E���J�/��+��I��!���U<�8�s��<��=�? �w��>�=C�( S���H=�Y3��ڊ;���<U*=�5
�L�A=�0�:pL?<���<0��<�K��A��n����;��k<M�J�}J�_�\=�0ӻ��<�F�+.�;��L�<g<�#	�C�������H=i5<�T$�'�7�����J<�1��ܙ<C F=؊���g�� �=��p=ۉ�~�)=ق�:���i=ZD��JV=s�O=� *��(�<�M�<F%<�l����;§��N��o�u=_�m��C���RE���	=�tY�� ��<��#/�<!1��3p������$��I�<߈��_iD�w&�<��C���J�F??=���<��{<��< PM��y�k�<�R=�p������6��m�=j��;E�=n�=<I��<�e=).�<�B���A=VQ����<��
=� m�	�����:w�x9xd�<*=�@?<�xE=�<=��弤x�<�a=��Q�R]9�2A�<�~�<�U0<g%���.=#du=E#ü��a<:.<��7<�޺<�	�<�"ͻ�1�O=5!!�
;�<FE
�.'�.����Y,���Uq��(7���Nڼ�����`(��s��_#="=_V�l�2<��*:������J=��9�],=O�T��(=*�=T���3��A9=���:<J�<|�<�"�<�G<qX<�>�=��<��7�cg=����0<t!�=3t;�`�������7<8��a�$��dL�[�j;��/�==,�<�ǣ�,�>=cI=�=�|E��F�;!���a��=_=�+=��)��.="/<L�<ؓ��T�<�p=;ԡO�ԇ��SC�ʧ�<߀��������S�_���B<V��:ArＹ�M�<$nM<�m7��d:��D=xĺ<�&l�@Mn;w<��������4=�~Ӽj�_��<�׼k;I=��9=�8=��G<W*&=�_=p�f�)Qb<��<9��+
�0���0=|>�=�<�<>�X�=R�/=x�f�̤��
��n�?��G�[<�.J=E^�a��:��;�q=�\�=;�����y��bt=9={�f���8=O� <fO!��3���Pi���/<1��;ћ:=����̒�?끼S�<3H<���<�[��x�m�������/z<���<1�t���U��F�4:g��M=���<X�J�l���
3=��}<����*{m<׉6;�W���==����#�՚�<��1=��=�<b����<�k��-5�3/��+e)�W���61��=LM���:I��;F�i��Y/=UWn<�
)=s5l=-�=�iO�!�׼'`=��+�c�-��Y��0�<Xb^�s��<��<	(�@Լ��=���<r�%=k��<�=O�F�[�����y=srM�h4;e��;r4��=$=��,���A� �=�vS=B���Ѽ�ݵ��f�<U���X�J�$�l]����_��M�����_�<�{+=,B,��om��䡼~����L���h,'=��Ǽ�)���3�<J3����<�2[=�o1=�%K���Q�OE=�ì�rм��q��lK<��7���8=��<��7=]�k<U��s��A
�� �8�P�=j�K�3�M1=��s<�%*=�Wh<g �<�P��p|<xjH=�1��`��7�<�����<HD�<�����<��%��a=����=����^=f�$�X�=[F&�Q���d���s=��$�g�k:�(J��_�<��A���N�Gg(� ��<�79�u�<$�B�E��;��.=ǐ=�@q�<��Ѽ*�\��x:�u<j�:ֆ;�4�;�F=�Q��N�=�z�J#t���;=
q<�|Ǉ=o���#E<^N=�? �i�<�1�<-E�<ŋ�;��l��Լ��Y�e*=��x�F�<x�t�N�l:��: 	=�҅���;�	��h[v=z�A=h!*��=�+�;�b:T�����%%=�:⼀�<�N�v�v<P`���݊<�]2=3qǼ��X<�M~<Vü�G=�u���Z�;��!=�H���ջ0�S�/�x�ż��<�Dc�<�=������5=	���Ҽl؀��D�<;��<��$����B:��#�<�z=2b;��:7t<�8=�Z�<R0�z�(�0��l��%�&=F��<��d=K>��엽��%�����,��<�4�<y�Y=��a=t�ڼ�^O<�Rɼ�;&�f��t�<���<���<�ʓ�Ŗ��k�;Z�"<$]�<s�i�̻�,F��?}��+d��8�;$E��bO�<�F1����k�<�c=��(<��;�l���P:@����,�wc�;���<f�伛6<�A�L���C<��ԼӍ�<r��<ݻ=p$!=�,<�U�<i K=1:j�we=��!����<�xf<��X=�K���8�9�l�;�ܼ��=��Y�������퐺�����N�50$<3<G�D{O=���<\��o��+a���@=G��<�>E=��G���d���<�%�\Ai��U��ι�<bc�<�m6<N<�'�;{�˺�<L�߼`ց�Â��U������G��m=��?���;������;���<L̀��02���:�*��g<KÎ<�AD=��<r��<�~ϼ�M�L?<�?>�aJ=�@�97�;#F=��:�O<=��ļz��<��f��l<f��<���=ĭ@=��r=�=�<�`��7�^�=8hg=*	������8	��7<a��<(Z�=��2��ƶ;3�<r�.=u���o(�;����g=7���8��C�<�K��R�8��<�s<r�r�ڰü�Þ:��&=(5�=�^;2Z=�m= ������<�'�<_�0=�
=�Xg�k�N��(�[˳;��Q�S�;�����C:G��<, =�":��w=��}�gb�s�w�_����B<L>�</��?ť��ҩ�I!=���<�]=^-L=\8���;��s��s�;�Ym���=�#V�<N�(<���<;�	9���x�<6����.�;��"=Q��<.ּ��@<��n=-� ��iv��SN=J�����(���<���<�j�<�N
��*=��A=؋��;�=o�F���	�+�?-�h�z���^�k��NpZ=�0��K6=k�+�:��<�|����I���V;��,���ͻ!
<�E���D=hrüu;<
*d;N��=$����,���w!��`��޵��/8�;��N=B W=;�$=D��<�����:��4�<!��r�#=m�&=��	�|���Ի����@����M�by�9�;��U=��*=�*^:���<c����<.�C=�J�<�p=���:����\<(6�wQ���ͷ��,o=d\�|`�<x�ເ�(������+�;�Q�2��=z�K=�u=-�n��C=�wj=�tz���G��N�<�=6<Q���}P<ɸ&��6�<�D�<W =a=GJ�<���H�=H�7=qd������=��<՗(=��<��<�V~=��<��S<�i����
�����k�r��ca=�WY=D�W��d=ɕ�<tA=5=�Un�kD�;n�'�{a=`w\=Cu��m�<�B�<�2=��<�lU�<������C�|�ż�Q��@���C��6E<9��<�`=�%����������� F���I�:9�<�&M�����}&"=ͷ=!;�J�Q=��Q�X>�9�*=�a��:�ټ�ᄻ"<�<�O�<� Z��`=�5<��==zH\=��3=lH =�L�ٶ;Udi=	zں6�=�А�wo-��w�;��.=��4��݁����-uH=jI���O=��)���<�=.=s�ʻG_��jh?��S� =&�=LhB������x;=����Jּc���<:Q�;�G!<�m<��*=�A=ڗ�;��t�㢂��1=_Fs=2�;O}3�ZSJ<ٽ=��Ai�G	-<�$d�ű.<�;]�$N����]�������y<M�X����BQ�-�̼�!=ƴ�(zP=H{<3�8B7�;�~R�P����A<_@缲������^�<�v<^�i=.}I��~�</C�=�(=����0ļ��;�I=�!��1���:�\�D��<^���p<�J�P��<��G�d����j�P.1='>�������9e�P��s,��ɺE�M�T�Ƽo�l��M=h;��W=B��:�1μf�=�X���=p0i<ș=�w���!��[��Ca=��T<kV=m/��ug=���������>}�=���<��&=�gS��J�<g�W�����
��Z�=�
.=C=�=��<�7��B=-{���;�{Z=+�<7���2�<.�<���;�m�<y��<L�X��5#=e���j�7�dV���ܼ�D>;Ni0�O'�<�L1���4=i)B<��m�_��w�0���=�ฺs�=�nL��	k��g;�ǝ��ּs=y�v��0�<�sA�!��%8+=��|��Ri=�0�0=��9���>���T�Yu^=Y��<�=+�^=`:#�A�<���<��&�O�e���<e<�=�H��Tj�; Ǻ<���A�¼�5=��n=X������p<��=VX��rE�,��ǏԻؓ2=� -�=
�W(�<{��"�E��-=G��;����:�x�h�0I�<2�,=LR�Cow=�м��뻓���n=��<�;�=R �;d�8�ޯ{=�Gm=� ��xK=if\���1<�E=��/O=����B'=`�\=�D�<�D��<�﷼�A=�H=��<a<��R=3D>���<Fڣ�	m!�Qcür�t=�(�H�Ѽq����k)<�;�2P� ֕�|��<hG=�=��;���=a96;�2m=���=]�:=�A�5����\i�:����M{=T�]<�wx�FO����<��D�#e<��D�8Vm��IĻgK=����rm=�����s�<�����<�X�<��<�?=��A��U���8�<��u<�����=Uj�:e5��=�=��f=H�f=��I<�:.��Y=?���n�,�;=lN�<����M��3���}f<�k^�B���ژ�;���(�<}�<=�$=pF�<���rJQ=H�<�(B<��+�~�<���<�h�K�<����<�f�;���;Mc2=�c�<m�K<W=�7�� <&�A=t����:m(�A"<� I�W�,�}\t=������I�Ðl=fF�<:�8=*X=z$	���#����;��=Jp=(#ú�l� � �ھ�<`:�<�Y����6�TN�;K��;v	�G�	���ɼa*��� ������/D�֠/��=���<�ȧ� ��<�#=F�
=�i^�L��;���W�+<ϲ�9�W���<{�,����<t�J��:=ī��sK=d2�<Oi�ҰO=bE+=7Z�����Z0=i� =Z-�<����(�X2J��p=�0�U�0��[�<?�=�\K�������8׾�EK;������<Җ�<��
=w��;Yu�<���A#��r�<F�p=�Ȝ� ���J\,;&ݚ����*= N:={�{;r_ۻ�s&������0=d�.��q=;��<r�$�7�=ȅ��ָ��`�<�♹��i�Ҕ�ԣ�<	L,��9$���%=z�z��V=*������,�)�:����=̾+;��<W��<��
�}�|��X=}�|;·�<0���z�<gٺ�HA�pG<�k��/�<V�@���P��B`=v���׻qpw<�Q����J��<V����\<��ռ�Z%�j߻Jܼ��7�+;�[U�=�<��&<1Ǽ��7�YU+�
�j��a��<�@�<�h=.B�<*�<�a���]�������/� <�E���w�;��(h���;�9= �I=�r�� �d=>"��ZZN���=����7�=W�c=�J���=��=d闼dW7=��z��"�b��<�6�<b�T=�(��o��B�M�;ˆ�<�҂�OFg�|�!�'P�<A���Px�Tv7�l$=.2�;�낼Sռ�N=��;�XZ���<��N;�4��)�=�u���;=}K��%qu=a��<��S<J3�ː==ԩ�;�j=Y�C<~�;=e�Q=2Ӽ�Z���E0=��)��-��/��t���9�M�<� D=D*��H�8zBH=}�<7=�<����A?=u<��N�;�P����;=�J��E�R�3�G<碻�_z=�i=������%�)_;%g��<3=�h)�u��;�>=/9!��1�<�Tz==���8�)Ѽm|;@�=aK;�T�,���q=[�<�+�<�8�U�T=}w��Ec���Ӽ1O�{�==C��JP���5�����<e��<HQȸ��¼���:+q�I)��^�<����J�J���z�-< �=�G ;��:�l>�&˻��(��Q�;�c��Gʼ�I����-t��C7=3�]��`��%l�<��2<�1F�����]�<��>���=�T-�����L�2�`���S���j=��;�c:��/;0�%=qC�=⥠<�/��_�8����s-=	@�<)7"�h�=i�D�M�q��Δ���<��	��x;/��<Ώ<G
G��F!���P=�����<�Q��h=���PT�<��Q���M�Z����<}�O=���	�;=j�<^ۻ��Y���}=N�5�&�6=3vM=:��,=�����9߼g�=S��Y0��0κ��3=��^�^��R�o��I��]C��Ǽ`�E�U�K<F���N6=�PK=K� ������8.�;2�==&C����R�7t�;"��<��ػTy��<[[��⩼5�e=*�Q�8�w=;���=��ȼ`Ƽ�ų<�<Y=ѡ;o���bS=푻ج=m�'=>�l<2@x��5="�H=�; ���=$��%gG;�p�{�.�A���ʽ�J�9�a_=%�<���9�)��%�������q=�YP=�!E���R=�U/��\�=��=�_��:�E=L*��m=+W=�=s����E=V+�=ԙ<wJ(=<һ���<��~�����d�D��ĉ=/���bü�;<,�.�A?��ci<�H=mD=��X;U=��"Hr�Ix��x��<�'=2��<�O9���=>"p=J�<��& ��<�J��m�A	��h�Q� �^w�:�}N=a�Ǻ��3�3K�:��/�����M=\�˼��5���E�N�[L =����'w1�J~Y���J=�=/�>=7YA=�0=ˊ�u�`=�~=8�%;��b=�,}�	�����=eMi��c����k�=4�;�"�3|!���A<	�<�_I<�����49�h"���''��<�u�;H��<�����E=H�-�q|^<��o=.�<��=�@<����<�T�<L3���J<�
�Zd��vU��K�<i���F���=6�^�5#:�GB��wռ��=�=���=��`=�T��q\�#hW���<��^=�V�<�|7�Ҧs<֞<.�X<�`�T$<�;q��-��+��7��<bz	���[��s9�UE��b�<`�=����zT���=;����϶��/�-=d.=/GG=��Ҽ[� =`����db���2��	6=ɝ9=a'8�| �<�V2=��=�W;�и�=B�<�R_<k�W=7%=W�/=$��:[N��g3�<_p#=�`<�A0��<.=�a?�2�=`ݲ�`�Y��,&�� <w�;���,=�)�4��;�ͬ��6��μ�����B���3E�<'� �-�@=Q�S=�=��/<�<���Pa�,�_��< �-��L��60���u@=	�^=�y�=�pj�K2w��-=��<�9мߓ���=�<���bx�`u��7<�d=9�;~wx<f�=�<e�<�2=��.=/
F�M.;�=�9�<���<�=�n�<���<�@=�RY���)���<C��<_� �8.O�RTͼ^�Ѽ򃺼���;;�L��\[��!=��ż~00=��7=�����X�=��x�<���<+'.�8 =Z�$=�>�˂�<��G�?9=�E?���>\�����w���%����<=�'=��>��ڼ~�������#�<M��<��S��c�<l�@��⾼n�b���5���;���;U�3=�C�:��;N����j�i�!��T=eʀ�����<P0���<�=~���-ʼ�6��b=�A��.3�Ո;�:�<U�=�|��켈9V�_A�<ak"�]�O���X��'~<��/=��=�/�<߿N=�ꗻ���:w&�Z�=��Ǽ���/�<�Gd��
ʼ�	=n�����A�+F���< �<J��:�/2�G��=������ļ��Y����!=�v���[�=Ϧ�<LB�;�]̼q�J=�[*<�*<�~"=��Ѭ�<�S(��w��z/=a8��������ڤi���=��F��/�<&Q9=o�:bh=���<	$P�)����O9=�w�U�,�N2=J�<��?_z�a��*="��'ʼ�D/=XJ=¼��A=�����Y��R�;�`x<��U/[�l3,������<'t;I���]���+g=��M�(<�< ����^V<5� =h�?���!;j��^~�n�a�f��<��<�59�[�<N��<ɝ��D��� �q=��*=����P<=Y��<���<�n���|�;
=C=o߼�y�@
���;� ���<�ER����<
bƻ���<T[��t�+<��P���ļ��<���	\=_&o���$���:�)"��n.<���v���<�ԉ��:@=`���]�	��J���h�r�d�zX�;y:U=e
'�n�V=�9�.�h�R� ���<(�<4��X�=���<a滓kG�M]l=�Zۻ�b���;�/G=+ =Q<��R�>=D:���8I=��*=�D��?�<��*=�p=��"=��缬�'�xƱ<ECG���R��Q2� N<�n=H�<I�!=��=[B=��;<v#H��w�� �<��<:�J;�ܼ��;�Ӑ�<���=pN�H=��E��cN�=HK��>�<����e�<�gʼ�|�*��<1��i�.� �=���=�nX�&�<Ҷ�<A5м��q=#9� ;4�;�-���&=�z��K��y��܂<��<���Tb=�X%<}�N<f�<�`_�p1��}@���<��g��W�<֑�����=�΋��N(<']S���Ӽ�AV�n��;\:�;����<֓5=���<^�<���: |���T-�攻��?=5�]9 `3�U�}�Ze=%�=b�<`b��Hh���<�+=�E�<"�;���<g�9����;�퀽{S�@m׼�I���Qh�P
<�6��'�:b�o=v�<�N=��.<b:���f=,���׼�@-<pM�軁<'��P�ܻ�f>=
z�(�= >��83���$=s�S���ճ;*���R�(��;��<08%<K76=��-=Z'��t=	{`=����T=]����f�=��<�̺<��$�D�Z�M�/<	ex<깆�	]*=�Ñ=[}R�4�2<�T��W'�<BMb<�RJ���D=i��Ɋ�,h=�G�<
��aR<��V<�]�<��"=�&�s�Z=
!x� �<�u�<��Z �?��;9�u<��=~N�<|�=���<��<���ʄ<*�^=<�|=���,�<#e�<�_6;?�R=��x�L�%��;�J=K�"�@���6�b4=
=<� ��q
-�����;��:=/2��L���R���xȼ�w�<�j]�(�<)���ϧ<��=�f����D�Q�Q�J��@�[��I<͡�;�Xj<X�N��A��4(<"�=������<��z�=��7=�M����<g'� .X<�E�<]H��K=�y���û��=��c=�_u���=�%�|������a��mn��uu�:(�:S���+s<��C=�T��v�jA�,3[=տ@���;��<���<?%&�iM
=j�Ȼ��r=�{����=E��<�b=�F=�h�;�A+��!�<��	<"�=����;	��F ��C��:C=�=�"ټw݊<�v0=qG5�B;6��-�<��=k�	��<�<�	мi��<X�ȼ�|<����e\=��Cc �6�}<�AF=4R[����dR����޼�M�|�1=�,��q��<.�u=;�	Z�<�1=��2=��[��>=�G�:պ2=	�;��:bbc=�E�s�;B��<8�g=�Y4�s��0kq�1�z��~F=��ټ�2����?I�<�3%�O]f��n���!�b�%e=�q׼s��j�_�_I|�Ǻ���K�A=�?>;�V=��5=O]�=Ժ��Mм��<�R<��R=0��<_�|� ��<t��{���`�-*p<9U~��_� b��cּ�I=�5B;Sx=��<��8���<�>^=��6='���}������<A>;���;FR�U�V��������<�Q0=�y3<�4=�u=[�:�OR�J�W�J�3|��qFB��OۼfT��<]!2�%�<�|����<E�m=�G#�QZ={m<C
��G�N=�r߼�.$����B�=��I<<�-����b5�0��<G�*<��
=�O=����7���<c�[<c! =
�F��'E=pc�<)�%��n��M&�<=�U+=�� <AaO=��Ǽ�t�==_<��a�	��9>�<G��=^b=w%���X˼>�,=���:���:>3.��%=� B��T^;�R����g��^l�X =��=뀇��M˼ ?$=0�=w�
;�Y=۽.;6�6=֬F��r�<��?LQ��f=`ڼ�r�<�A="�C��O��/i��N�<�1n���>=$�<6�j���(����<̌{�O�<=N��
_N��Sc�&�b=��<
D=�󄼃G������0I=��$�
��<���ށ<P�:=�r�<͘ؼ��=�)���Ђ<Ԉ����Q���T<�M�<�VM�N�����d;�]�'W��=��n��xD��3=f�6=��_�N�8=�ӈ=��F���=C6=� ��)T�:�N���#<�N �!v�<�S0�fZκ
n�[�o�ݰ�<=l�:�@J�=!����"����<8�<�R��x{ = =I1=B�<x��G<��n��)!�|��;�<>;��<��-��	0���J�&�<= ���o�3�b���.��Qw���<�_G���U=�h�� �B=Ou=1�=���W�	=�*=����{�6bμ3�r�l���B<ۦ�;_,<���_O��@��/'�<qT=U����z��=���<W��	�<B*��1�^<`�\=�d*�`��l*�<��h=l�Y=�F=�m=��� <�N%��Y#���:�7�;��n�c��Ť<kJ
=�+t�9��!:��T�׼��<�<�f-�Ր¼|_ =H��;�u���m =.�6=`���}�<wqi=:	Ȼt!2�LWҼ��<)<� ��L�:<���<M�ȼJ�X=�6=�q�=L�<V�-=���#�<ўe�X|=�9��S�<�u��i�$�{�2uͼr1����ݼ�t,��Oݺ�h����8=������0<��T�Y��<���<q��<�@��3m=�@Ǽ�<b���.9���G��V���К><�={�e=mH��B=���;<
üр=�@��Z�v���]=}k��b��<���; �s;1I�<����庡�ɖл6��<1k��� �<�<�=�f���׻:`>�LD���;Grh��h=���<�..��F�"s޼�<n缫43=zm�8��;����lW=2vh���2;7^_=���\<�|[;��x��	O�ju�<6�;��U�#F��0�<��=K��cI�<V;L��G�����'=�=�6)=�3N��A=��(��*��C|<�̓<��)�v���J�������<IM�z��<Y�<ٙ5=�Aл��<���	=?q�<�Q=����==����M<o�*=h�+=��9<�<��N��R=�K�<���K[�/��<ώ&�l�<�C��h�<����T=	>=)��&�X;#��+=���:�u<��C;}�a��LS�j���K'�<�@��{,=zbM=��3={�[�=M5����<�)�<b'=��W���C�G�9�,Թ<��׼��y���-��9_F���U��H����6��
=6�:��nB=&�4=�'��p�<C�H=B���"�?=�p=C�=}��M��<"�l�!n�<�C4=�׼Ҏ������"�<퓯<��f�o��J=4�,=�<�N�<����4X����3�=��b=�&f�Xo0���v�Z@�<>-I��`��`��<��k=���< `@���C���l�u=]�^�~/���N_��*M�#va��R�����Tb%;�1�<��Q���=*�\=`�ݻ���<8~ ��޺Hm�<�xA=+Ĥ<�Oc:^`�)�=���O���X�Q�}���d=��(=���<ϵ=<��q[��Ҁ=���}T��$A��ԻN
=y�y=Dx�;1�{=wsd���<�����KD���]=���<Uϝ<H�<D��d��<�
�G===��-����<ܒ.<�.=P|_�{p=GqQ�ƒ�<P"�Թ���=��Z=#s�<<c=��E=d
8���>�+=���<�(= P<=ƄH��5�Wz�C�$�@ɮ<��)=v�ʻ;� A3��ׇ��di�唍<i�(�<�&��鼻u�<��'=�꼉�(=�KP=35��O�V=�=��9=�C�<��Yɻ��<$p =��<��!=L`���F=�7�'��m=G�+=�n=X�p���<�z��C�$û��r	=�=�9'=�WX�Zʬ�i�M��$Q=���$<���<���3D���#N=��<y����U==4.��$�ݻe,��ճ<��Z<6<@=��K=5�<?�9Ef�;V��<S_><V��<ue=/�N��h��d���%��c˼�?��>$��׎<1FU��ẻ�Hp��C�;��<��y�Sc�6BA���V�������(M�<PGm�:\���<�t���w����<�@=�ȼ�)�;߹�<�4U<�o^�N�P=-I<ub���Ď�;2�<��w=~B=S�=�:<���hP� 34�]����Ӽ�"��|#!�s���Ӵ<���<���;-�=��F�'B�<�,���W��;C���O9����A�'�=�Z<����M<~��<sc;��H��>�q�0��.:e�������x=�l ;:�=T���0������/ =��Ļ��1=�� =���<!�����<�n�*=�<8z�.3(�N_�<��U��m�<�p�<bټ�h��5�<~��<����
��<:_����$=f�m<q��<qZ�wG���T=����=:cs=�LG=\�;R�(�����d;��W���"'�,���AS_=�7=��,=�Rx��������<���<����X�<.=��(=����W�~��戻������36�<�^=W�?=���_��<�n�<E��Q�<�����!���W���<o7�;g�=��V�	��=�m����<��=�x��*4���B�d�<=�n�<�Sm���
=Q�=~�p��I;��4=g��<��<�GP�Jz+�*DX=���<n#Ⱥ��*�#j0�3�<�?4�-K=�.�H��;r��Q�� K(�����xV;|�3<�)�;��0=~�4�=��C=��:��P��<�IL�Ǩ�;����S����=(X=����|�q<�*� *=C�<��8�(��<ҍa�����w���e����<֟=��,�H>=&=��+�؆+<1�ɼ�ç�Fh =IJ=�˼)��A0���7=fv<'�=��=�./=�3!�Υ��V�6=�X򼙆@=U<�<S��_/&���~=��<��<�K����</����.���B��YF=��@=��< �C<�Q��� �<��I=/&�<@i��M��v�=a <��T��<�n<tȺt==��>;
J<���=аH=�HL<+=ۺ�`<f=�d}����Tƨ<�U0<�N�<�<���;���u�Ƽml=��Tt�<��<����^t�iW�(p=R�V;x�E��e>=?�=�C^=�YJ=�V��ԭ�2��ʀ�<ٚ��Qe=K�J=���<�@�<<��<�[�<��E=A8�:�����
�<���������j�<�Q��KK_=�n<ѳ㸾���P�>�(����Լ�NV=��<�QU�N,��6={�ʼ��o<����l&�;�<iZ%���<Pr�<�l=ޗ���U�<a
h��%�;oԶ<��;�u=z	���e��P&=��|����н+=��1;�mD��w��P���X%<H�r�h�g90�e�����<2���oR���w�P�=��2�X�W�hv��=ռ�2=��<3A����B�X�&ülI���U<�-}<r���#�C�?+9=O�-;�����` �4	��՗`�+=�줻�<(����˖<#�N<��
�*�|=.ܼ1�����=[�<̓��W�8=��l��9=��<�߀��W=��8�{�R���;<RC���5==���3q�C�W=Q�u���-<���Y*�;��;�@8�V�$=�+=��t��		����TyN=k���<=�	<s��<�Ԟ<�å<�<�<��g=˴`=�R#��J�<�8=�w����+���9�뽼!��\h��^,=��;$2*=�8<j�<��M�d_k�CH|����;N.c�@��<�3k=G䌼���?	$=P�,=O��<Pt��zy.=��)7u�uw�|: �ꈳ;�e��w14�l���=^\��;�w�o�Z�C<�T�>�%�]�Z����A#=L$��f�ּ/�0=��ϻ��g�
��
;��\��E=\�;�\&������:��2�y�<4�Ҽ��Q<O�5��n��S�<X���x�<+{�<�$7P��<=�yad=p�t� 	��!i�<�� ���<Ⲹ�
��ZZ<\�.=��y��漨�<>�"=��:���\�?:=c<3p<y�7�O��$�<�>��0G<����/�m9=����z�����<.G*<f8$�J.��z�;�.5�Q�<��$=g�v;��C=�;=�<	�i=5=`5l���� b���V�<p�%�p�R�1��9�o��*vv�e�5=t���f�	��<�!=����>�S�=��j�,m�T�=&F��(�Y=�x<��7�l�Q=�(�;R�@�K���[-��;��g����;�[_=Ib,�>	T<�G=Z�82]-���R�39d=*�=)��ud[=�� ��\��� p=�@����7o�<\=$�;��qh�Ɂ�<<�=�k;K�U�?��=KC�9G��<l�<5��<�ƅ���Z�T�Z=��X�]�ӻ�<��0���:MJ?=�y����<��1=�q=��+�V@A��w��أ��Y�� XW=zMd=�Y<�=%|���E=���;�42���(��o1=�����)=x��<.�Լ�L_��z=�T��Yq=��z�j^�<���?�<�ȼw���X&=��Y�U0]�1��<���|���=Rμ���:/U	���^=eG,��_���$����<��=���J�B��W�<>SA��k˼p�c��P�9�}�����3��E�4=��E�l���A9��=���=L8+=�(=z\����G�2��F�=�ؿ�̰�<B������<[���:��SK��<M�'=��G��K�=�v�<�ƙ=ZZ�����;�2Q=�Qm=���< G�����mF����;=m�j�Ooϼ�3=;K=��1=�L�<��&�b痼��_��L$���':�����<�Y�D�=Y�L�=�D�<�<����p�Jz�*I=��s=%��<�!����1ú׳ =�dh=�=Dl�<������/���w��3�O��t)p��u�<!��<{��]��[�5�� 7��RE=�D8=�^��رj=�B�����S�0=����(�<3 R=~�ǻ�<��x.���h�<�`��\
��:3=��R�ou<6�O�$����x=m��(+=y��<�IO�S9;$nU�Uw=���`�/:Z�;����8�	�Q�L=Tp=��ż} �<�ca���;���T��K�j��'��/~����<˗�<^W"=~=�J�<:�ȼ7�='�V�R7=��:=���Nk����:�e����K<�����<��l���K<�i�<UП��=�Q�@=��c�v[+=r-'������3�B��<߈�d=~�Q�߻��Y����/��<�ك�̆T�_�?��#��n
���>��P=$I=�n��R�u�ü�r;9����C<��;�@0=Q|<	%<�M��	s�kA=m���"�k=]'��{C��Uټ���;��߼��=�UǼ�!=-B��ܾ�d�}=6*^=�د�w��:�V=�h�<�j�<z�%��PQ=�>l;����<�?+M���;����[*�<��<n��p�6=F�<�0��-��z>��3�*o����߼c	f=�Z�UC�<�M=��`����1�T�u�>��=QVk���,���<�8����w�,��$=��"��U�G�G��<�߾��QM��7�Vn�<>rL=���<���*�����4}��f=ur]���
=�xr=���m<s�:�m�n<i�L��w����
=�/ <ҝ<u�ʼ���<�&<�ҍ�B�:=B��E��
� =��#=�A9=��B�v.����ђ%�X����n�No�=�y='�=$L=O�h����#��<�W�<A�'��Q������5<
��=��#�蔅���<D$�a�=��<��w=��=�=:�*�~����S�<W��:��y=�zN=aPx=Ж�g<��(��J�<qd���B=p>$=�&=�r�<��мK"�픽B9Z=�=���=e��<���<��;��=H	��l��Y�<I�;c=�Dc;�<޻�GN��R�pe#=�I����h4��[��LR=��ּ����T[��AE��}��'���h����<6 1��^=�����;*�Ἣ;�<�a�<O�!��� ��H1��vL<�?<&��!�*=s�<Qw���c�<��<_��<1����62������=����x��	�A��d3=3w=?�4��	��-�<`��1ڼ���1��*�~Ҍ=X�Z�g����&��I�;5������<��=��<���<ڑ<�-Y�iC�;O����#���Μ�����y=�� =���<m�������LS�=��<���<�K̸~�W��7=|�==S� <ܜ�<'�=�=�E�;��¼��=0̸� �E�g̼�����v0=��-��٪��y� �`��<(	D=�`��6==zn�<�; v��[�=ۅ<�(�9��8����P(�<8L=arW��$<�m��{R�.H=���<�K=&����=����Z �<�q��Y��՟��c6={��<Ƽ��=������<b�Z<�9G=:��w��<P��>��9^��) ;�W�<��P=��S</y-�X3Q��h�ui�<�/�����<C�м��7<)�B��G�<Ѕ�<�<��9=&7�+�+=�MZ<�h=��<�PM;/Y�<*�D=��:=�{�<�a,���<si�c�l<�4�<�逼�y#����nSY��j<�C���<��C���<M�=� 缹J�<�v�;#Q�<����M�i�L�|P�<�`=(�=�LS��{o�U��%決hi]�qH��h)=�4���"=]<S�L�me�;$k�<��Q=���Y�2�����K�����<.M=�B:z����o���=[Sz<:=�=@/4���G��r�<!K~�2;m�Z=�.��I=w7F�g¼�J�<St0���;�	�=��f��nK�6U��O�<����T(���:��;��v=c�<{�A�B��
KS��b<qH1=�<�<lU�<Z1�;Є =9 �<b"�������(R=8P=J��q����>��
R��G�l��<'Y�<?�$<�Q�c�a=Q��<Bh=�C�EW'�㽋�-z��N&s=l0k;�->�ҫ�����&�<�����E=᫡<���*;�s�<�`������&�a=�bܼ��G��n��=��P=�!
�YKy����ɚ̼o�#��̈́��x��Z����5=���P�e�3���@���8q��=��E�68=�4z�K�=<�}%=G-g��G]�ɦ����<y;E=�!A�޿���A�;��o=���<�FԼ�B��Z�<g�=�vY= c����,�X���=�Ib<�J�����- �V��<O�`�~��Qu,=�*��;Ct<�1�<T�E���J��Se=8�;i�<"J<����M�q|$�r6�<"F˻�v_�����j���n�g��;��\�4c�;,�
�9d���߻�6<�X��c����;�j(�!��<Y�&��{ٻ톰�"쎻V(�<�'����J�2���	ǻ�7�<h6P=�[=��3=cD=+�h�?����=,�>�e�;i�A=O�*;w�<��m��)�:A�~��!���<�z��O�=�����{d��y;���;ۗ�6�=V4��킼�S��� &=OA�;�ר<�z�<�;����p=j=�m=ǰ�<��='��;�:v��5Q=9ǋ=�u<�S�9����Y[w<5�=�E�Ԁ'�#x���N�=�b�<��<��p:V��M��=Pa��帛<����J=�J?���<ū&="\n=9�y�����ɡ�����6�<��:=h��<�>o���/��F <ī�<i:*��\<=J��;�d?��;�;Kg7�Y�L�+9�0ԍ<\4��t;詑�Ӂ���TF��G=tϏ<���<c�k=�!��P��}�	<R/�Y=�^ =�� =�Lv�Z�%�Xnv<�a=,�n;�@�9�Ko<;�6��D=c n��8c<�ͼٌq�W���,=�ͼC�*=�������<0t�	�+=Ite;���<�D�;ը8<�Ƽ�!��S=��A��10<����W=	t`����\@=Q�=2�[���<Ɩ]=>Ӳ��9r<d�T��Y:=v�=�D5����<�<A=�V;����ּ˕)��H�܎=�����d=2��;;:	D{<�̠������U���:�W�;���;q�^��T=pL$=��3��_x���{<:R=&�p=�~�;	L��У�<b��<t�:�\+��r/=X�)�+�E_���;ϵ��=r_�<��7�=���d����<0`��\=�`ż4���F;�i=���:��Z���F��=�� �=(�k�{��<��<�X�T=�D�<PW���7����<W�=u�~�6�=)��tͯ�Lo"��;=����"`k���=���<0=ҕ<8x�;�<9�5�{�a�"S1�	V����:��M�l=`�'=�=^< ��<��N=DP�<j�=�v0�G�=�r�=�?=��ȼ6]��^�dv4���S+;ƪ^�A�<4b�;��<�C�:#=�<��ջ������#<�d���y<6�!=l�ȼ��<�&����<��o�v��<��<�X�+�]J^=���ﲂ=�����<(Q�<}�N�����(��r� =���<�A�;4�;'kD����<[k�����;��y�!�L��eһ=�'��t+=�<�e<��,�S����1=ނټ��z=�U	<��=^#=�­� �a=Z�);U�<,�8=��üW�|���=P!�9�<�)@��n�;�!ڼx�O�~1�������XW=�uU�ݨ;�'� -�<IW=��-�e=�kv=�l=��J��S�<��\<M�4�TB�<��0=9o'=��u���M�����"����*�<���;X�fk�;�$=�s2�qFN=u ����9�f��6=��?=|�;Ա���j�M��/$�;�^<9��뿼�\����v�h=r\�H=���M� ��=9o^�;1����Z��dɻq6=6$e=�ȣ<�<ګ�<?{��V4����<(;�9=ɥ!��mO��=�<h�y=�S8=�9V:��[���b=�`�<~`=���R~�2-�<����y �AUG��6=s��I���*=�Y�<���2�<zQE=P��<Fq ��9�<���<�'T��Gn<¦�*�x�ۇ<!�-�(�Ǽ�C���@�`� �E*(�3��=Ϯg�k1��y.=E��:@������H}��rS=
�Z���׻F#�0�m�$�\<��O�<j�����B<E=<
���==C�T�`��<���DX=��
��=� ��0� ��+J@���P=a�N��Rܼ��;B><-h�K��<�?}���g����;�饼&�^��h���yS<�&=>�=�ªD<\cH=��D=�'�<MͰ����:#A�<�G�<�y���C<����&����<�p�ş�<��D���=��+�x==R@%=��1����;V>�<�g=�;�<�f����5=K� =�pJ��ڀ=��n<æ���<��|���<m�q=�A9�2=�� =n+��E�<���<��<�	'�W[O=w�i�W|�=6�2�9�_+ =�F�<�<Qq�7�=� =��+��D=Q�;J�f�z~����;�F���؈<�F�<n��9_ἔ�/;�����7��"=��(�����Be=���7ʼ�h�=,x0<�_P<f^���Z�`V<Dq�<��O�iL=�姼�N�<�1��Ἴ�9!=�8��� ���	�� �<�&9��Gq��+�=��3=_�LXG=��e�a��<<��<������.��lc�s�F=� �0*<���<r���_=d���(�F��_��+����=0��;$�%�x	�i�X=�<=��o<�������"�<��H���
c	=��+�=p��U�r=�><�N;3�%�}4C=^�:��<�漦�N�к��ݍ���"(�c��<���<Ӌ��Ю=�S =&�r�������<�$ļ
0
�"�=N��Y
=d�c=\�<l`�;�'=%`=��V=�T�;�j�Ͷ�<n�$5=},�;�8��r��/]�3����I=]�ڼ��D<[�<I�@���\��R=L��=�N>��QD�{V��0���,��0��<%�;[ �<W���t<<�=,-��ڤ��� <EWP;vL,�2�?���f�i�ϼ��<�$8�)��?��*db=�W=hμ�P��i=�[<���<9b��'<	c���{Ƽ��˼�\�<�Z�����Ds\�X�<ӑX�� �f<��%��?�<7�ܼ���<�A<=q��� ��<B�a~$=����/<�4Z��%=su�9f�g�^��;k�;|N=��=��=�ջ���b3=[~=�wӼ�<�=�ɳ�d�3�P3<�,��%��2J;���z��<�^=�J=�z;�)����0=��T�um��G�6��w(���==3ag�N�J�y�/��� =q}v�G��<fcn=�S�;mU���ˡ���!�]z�<X�W�}Ơ��ׯ������w׼sx=&4P�4=/;v�0�S(�¤|<WP=.���%�����;��O=�Ei=�ߵ<f"��aLx�i�"���=�>���&;ړ����<~��=�K<�-=�	���,��漶�7=i1H=S�ڼ�#�;XpѼ�&�e���S�=�e<��3<��Y=I�����7=���<)z=�4=��X�\�4�t=](��<r^��=��%=�h=���<��<7��8���jh=�VJ=��Ἄ�$�@�5=��U=��O=J�<�X=��ͻ6����P�<�/S��L
��8�]�*��A�:��c<�t�=Qf�:�=��<�y;�}u���(=h�=Vc�����l<�?=�� ���<�ͼ�{���W�m=:�U=!�<��<f�.��#�:��ۼi
��!=�k���TZ=�+�<S=�:��\��<��+= 
����;�H=�q=Qww�!!��df$=S~=�X���*=o/=�$<�I<�q=�K�vt=a�=�=ɈX=���z[9�CbA=Y�/=+�F�@��8��=��<<ռ�;�U��C���[�������;!�����<�- =>���>���h�<�O�<E�����=|<�_<��<� �<�=�=/ֆ�+ ڻ���JK��C��<2@3��K��<��ļ��Ļ�n=��d=��&���6��<_�������(2=��(��Z=��z��z��:���K��?ռj�=SSN=�7�;:�׻�.0�|�N=�x#<BZ�����bW�Z#�V"~�"=�����e�;����5�{=�&=��T=�����.������<8�#�Z<���;Ԛ���<ܺ��l����<�[9=�]��;�_|����;�9�<#&�bU<=��y��S)<��<pO�WN=�v��Ƨ�qq��$�o��Q�<>�~:Р���=�<�;�������XU0;rq;�"n�@]���]�<�n��*CS�/}A;���2}�.~�<+�����F�\�g��-�0��<0�=�x�<�� <">.=�����;7��2��0��<=ŭ����g~=�1�\6N�y�����<h�p��ȼ��<G��<%������:&>=*�M;\�B��.�@0&��ݯ<��^�no=D�<�v�-B�ҷ>�)�;=
��D"��X�bG
=AH����(<�$��'Yh=�JP=K�Ѻ]}��.���|�I=�|j=���:A��;`�f=��:7҆=(׹���<z�C=�<�Tw<_�;�=�<����B�l@��m}$<�mm�S|�;��<��\6�<b�#=+]���z!=^b����
=�*n=z��<�.��伪�m���~<�§;@��<0\h�Z �<��:d]<�Fq���ۼ��R�;�d��aW�Hn�<:�<���<S���|��3����������	�׌P=I%�����+��\��|����vp�<��G=��[�`�<a"����=H*��g=8�<��H<#���T��;��<�2�;��d=�c�;��-=�Sp�D"0��cD<�F=�=Y��kϼӌ����<���<���;����^0˼�:={9��m;Ϝ��������;�Zn��S^�"�����<	%N=]2<����<���;��L<3��,/K;m�^=Yw7�<%�;�Y����(<À�<R��<�h�<Ffd�i���v������=
��;�f�</�B=�=�r���P< 9��"���f,=�/ϼZ�[=>H�NK�<ͥv��m&=�м;d�x�i�}V=ݙ�:�T=KD���go�b�ʼ�+�<���O�o=}$L=1�=_��°�;D2:eSȼ��<I�=_�p9�DC=���H;�<�":�r�s�"U:@�V=\j5<�)�=p�2=MX�t� �+�:B��~@E=~oK��?==o�Y=χ)�b5:��U�`V@��	���o=�{D� ��T�U=�T�<��<�����P��ӑ��]A�N�Ἱ����n(�l�̼�T=�
�<R�o=Le�=�)*=��;5��<r��%�<���NGH=����W�w4�9#=ߩ���~=�s?;��<�P�<�=me�<:@���9[�eH	=u�l�U��P��<^sG��]�=�.v<:�A=Z�*���=�J=�8�;�%�<�~6�F�"�� �<*6\�v����,=	L"=����?������&���y:ҥ�:�·��V��a}O=<0�<O\5=�����ɗ� -d������<+�S=��)=DC���:��(5=a�U;|�'��o����=�jd��=q��;��7���=�Մ�6�)��z�=��qX=)O���B=��]=�G;�y�ѝ���x0=$!���2G;��/=�AY��\��M��K�=_�I����< 3��R-=]m���c%=��~�;�D=[��l�U�ۼ�q=��Ѽ�AC��=Q-�<X�q�����K!{=�#����u=d��`7=K�^a!�'I�<�a=�*�)h��[4K<t��<��v=�+=��<	�
�V�6<}�e��cU���9�������<v�<ƞ1�+�<�+��b��<%<TQ=�м�#���\=Å�<_߿<�y�mqJ=�Ø�,eg����;�&4=z�<ṫ��׬�*ۼOe��K:,=fJ��DZ<�?<Գ������¼�Y;�`/���<�z <����C2�Lo��4� �<�m�H�A��3@<n{����=�f,=Bn��t���<n��eX�>�%��I�';������O!���	=��-;G�ؼ?��<}��;;�;]j�;��6�@?h<Yz;�,���
=�1��SH��_$��g��E�=dü�y=0=v�Ʈ	�����=��|��J:Qü׀p=�C�<��M.���+=9[u��;_<�c��Q��4�̮X=�o<�Ә��s;VrM�@������_L<��#�,=\=S�<�}�<~b�;U�M=����F�;uk����;�h��=�m\��FƼZ��<8��I�(=U��<p{ۻXhV��t�<���>x2=b�<�<D����<m��<E�
=%=��Z=�#�P�=핼��d���L���xμ�CI�&!����;�� =4�zY������`Q=G��<uŔ�&S�$�;ܚ<����Tq����I1=�6=3�(��1)=�VB����t�<�근�<$Y�<˨Y���':�7K���=�5�<±�<N�-=�;C=�tY�g�B=�@�Fx�j=���W�
:=j��:��,=�ƿ�"�=����lg=D&=�!=�M��<�=��5;��#;�8�%{L�rT�<�L��ڸ9=is�\=��s�FT<�o��A�s�<�i��֩��tغX�V���&�$L7=s��;�Y=��<Ӏ��h��(��/����+ =P|��ʮ�,"=/�=#i��\=p�]��^<�3�<�7�c�鼕CG��x@=��=�֝����<��=�Q�;I�-����<�S=g�����%<�JI���=�S='-G�&<*��;3�� �`<���<��;>�]�<s3�a�b=Rm��i#=ݵ�*��ֶ<���Df=��=�����<Z�-=!@�<p�a=��`<��A����22���8�=��<���<��F=�E��5��Lt=�V�=*z1<�-F=
��<�=���=g6��H�l�W<��<w��4���<˟�;iU���#+���8�<�)=g�.�AJb�������-��*$=m��<���;ٸ=����2�R;.2�<.�b=M=`>�:����<͋j��_+��^=4�="�8==��<��N=�=n5=���<��<=�[=\�����=4?�<�����@<1<żu5T�.g��R<s�0<F�<�D�<���[�=�����ZV=������L=�J$=��,�f�R;�-�����~0=B_y�l�T=J=���a5=-{�x�<��?=8��9���72�MvX=ضS�6cD<w�<� �<I/���߼׉��ҫ<.9.;�g	���l������	<V� ��=ס�����<���<t�+=��B<�電a_޼8+�<�/=��W=�=�~�G=<C��4��<X=v}���g'=b�=�~)=�|��q=C��<������mk���"<�A�<�<+=`=���<��8��zJ�Okۼ��h=�	��}�	���<�4{�ݍ�<�
>=E������>�#��:��=���Ѝ�_9��U绁�<=@��<��==���<B�����?=/�u�ȡ�<��I<).ͺ�<M���<�G5���u=���<��9=�Ow=5���B�;5�����\;T�V=�+����K�Zr�<m�D�M����01=�Ѽ*��<�)�Y�J=C����t=��7�ϱ�RG���b��$T�;�
�>ܩ<��7��ۀ�ř&=9��<q�/<�p�<��2�%=��<n�2���ݼ�tp����҉F<�r�=m�E���@�N�� ��<�\@=w1���=��D�i��{�<v��<�Z7=']=&�<��0=��$<U9¼��j=>��<��<R�B<�<v��!= ;7n�Gk��ki�;�=��Q�^b�o�<9�ĻJz�<�}����#=��;C��<ξ��#��Ak;�a껷���?<��}�^��<Wmi=4�#=��_���-���&<�����4�Z������6[��+<W��<�'R;�R=��<>5=�#S=�A��$�:�T�<R@�;g�B=�Z=F37=��ּs_��ώ���\��¼	����=�m�<�;۷\=�of���V��9�<�=T���p�ڝH=��.��G&�c�Q=\�';�bh<N�];��<��U�����RxM���,�z;=��<��=G�����<b
���i����/�=����B\��,C=J=�ʉ<��N���Z���I<�?��`��v��<s�/��\���Z���U�:J���м{�04ż���1V�A-<�g/=�@�<s��_�:4�w<v�輠,�<�j�+��<~� ���;�z���0=�8J�k�c���K=_bk�b�=�����<��<���-�E�<-8�?��<¡�<�n	<�����2=��q��Z�J<��X=�6��� S<w��s{�<^��<���;
��<A`J�}�<�s���O���÷��^	<$*�<�aƻ���<���"������/�ź�ּih�<K�1��(���k�����0�ղq=᮵��ӎ=��;�$=��^��O߼�R|<�o6�j�J;=J�<]Z�;Wr����^=�T<_F��{�m=2���� =�	�����C�D=���n{�<�+*<@�ռ��%>:=	��=㠅���R=���Ao=ڏE��E���3�R�h=L:&���<n)��@�=]�4=��!=�}X�$v4�T6=���=�n=Ѐ��OM�� �㼞%�Pyx=�Y[;�8=���g�=��O=�tE=X�H�y}�$!�N�=HJ'=
�x���ּgų<�N�;l�}�i<��-�+����,�;�o<���a��<���<��=qֈ�N�0=�=��rD<���.w,=U�<�y=��:�ٰ<927�
h�;_h�<W�L��$�;�Kh���L��n���z���l1=��";X�2��.��6�
;X���x�;˛<�K��`*�Jѯ=#>=G�뼑���Q =��=�`һƑ=`Go;�ً�u��6�<�pF��,R�ne�+���6?=����{��OS��O(=���<q���'E;3�=�"�=]dg<)�Y��K�J���Ib�Q.;^�S<��=��;s��(44=�<(�;k��<$|��6{6�#�����<�K <�؄<��<�K�<�^�����;�<frN=��<�=�K�Zw=%м�7t=3,�<�R�<#)�;�����<��<#:=���;3t?=�y�%J<�酽�r��<�<�P`�R)���+[����܊G<K�ټ��z�υ�7��<d��;ޢ�:7=�������~�c��2	��j�sӾ<�r�<��R<a,=�3h��u<=�X==��Y=�_=�-�<��ػ.�U��h|���W=��3=%m<B���,p<@���p�2=p2(;,�N<�����	��z/��4|�"5	�P=�<�3��k�s=��p�Ѽ)=��H�9;<;?J=�����lN��lq=,-�
����߼Z^�<���`\_<��=��S�5
ü��A�\g=���<n���m��$/���Z��vI<��������w/���0=�a,���\����<+�����=��=M�a=��K<oeҼd�3;���<�[��/s�=��<�o:������19��T�*�-�d�;aR����<{;���|<�D=E��;^�D=�T<���<$��</?�V<4=�t=�b̺p��<M	T=
�ټ��<�_1��
-�詛��򰼕��<I��/]���&h�K� A=��n=��v���d���7=[�pT=�Iü�$ =��2��=.n�����tx^���=>�l=�/N;DU2�S��<�� �5=�t-=cRz�m����؆=�o�]��ס=&�\=T�x=� �<Y��<����C&��4`����<���j?'=ϘV��^�;x6F�{=%~�<�+S=e�*��] ���]=`�<�y=�⵼>�^�2��JZ=c�S�+֨�j;��@=5�<�������2x�!�[=&�J=u�o=.��:�\O�����gR#=@^� �<� �$59=G� �O��;���<��I<���;9�j����\����_�<Y0b���;@��PǄ<7�'=s�F=�C��=�ٚ<fS �-i=𸙼\�
=�-���A<432;1�<��S=�9���Gb��D�<3Up=N����u=���<�8���8�<��D 1=���� <?����<�=4ļc^5�j� =-�H<y�1�u���D�V<�i��c�R=q�$�X�]�3h�=A;s=47�<���_���<����:=ͫX���7�%��<g5�+(,��85�x�b<y�HZX�bV��
�N4W�𣶼�k�=�!����*	ʼOǯ<F7>=wu[�Ԣ�<�ż ��:�����$= qL=���<�_`��,�;L�a=ɍ�NB4�O�<[�Q=2�<����<ϵ�<Ξ�<��J����<�S�<��P=��=���<aP1=)��0����<�[C��_o=M}<�	U<�]�;1.<���\�n<�D=ç�`T<�u�;�ZT������Y=p�g�=��l=�A��Ub :��<&̴��}�Is�ϵ뼌�v�l�^��鿻~dQ���2�̒_���R=��4���D=NO<�:=7�W���R�ж�-��:}J=̔�:��C=:���:=~N=��;<̛<�e<�z�<�g�<%|Q=/=��=�?���f=iL|=f��iۼg.�<�By=�]�� �<Χ=N7�A8�&�	<K@�1�/W��$�H����ڼ�>9D@=8�F��󍽬�=�D=F�e�j�D�%"C��A><�%�=C��<�Q?��o(���G=���<Uk�(Q&��er�>�qU���F$<{I���3��������!��"=��=��������6�=�����d�!��ћӻ���Z<�E�<}�޻/[����=�wO��m=�#��[��C@<F�=K��<�.�0� :�K��L�<^a<��O��X~<�G�<�ۼ��<�k���$p=x�b�8;�������tR=0U���L&���j�=�=4û��X�(��<��<����Pf�� c����<i ��
t˼`$ͼ���'6��q�.����d��zà<iwP��C=i��<{�f����<r����j�<`��l�-<�X�F��� t[�W�X���<���;.1l=k�=J�0���}<�f)����;x'����<� �<m��<*�);X����+
=*�<B��=��{��5=�J�ܩ����ڼk=�'=3bI=�Xl��`���N�f�Y��*�<�0�<.��Z*��Q��l���]������eW;�fT=�pz�I�*�i�Ǽ=���8	=�����漒�q=�pN=��=�y�;�;�;Y%��D?=>F������);*=)F=�V�	j�< ����$=���	HO�4���l�	=�$E��?g=�ɼ}��<|휼#�w<����t��m��Ĝ=���;T��<W�g�k�s�y�6�|᜼�¼g�s�m����<����� j�5�<�
���b<&�?�N�c<�L=h �<��;=���<ҧ��5=̾=��`�%2�<�3��V�<I�=z���bi�ð=�����6�ۃ�<��úI�=� ��=j�X;����6=0��<��_=RX�֍2���ǻ;=�Ǆ<9c=q�b�v��<�b�=D6�=�g���"�����^�,=��ϼښӻ:=^s��n���2�<��=�D>�,���HA�<�Ҽ4�+<j�,��W<gJ9�&�=~�`=1�ϼ�A⼹`=�H]=`V�Gr�tʪ;�tK��|ٻ���<��(�����=M�,=mZ�����hx=���<�<;�*7��5.�=]͐<U�����J=nd��<�������K�z�r=a	�<n8=�͵;s�Q�:�߻g�����<J3�k:��)=�0�<����t#Ѽ�P|�̡;qV=�$���%ݼ�ڪ<��q<�j�G�#=D��R�a��ԍ�l�S=��k=��T�a0�e�)=�t=��;��<���Tw<_Y����<���r��C�� t��P$< =���6b=W?8���;Ӥ����;a� d�;H��<&�0�7@�;�識��1�g|���
J=��,��A�<��S�C�J�Z��X7���ļSe)=�,;�E<��z���0���B=~��<�h,���Y=)�$I����<�L	=���RD)��'#=.����L=�� �Tg�4���V�<��P;@��s�	�%��؟��Or�c�<������&��Ye��d=j�ݼ��<k��<��;��<Ћ��K�<�53=K8�<�I�<RX�:o���l����<[�=�<2�r.=-=='��=�$o:�%z<P:�1�J;검<�#<|�]=���a��+�C<�L���`�;�
��.ʼ3�	=�:#�$<(,=m�μ��<�8��(��7��R]1��2b=��P�yf���=�g=�kR�Qb=�2��㼁m�4!=[��=��<gR=���ɺ/���H=���t�+=p@�<{�f��WC;|�q���
�L��7f<��)�A���R=G���Y|D��O�<OC^=��<ݑ;"k�1(�;z�����iK=�e=�F=q���L<<7{<.�j�|�I=gk�<��}=9sQ=D�A="yͼ�9���<,D=�	��o[�<��:=rRr���<b~�q�M��� =�@]�CQ{=���ӵ�=�w)�c�<�</��<��<��==k�'���=�5�c�7=;3�<��=<�%��& �L�^=u��<��,����="����<�B=�ߝ:⭻�����y=���T��^�g�5�L�bP~:�����<Ot=p:= ����$}=}�;=}w����"=��=��-=)S3�a�=��<��ټ�>s<�\�<��<��J�6{s=�A=���<3���5�<�B���	�CJA<��(=�JW�4�}=΃�<z��<�9=��̼�qƼZr��.�=%�:=$�f��xǺ�ި��<=_�::���<��k����;F<��<��E=�u�16J�<��;����Kû���/-<D ���Ƽ���:�C8<9����h{�<�����s}�1X��Y��M,$��0X=_1=�6���V�<�LC=K_缬9$��Ia=%CO����S;�^����=sN�U��.�o�ܼ�8<O�A���ü�0=���:�,5���T<}[޻+{��E��8=��F�S�;S�ј��aϤ;�eb=�O�<s�]�� 5=�	==��j����՘6��dK��� =F<.=�<Z��<�ϒ�Um�����<ά��Vt��:=�4P=.�<�~+���C����<P@�����:��=ח�=���G�<��<}%�;��:<�5���<=�=g�0=ޭT�ʔZ=Pl�4UR�+��<qu2�OIb��n�9�H�<sw;���c<�X��������=�8=躲<	Il�Or1�V_<?�Ƽ��A=��<o�0;��i��(b�P��<�䋽���<?�v���=���<�j�<��H;Q=&c�<�ƈ����=}�H������I���=��3�G1�x�f���|<(4���\�;��<N��<�n1=�nܼUi�<V�����=F�D;�'<�N~ʼ��H<��#�Z�<%Y�<j#.���;,�q��Q;q��;ƉI�PT�<@=��89TF�:��<����ʴ�c_��Ԫ�<�<��O�(K�6�=�λV��&-=w/3<VM�;F�t��&<6�'<K�7�G|=(��;N9=^<��
��٥�v��;�TQ=�W��Q��<@��̥�PR�<�l�<�p׺��mI�<Y�Ǽ6  :�&�;�����=ylT�P��=���<ګr<��v�B2�G���!�;�&󼋵z���G��4O�)P�<sB�;=�\�V��=R�>=3�~��K�|o<=��/=X�+=���<�.�B�n<���Om+��7i�=�+���%��U[<
T������<@�u��K�<v�<��=�<g�Sv˼XG3=����㻥�)=�<_<b,>=����ݪ</	Y<+� =�#�<k�=%p�<k�:u�;�X&i�"t�
���l��<���o��<��<LQH<�F��O<�&=Ȑ��X/�|�=Ҩ�<��c=���')�<Sb<
��cBq=��o1	=m�S��c�Ho=qš��
���x=N#<��
=�?I=P�I�O� =�rm���H�շ���值��#�?2,�̰������Ƽ9ټ�`���~G=�1���V&���<ІD<S��81v=�:=�8���ro< ��<=��<:�<�=n)j�8�(�|e�;*d	<.,=�����<���G&���^={�=s�R<
|<=��A=Gq4=O�<�6���&�����0'G<p7=s?=��N� "�;�����r���<��SR�<�֬��@<kV��z%<����;�9<�	=�]=^K�<�إ���#<�6=Xl�<e�`��H�l�º2 <�i�?�=�3<r(|���M<#��<��7���B<w��X���.�2<�ռO�f=�U<��d=�=�pּG����2><I��</�˯B=Z�<k�/= �	=��<=dC#=��=i�<H�<z+=#O�=�+���M�rRx�o3X�V�=�UB=��Ҽ��r�f��;�k̼��E=҃�;
|�=��>���i{�<�G+�*��<���<Ƃ���d���$=�U&��I�L䖼�h`��5=w�p=Lu!�_�=�i=�Km�+s�<��ڼ)�<20=ӱA�f�%=4�=��~�.l=&2:�A�
��{0��;u�-�|<��L���=D��(6�@��<\����"<$�<M�I�Z����A=���<[^�<9���P�<��=�8�=�<�<��3�M�-��(��hq;Q��<J>�<��>�&��<��S�zp���J ���,:�.K;D_(�˦=�|s�E�c<�V\�j��D�=,�K=���<���<	�K=%����%<Ҭ�;8y�<%r= $b�gv=�"�͆�;OD<��k��7�<�8�<�m��<��n�<*���)�[ �<r���.U<�k�IVC��s�;��M��ɠ<K����K=BR���<ii��V���RѼ���d=8����b<�M�ɧ��i��Z$>=������8<�s�<��<PX<�~I=�LB����<�=.��<�JO�J,�<�EU��I�<tS������t��\<�==k	5���(=�>4=]�߼NPK<�M=f�F����<�l�6K�<�g�<��-=�t;F����"����k�,�a�X��"=��t�;����R��@c<�� �"�<gF =�@G����<��w.=��|�W�(�=��ֻj�9�ʿ��Ү;S�-=���1Y�;��<��*=�=}�������=b5:<X��<#:=��G�6�)_@=��E<	����M˼]M�����U�= �_<1�����=U�$�hݼ�m��:b�=��g<5tG�Y:�~jX=)��<l�<��S�e/+="Z-= Ө�=�@=��%=��S�p<�6�:��<�3O�\�h<�E|��2ڼe��'��<9:�����<5F�<�,4;�����������Y��������ծ;�F.���|��NX=+$8�Y{y��
; �>��Ġ:�׸��n�R>o=�&�N�� �=�=���ևT=�=��&�¬@<��}�����=�L:n=��t�~�r=Nh{���)�I��<��4=�G�U�B��9=��{<k�;SF:��X<��$=�%Y�	��;뜃<�;�rڼCP�=h(�;��%:d�H=�CG;�2=3=�$;�����kY=3P������<9����<C�=d�=b6�#m�<y�A�5O!<�@�O/�<�:=� = �:�|�=#8�h/̼ٟ��K���ja:I�F<\�ϼ�<=f(��=i��Ʒ^=�<=�aR������\=��%�h����&�6�h�X}ϼ�"ּ���<[>�}�L�C��Ba�s�)��,=�_��b�<d�V����JD;�6�c��s�<�r=�sI�ǻ�1���y̼��;�
�#�=꣬<��S<��	=I�C�(A���=�o&�<D�F=��=V(=/1A=��`��`׼�ƙ��?�<�[=Nb/=^�߼ߙ�<�d��'����]=�$�<J�;"=�qR=�A�i��t�<{8=���'�V;���;�E�NL�<8�O�8Zf�$�Z�ޅ =��Y=_(��VY=�t<�L<�@5���S=@��<D�<�[�<�+=I��<�T���_=��%=��<3
=p��w��<%�Z&�7�1;g�@=����h=��(<�"�<ǑB���;b]	�贳<VW=6b=K��<�]�=��E=L�J=EU�<�8;GQ��d!h��n9<H�?���D�m�0�zf�<��F=%�f���5�Wh�<���<a1{���`=B�����;ŷ��{���<�?�2j��Ɵ����O-]��K�>�
=�˻����
d=%t]�"]=���<�E'=��H�y��2�6�p���J=k��<�YH<�ü����e+8�]�<l1+��r��Pf=fU�<��t�@�ۄ,<v=<���<?��<��\��0=L�c�"�����p���K�R�<�6=�@6:-A=�3B=��F<��J��w;�|�\=X@�<�q����Nn*���G�I��<:��<���LV
�vw(=K}g=�1>��(�<U�q�)�,<��<kb0=b�=7�#�y�)�Q����G<0���E�<�O=����k<���r����k8����<k�n�%
=)
�m登�&�=�q��h�;`��?���4�;�9���<�<^��<����:�<��(��D��5�1=!0=���<[�+;�Y�<C�A���'=1�<��}���YK��a��S̃�L4=Y�*=��O��ἣ���Y!�<\q�$A=��<J{\=ݼ��J�����O���H���9=ӆ<���;M��<0Q�<^)�<�N��5�����:�=���;��μ��7���R=QȤ����;o���e�,�V�����=�$^y=��t=e�����<s���>l=�x�����O�<@�&��,=yg=��=�W%=%C�<�)�.=�U�%�[=��r�{��=>Rռp�5=�s=�+V;��
�K����3���U�:�/� ,A��B�<�yC<|=���u�P��1
�D���r7��3���3��0�C��ּ�-m=�y׻�u=�.=��R�5o���<��#<�H=wR=(�Z��"�=-=3P��a`�]�wm���>=��p��)#=����dǺr��-����������:,7H=~�~=L��<1�Y<�t�6�Q�7	����<���������$��u>��5�]�a<��8=�l�=�%=�Q{��Ó�7'=��<�kF��{�<�}	���缐�O=�s=C(���<�7߼M��;��5��%�<��}�k���n=F���@>	=����ȼ�N�<ItP�N�O���=r'Ǽ��=D�/�T�K=���<�G�xW<W˃;��R��N�<�̻�?��;E���ּ��P=��<���=���ا�y	�;��=��<@���6`��ˤ�<����;ĻA�#=��<>A�BX��{<�
�==J=�@(=hk<�e=��C�k�r:g
<���;%��>(м-󁼘M���i2���l;,��L]�<Ki�<��x�xT=.+��Ս�;-$E�vK<N��;�e]��e=~�;�����6=tbR�����Pʀ��q<u�p<��=�;���?��:�A/=��v=��S=��
��I�<���=SG=S���m��C=D�;���9=�;�z<Aͼj����\��4eT=X仺Mp1���4;��T��/�<���<a>===ԁ����=;kq�%��[����l�m3�< �<���P=�N��1�;�l�#;=����'�2f=Uq8=�b�;#�@=��R"]=���;>A�;�1���<|Ca�1e[��4�;6W�v�o<��]W7�VG�<P�����%����<�u&=����YxQ��'<�w�<�uw<�ܼ���F>=�]=�;�N;Bg5���9z'<��X=�'=xw�<x�[��K=)(.�Y��������C=�S���<I���N���A�u�2� =V G���M=�t=�ݟ<�w�:u�l=�4@=nSѼ=A)�|Wm�o��< �g;�&��x�;&�= L��+d8=�[��A�<�߼���<�����<�&c;�It��SC<���q����<Wa�</�=�7=v����jĻ+Ӽ8M}���>����<* Y��/�<^���1�g���A�ÆP�@2�d B<��=��K<�LB���'<cS�<�R<����<^}�<�`���^��� <�%���T�.��g!�:\T;���1;c�3=|�3=�r���$����k=���e=8�x�� �<�g=	[7��F�\���<�
D���
<<l�#��<��5;$E��l/����uڻȍL=���<���;�_=��<���B���pT���Y%=H2���6R�0C�;q<=n�<	�:=�	6�*�8<P�^��w?��eG=�~˼;�:��3=\g�Z���{�<��5��-�;��;����OE;���<��2=�&
��H[=���<k:=R�h=�<��j>�C���F=~(=��=L���'= %J<��g�P�2�YF���X<��=���=;��:P�<|�u=F���5-=�XG���/�6v)��(<���M�b�b�.�_O�;�'�<r��<�%F:e�h=�j��������y�)e��������;�==iѼ�Tt���.=��޻�r�<Pԛ<_"(�W�=}��<��!��H<M=����@�X=E�p�:U�A�z��g���<g����<�<'0=��A<< [���I=��Ǽ�z	� ,�.6Y�:�=->��VO<�s�<s�R�9��=&��1<ʃ�a�U�.m=�A�<��+=;[=�;?QE��':�:>㻃w���}��|=)�<�<�9�7�$����<�� =$�%Q���+�]�.�Qt=����	�!e�p���\b�㤶��mw<�1�<ޢ��0�ӻ��<����%�&�
༭U��.����<]���ڔH=� <�ǥ�vn�<����=\�=<lt�4�5���L=�]�<je<�==�ٗ<#>�<ғü��=��W?��s<�=��1����;8�,=-�μ�lq����<x���$�y�>p���-����o<���<ʇ����M=|�=P<�����-��������;��z=���<K�O=Y��;y�=,Ж��d<��μ�pP��L�����<�#+<��̻�6�;��<��'���#� 3=��<���qI= f<�%����;�
�v9�<�J_�Kc=qC;�5ż$�(=�_����<�E�3M��Q�<݃��b}K=�#h����;<�&�k���m]��>&=ߧT<��"=H3�<[C-����S'��j򼏕=��!=��2�3�g=.�E�[S���v��=��׻�f�<���|T=?�a��s=fF:n�M��(A������<�X=v@ ��%<�x.=���f!%=yѹ�/^s<D�����ρ��h�\������p$��r<}`'=r���/���6��A=��F<�,3��`=�b"=m��<D�+<3=�)X=&�="�X�����D�����C9�#G�<�_=JHͼ���<e��1Y�<��:po���<ξ-=),=�<���;���<��D<e������.���!����]�Mu𼉃@=���9<(Q=2����<H�:�D����;�8߻7�<�p����<e�)�D-4=����>�G�^�';�\Ҽw�:��.�\�*=$�l���h]c��tB='�7�m�����)�a�d���<��=M���f=�Q�<�6=S�$�>�	=��4=�r���?=?��<�[�#T{�v���s��:�ۅ<S�e�衼��g=�=Q�<��'=����E�F<��d� �h��b=��;p�;(�̼϶�>�</f�<�\"�l����л��;{�<�2�<�=�� =��:���<��	<2����ʼ�#W;J|����H���d=�mM=f�Ѽ��S��MX=O	;�R=qaR<R
��<s�=�%[=~<<��+�S���N�<�<ŝC��^|�ay�<m�3����|	��7�;�Ae�ZG�<M�];t		�BqO=�����K=w}�<S%b=�Q8�m =��A|���[4��~���H� ֽ�$"X��rs�'�=;�+=��=Z�<�o��L
h=������5=��B�p���F=s�=Y�;z�d�$&��R�W<�dT:�����;h��T=v��~+=��ϼrn�<��l=�Aռ���$�X����#�EC���w,<�Bx=�@5=��s��mӼz=�3����<�wl=��C�(����S�<j)e=fE/�6  =��伜w���W�M�}�df�L���*�=�A5=9;�H���/�=#O	��us���=c��ܯ�u\=���<�=e�� ������<?��<P�=���<\��<,?м�%�c<+=�H��Z�`=ѷ�=Wa�e
�W�<t=4.p���t<����#�<��1�&s�\L���;���;��:93�<Rv/��]�L�����;�Iu�e��<�<���u�U�w�=�b=,�<���<O-]=��<�<+�.��� ��ז<�H���A���U=Cؼ�:��<��1�D�8=M#����b�y=�}
=K�<-�;���;��N=��[=X �<���<f5 �ˀ8=�����+8�b��<�G=t�[=�!�< ����3�Z�2=�<V�� �<�(޼Q��N�:<Z&��!Q�	;7<M8i=��P=�ᶼ�V%=�����t8=�I<�Ŝ<w��p�~�h��ɱ�>�y=�d=]Ǽ�]=�5�<��ݺ��<�\!��d&�ݑ7=��V���{	�<Fޢ:�ϼyռ�$���]<� I��� �2K(=`I~��-R=JS=�=��%=)���k����<eQ���=$)S�-Ǵ<�5F;M�Ǻ��~�n�o���0=,�U<��.�J��<��Q;"�1��2&=��g=!�a����و;}ɼT� =��5�3=>T=�o9=�
�[z���;nA=��f=p���jso;$�X=8M+���<��Q��mj=ߘǼ4{[<��;,�q�i�����<��4�`W6�m=�BU�����P��C�����@ =�.U=2&�;�M�;�p��<�X�<��>�]Y�)�t�f�\�j��֯]=4��<ӄ�;�<*}̻���<�5��f��<K�3�Z�=V	����<&�ļ�RH=�i(��=|����S�v< ��%��^�λ��p���P���:_n�<�Z;=��^�Ӕ�<�&-=H��<Ȅ$��l�;�+=ڨ�<��<�$~���U;q��Ԅ�lp�;8�-�C1��BY<�Xy�{�=��+��3=�����V�;��<LH_��V=Q�9=#4����<�������ļT��'�ʪe��+D<���<�s���DQ�&�=0�ټ��P��;����rB�b�=L��ʢ�<`eg���;��ϼ���<WfK�<OO=O� �<�0<�m=���;,��;�W��N���]���q<�@>�$uT����;E[N=��=��*<�[ּ�aS��=��^=3>.� q�<g�?�����8�� p�<1�<V"=ن6���+���=�m��p��6%�5q^�3 ,=3�G�U���d�t���(���U-y���v�ŀ���Oκ]�6�Mn<��e����<c���E�W��<`,����ɼ|X���$<P�¼ܼV��|H=��$���ؼ_L�#A2�SgM=�1��T�<-�Ǽ���I���Vr|��1s�d��@�*�1Kظ~�+=cכּI�;��K=4�=��3м�<D=��%��9=�m��-�b�Ԟ��П.��$��g�-᳼�n4=�[\==�=W�d;A`��;�O<�����<��NQ|���0��$o�F���-�� �<�%�^Qg=��;�J�;!>O��LV��L���DB=�$�<�~{�(-:0>�<6u[=N�=ӓ==�{(=\��<|h=:�<Q,�<�=����<X�v<�S�~�@=�#*���I=��6=�\��-���( ���uS<6˼�_=Q`��Y=G�<�"�<�
�<⢐���=n�o=%;Ą��u�<̳་�1��y������Q�<�!i��μ�������Le"=�y����H<��=�t+�j�'��������
p=�낻{K�9%����B<.7f<�c=Yх<[�h<�S�4��:G:{����:�����NJ=s
=7o=8�{<,9e��3=��=�Ti��-q=l�O<c����2��1�:8���t�={8���V8=��ڻ�X�<9B?=�h)=ta� �;	'�<f�n=6T=�u�<BVA�ǀ	��s���<���<\�R(m=���<�R=�[�0=;��o1=�=> J=:������'��إ��A�&Tj=ȞW��N�xH=[�<����cTh=�Tq�b�����<m�U<�����+��w2=�7U=rS������
�;k,<��<Pa�<KAۼ�(��KM����"�A��X<8Uڼ/���o^X;�=�i`<�oC�a$��2�¼�kS��!�=[<;��e=#�i�����=F��0#��B�J�g���4�2�Y��YX=s��<��<��D=G��=�L!=4�[=�1=�:���)��*w��K�;��=m�"=�v=�㒼q��i�:T�;�=|�_��s4<��ۼQ�����=�<ǽU<�u<<�<^�4���:ޏG�����C�<Z&5=cT=\��<$/=���<
���g@��Ǭ������T="T=���< ������`8<�rE<= ��Ę��Y!��6żi�^��i��I�����=�;y�+�B���ܚT���K��/=�
�r����`D<��=Pn
��C��+<��b=�߀=�W�����W�K�8o"�I�׼������;�e��������<����<��m<J>L=z��<Bմ��Z�<��<��M�w^���Z�M�
��*��>���w��@j��+=��w�7D�L`9���&��������<�>=�H�	}��w�x=�]���~�D�=X�W���P=�	A=�oK=��<󢲼䃅�var�x��<t*�7��Pn��|���!��ڼ�gb��?=��_���5=��=`��D���z<C�<�y����<P�<BI�=;�G=�6�O��<?��<���<�t'=�#����>�ð<���<4��<g�=��<�Z�ȑ��(Y�<�T'���!�E�V<��E=f_	��p�<0{�<>���<"�27=���r�.=�%$�#t��{4<=O@�<��ۼ�9#��QU��<<Y�<&,���]=,��'����JV=^��;��h��Q�<1�y��}�;~��Ř�g��.�ϻ����.��p�P=eJ�������<R����7��w$�9Gw<���
"W=I�Ƽ����vR�&n^�����w��aYR�l�:�o� T��(��k��<(3�<M`��ѾE� W6<izK<��K�iݼ�v��8Q��I��rJ�A�u<j[���:/�a%�vpD�s= �<&����	<�7���S<9��<�y��e`��;���<K�м����"�=���;Q��{]��.o<�ɼ69R�<�2=�==�M�;�^=r��f��<JZ=������^=l<�W��~�<h3��
��;ճ��hDJ�3�/�Ӛ�:��ռ�rʼ��<�����w-���#�|��D�7�;�<W��<��	��(�<���@���<��<���v���X<<f2���J=�n༯�V<��<}Ǹ<|?���V�������<<�;�<��Y��T�����l�<��G����&����<��ͼ(�򼲪D=o�켋�=�@f�a�Ƽ�V���\=���<�g=��*�����:�����D=_�U<��"� �#<;�V=�/���<@�<>���C ��t�i�<�8P<�δ<� J<�h������E��'m<�(=��Q<���=��<`}ʼ�Wؼ�����Jp��<��=T��������λ��^9���E_=#��<�����=�����4=件;BQ�<oA�&Q;;@OO=�tǼ�-�<��=j��;��N=��'=E=�%H�`^1;P_K;U('=��ݹ����dѼ��b���#�g=ț;.�+��]<y��_�����\�1�3<�("=��-;?�����y�<x��<jx~�Nf=YՒ��Y��x,=hMj�"�<���;��1���#=�JҼX�="=&;�Cq=�k�;η'=e�`��:h�=<�$�G�A<�i:=��i=���<J��[�<�ϼ�G<=����7o�猺F�p=�~2��ܼٗ<��A���<=ۥ=L�+�V�<JM<Q+�=g�=F�+<����D�6j3=:��\�(=�o=�e���<<~u>�������;I�<����˫�tiJ���<�Ź�b<�j"�<�=�H;ϙ:=Z!= 7��V��t�=o48�ZB�<;�=4��<@�^=O�ϼ�B��Ɩ=��e�#!E��<�xD=�)a��+��?�;�߃���a�!|�<*�<}�����=���:����4=c4=�U9�B�=>�#=:���(=eUT=Z�|;��==!�-�;x��㰾����<�	=�>ze��1_=i�5�k6�9�P������<��{���e�`�8�)�`�^�
�M=�s��Ҥ�=�U»<5#�E��z	=��<�w<��3���<a�<33
�)s ���E=)>-=��n=!�;f_=��T<x��<��>�yAT=8�<X�=%��4A>=�'�<$�Ҽ�=�=	;b�'�ט�����<7E=����#=�9<���9�}�����9<6�޼�n�<}	>�ΰ?=��;�볼l�=�ĕ<`H�<����?"=sGx;TP��ݓ��	=,Ƀ=��<�2�<�V�<�Ř�A4m���9�3��T8��HL����;BB���km<��&�b=��0=6�H��c����;����x��&t�>x<�8�,C�}��;�_2�����-����`�������軎�1�Y_�<0(\�C�f�h��6�I=�Z=I ^=%c=���ƨ=p�� �=��s��m����<dL<eN���#=ps����<�����<�p$=iDD��0=\z<�x��d'� sU=�9u<�F�<�}a=����B�<�r;H/�<�?(=�-��>Q��Cք<K��!��<lLѻaC�<OV��|@V�\��<`.Y���d=g��<��<��B��A��[�	�;O���L�^�4=��=��L�HS= 	=j�'����*����5=�j��\=L�<���<@;�=z�$=�l{�d���?�]�@^/��QE��3��#SC���"�t�S��W��ݜ�����;�'��}p��JҼ�M��R�݁ļ�o�<���<���<�(�<A~W=�)�
�<�&=Q�(����(f:t$=�6�[4P<�Iݻ�;�$�H��K�����<�bX��J���U�>"=�J=$=�< t���/1�����y=�X=Lμ#'��� =庒���d<59����7��v��O���u�<��!�3u2=9C�Ĕ�<�#�< �ܼ6�U;@��<�+�G1=A�G���=���<�(�#��:�p�=.�?=4M<Iя��[e���9�c��<�`�;�~:��;��<0��<uZ��Q�1=y��Q�<����/=�qǼ1=ak�<цU=�<<J�==&d=�n=� ���Pf��iu��>�����~"=�����R>;%_D;m9w<D�o==�<MB�<��=9@���3�ka	=��$�A��z�}\=&�<�}��l��\/=b�>�Fr�Q�;�d�<�� �W�X;憮<!t4<)SC=S1%;�Y輼�8<o�<3�*=Zpf={�b�'�-�����S�$<{��<��G��ڬ<k�!�ͳj=�_A=F輒]�<�tO�v�N�*O6=f6h=v+(�|b�<h,�4O3�@7l=����B�\w#<Ѡ:��@�)St�,(�8Q=Ʀ4�PQ��r~����~��zؼC䅻 �<�%�������м�l����r��&=sX�<&2�A=�$*=[/�Ph�;U�R��<%�D<.�����*=�9<<�tf�k�=\�u=��|�tY=�Kq;�B�v�:=������?�i�Z�1K�=��W=�ӹ<B�<&=h���a��WS����<�P<�M=bc�<��I���S��\(=��8=�5=�@ż��=�d��<��~=��)�V�F�ʁ��֊E='�?��u������9E:��*�<d�om�������,#=�I��>ͻ���L��<S0�<�}�<�zS;�j#<��@���djo�:(�:t���);�8�$�0� �h<�9�;T�@�Q����Pg�;���k�;�����+= �2=v� ��x�Æ!<$P	�}��<��P=����tټu�ޢ��m�-=�t �n]~<i��<�}7<n&���%����B$S��=�;�W�ۓ�<)�c���U����;#������'��:)@|���K��.�<�E�y����Լ�;Z�}�i=���<y�2=Ȝ=��;�A �{�5���A=y$�<�;�r.=����d;b�-=�F� ���<y*t;�<��C<^R��Hl:۱8=:M<��ѻh��<����r$����;�V%<��W=l<+zM<�=��p�0�=����%=lT�ʙ��J̼�3=ѣB=��D������=j���誼�����0=�L^=�w�<=�<G�=i�1=n� �����#nk��')�L�l��<0d<��'�p��c�)=�9 ��������(�<�Mz�,VG��~?��<U�5�_�N�X�=�+��5�<���9d=5=��C=g�x< �%�X<K���<�<�==F:������@��[^=��;�>��Wͷ<�F���a=kb漾���vH��x��`�ˬ(=6����Y6�C�<��<�]0��[S<p�����6e��ҍ��,;="XP=j�=�	!�.�?=���b�t�<��<�q�����<i <ҿԼ��;�>P<�m�;w���8��m�<�L��=��<���< #�<�4���Q=@� ��=25ߺɧ=�� �S&<�U���A���-���"B=��;�=�U��1*=>�;���B�=��Ἓ�ɼ�-(�_��<Ȅ��e=�����	6=*k�<	�D=&‽�}��8��s���1���@=�j=�~�Z�����m�=���$P=�QG=�e�tG�B���dy<zR<��K!���<��}��X=V��f>9��ؼ����,��<+qM��a=@;��x��� W=6���n��:���<��ݴ~���5<��<���<gh<#u5=Ԏ\<o&�=P=��μ %=~0�JO��z����b;�(=�7��P"=#�H=T� �&��p=cp��?q�<^���/�"�<��`��<󙖽�'��5�;=۝�z. =S=��C�� =�A=���<i�h�|p{=�
���l=����"S���<}$��927=Z�ü�+:;}�u=W�;߳˼J"���G=B�ݻ�6���[#=�Y�<"���3TT<}"k=��)=hI��53= Xg��Z�<�*�ΣK=jQg=�=V=#<fΩ�99���fD�*�r���{<��\�u���i=*<�<�%"�f2�WL="@�<�^(w<��H=2�⺏�式�;�a)���=h�5=�T3={�8=�h�<�.�<ãE��9� �"<b��<��|=!�W�k���S<6��/�j=�ȍ<��$��<0��KF��;c��+<�p�;�<o�0�t�<�<��%<�,=���vP�=�#�<�$�<P�<TQ�<�v`<�	��gO�����v�+���ؼ�&�|҈= h�<���U�=��
=���;�f.=M��;�R>=`��I0�:���;�r��ކt=׀�<q9ȼ"�6=�:��6���Ȼ/⼢��<xO ��1���(�����;�鼥=���������FҼA���v=l>(=��#���D�i��<��� �e�,i�*h]�3=�=�wȼV--</C��d!=�o－�W=9^_�m����<p2�;"$!=gU�<>�/�ŝ���=��<�fT=`#=h�^=⿚���'���8���<���<����k�J=`�=a�R=C�;���=y�'�>~��?�f�Է
�u�=
�4�e ��k�R=�xI��	��!>�KR=�Y�a�9Y~�n���3�9��,�����.2`��&=��"1��ʬ/�����!�9���=W��91=xw�T�/=]�����W=�t@=�
J�ы�<�s6=i���Y=aS�<��¼��7<�<�&e=��1���ռG0�&����� �O����n�<@O�<��2=Pϻ��RK=HW?=g�I=�j�;#�=�xq=-�D<�/�<��ڼz�ѻ��Z����J% ;'��x=��9=�Ac=`r�:}��<��<P�S<)��T�<t���=](�+P�ZI;�e���/=Y�v���`��]�<?rB<�<�M��<XJ����̺_ <�5=p���/f=�U<����$r==X��wܻ�D=�<b7�<7����M<=���;������<�U=�h��:N=��=�I �`����<�F|�q^�<.ǂ��	��������~9�0=Vt|=��I;����x�*�=��8=�d(��W?�R�Q=�l
=!0��87�0H�2�<YH��;�=��-=��a="��2ļ'�I=�D���-�H^o��&n�i����x�¨�<�>���N<�h�=je��a=80Լ��m���u<�XR<�3=�����L�=}|�<�U_�m��<�I�E�==u�/=)<ü�[3;���<j{W��,�<�53<�9+=���<$�\�</Q��K=��ڼ!�y�Y,���|o=�#��u+<�*���;���Q�M=)Z��O�C��C.<��2;��=,����<)q�<��ź�~&�#Z<�J#<}<�f�=C�U=bW*=a).=���Õ�m����b=�W�J<FD�<��;<���6r;��T=��u��7���V�L��<��r�4�s�w�S�l�J��i9=��/<y�7=�,�p�[��>��i��J;;��<n��<��@�A�5ˤ�QJI=*ը<�#�?f�<T���g�(=!�'=���L =��[�y�0��5!��t��QvP���p=�;�d@�G����'<B�����*�<�m1��~���Q��8�=rH�<�?��
�=q��̴Q�,f=X� ��e3=W����B<��H��z�<xvR=���<qz=e�=O�?<I@��f���$P<��3=���A��<ux���$�=R4=�:\���7��@a���حC=�>�<�=�{�;����n�<�x<�����<K~=��O�%-��@!=�|=}V���@��0�;Ŗ��\�kl�;Y��<V�<t��<6+�_�,=q�ٺ��7;�$x=1�ݼ��=ih�<hU+<��kR���
��?�<��	=o�`:�v���&����<rݝ<� �K7C=h�k=t�'��HļB��ݼ-8�;1��<j�h��;<)�8�<��O<��-�仔
>�0�6�a=(f��6�!��l��=���<����m��ɱ��D'����:5�j<��\=)�.���hA=Ea=��;=�y|������q��+��*)��-�;�9`��#D=o�Ӽh�<l�3o��yo��h�<�i�<��.����4
�:L1=BM�<�$�� �<��<���bo=��@=�p<�<�d]<���<�l�<X��=>=�	n� ��;��<=��Z���μ���<s�v<�B)=
k�<�D=\��<�=1<��:�aML�M]����<�Dj��5=�6<!=��*���HƻK�<opA��V='�!��n�{��<���<��=zz��iv�q/N=t�u=e�=�]939 <�4�����<�<�W�� ��Gh=,@����<��<�n = ���j��qG�c��=�%��� =��*��F�<�/ۺOD����0��<6��[�I!<.E=�&��ig�P[ʼ=�@�7=�hw=O
�<�*=���<9�����F�ѼUNc;g� ��.���)��g<@\�:�:��*�W}y9��Ua~�����'���w���5;����l�V��;Ӗ�;禐�K�����<nv�
�� o|�A,E�v��<+�g����� �'<Q;=�1=$Ҍ<�=� �;8s=4p<8��m�7=��=�[)�h��<pjm�7�=��.�=~H�C* ='�=L|ݻC��^�Ҽ&�x��c�;���<��'�l�3=��<R=�<���h6=���<MF$=���<@K�| �sPI���� 9�{�<��<�U%�/�Z���r=;��<�B�<P���O�j����;��<N�F;k�缪r�u&�;kT=1�r�b�r
�����|?��y��%r_�۲ռ�;5����?<�x��d�<��������q���4^/����<dq�<��漴�F<\�<��If�
�C�W�'W=�x<�U ��=,�9�u�<��=�/=���<ґ�<�R�<u=5iF=�oe<U6R<�]��h����<Ԡ@=f]�m��:��<]�<z��sk1�0g>��a���22�K��mA�<?r�;��I�'��<{�P=D)W���2����
�L<��@<��E<I��x��<R�C��#x=5Np��?:=>��yq��¼���U��k�<<}G����by�<��F=���jm�6i�^�O����;�
R=��
=8�<4�<lJ���=�R��q=V8b=U�	�_��[8�?�⼐|!��忺2�c�4t= �޻�J#�wZ=�6@�eh��M��@ɼ��5�`;��6�<X�z=YW<�o�C���<EF��n�n�����Jf=�e�<M�.�4��;��2�</?=%�c��:p=�������<��i;AO��T'B�r�=`k�;�:=uy<���<����	�< b-��~���[#=%_4���ȼ���bM&���=u$1=��l�6�n�^;���� s=��J=5� ;3KJ=�@l�󝞼�F�����<�+���Ք��s<c�ܼ�	;�d��b�<?Q=��M���?�I��<�K���kX�*�K;�װ<�<;=z�l=��(��g#��7��x��<��s��A�<v�b��dT="8= �^�qM-==3<��݈ =~�"<�/L��W/<K�<9��<pǼ ���l��PH=f������<��#=sU��ٜ+�{j�
�<��J=-�<n�]<��=���<���Y��<��3�F��P�]��Ģ<���m͋<�"�%����_����zd`�%���Q藻u>;� ��ټ�N^�ϖ=W@����<i]����_���C=��<@����B�O=�Z<9=9��;ea��7!.<�H�;�W��L#u�5K�9�돻��	<~#@=2Jѻ�/^=D�����O����4/=5| �P.=���&sN�c�<@м24�.�5<o��b���(��4��<Z�h=��;������;�M�<o)���p;]�#�1��<�6���z!=>�@=�y<�W=`h=�'��g��>=N�(�,�y�fa�<)�d���ļ�=2��<�:+=�]3=+U=�Qt<g8=�d<�S���k&=�ܬ:QI��08������T�;�F=��a��X;[v�j�Q�@�@=C�Լ�x���=f�+<���]��<=&����2=��Z=�=+�{<�������l�=]m��q#=�S*����;�: �F3������&��w���EW=�bM<���jԼ!�<~�0=�����1&�~Bz���A=�Um<z���>JA�J�:��l=����~�J=���9�B������.c����<h/<�C�;e =`ps=��;=8�];@��<�Tl=+?,=X�U=�z�<��`���F�>���G�<�e�:"lO�~���O��<(p]=aet=t�v��^��^Q�!"�<��
�T	3=���R	=�����E'�π�<��-=��6<+4<��6���\�z�K<~pq=q%Q���A�a}<� (�9�G=Ća��w���%=%�D=��W=�i?�獢����WT=�(����<��e����<���z���;Q�	.����ª<��$�<��h<�O~�v�?�#��;���<J��=��b=�.q��g���7�<+L�� ��<>�<zf!�����?�<�n�</X�=��k\�%�=He�Dڼ�{��0��;�T%<;=s�2���tR �y
=�=�����im�� �792�r� �dN�<��Q=�̾� �H�����B��j޼_������ܒ;���;��m�<��=l��Ս�:c��<�D�;���;�kN�������<���F;����<��g=
k@��ZB=�>=b�6=�S>�9(H��[�<��;����\<�;�;�8��w=���<)�<���<�G=b ��[d��&
��pH=�}ؼY�(�: �<��介IW���<"O�M3�<+.�;�:�<�<�<Z��	�<v�Z����<�;����;���<���<�>��Qo��dӺS�˼��<��L�c9H��<� =S�����<�c�=Y5��	�<��!���ʼ](L;�.'���2:9k�;G}3=:�h=��<�%�;�<����ɺ�s�=��ռj}�g��<L�g=�P�J�a����;��6?=���R�Z=a���c*Z<?��<Æe==�-=`�<k��]wL��XQ�d�o��J4=Bn�;�E=Z�:�[=$�=�V=sJ����O�<����ȯq=�N~<��)<h�U��<6�y�*=NlR�tm�)
=#�6�;��=�A˻��ڻ��L<��*=��(=��X��¼�*���L�=m�����K#��7&��\��	k��<$�<ƍ?�+I��s*��b=���<��H�0�ϼ�J��Z���H<;��;�d�uE����<y&Q=�m�<�׼o�'��v�<N!��d<�o��<کI�1/�;��=D������lh,��@����i=�@[=�n='u�::v�8 L�Tϼ�D�pO�<��=R�K���M=Si=�Ba<�n=E��;��=��	�kI+�%�S�<< �!��1;O����<��/=���/�8�Xc��J�"��5=��<R%-=��5���n�f��<ݐ=�¼� H=V��<.=��M<��.=U�H���=��μ�8+�v�=��;n?=Bg�~�<�s��3�<�-��TL=�}(<�c=k�i=8"�;U:��
���:1��:T)�<���g�1=�Q���f=����$M���b�vW�;�,�A�+=��<��={�N��p�<��u</�<�q=~��[�;.=ُ��y=o�<v=�G(���=b�E��_;��=��\=g�ڼ�̽��PͼGH������a�<8gK=�w����ܼ�K,<h�<��ͼL������O�
�$�_v1�a�0���h<��<Ź�<g���P0=�<��=��$��)���ȼ�I����<g'�	�P=/y	�Z&���JK=�b�\������8�a�'��@�=O�<&�>�k�<���<W߼"��Ъ�{�	�Z�<�M���^=0�<��<\M��7���^�����;��K���R=į��`�=�^=�/��wL=���<�_=R0�|>黪BW���)J��ʴ���y<�{<c�=��v�Y=���R�'Ɔ�ob<��+�Q=�^��r��<�H=Q"=}0�C�h�����~<(Q�<F�� .�S�;J��;�~l�n����|�)e�k-=c �<���6�=�{=�z=�g
<�7=�'�;n)�� μ\��<"��=GB��z=E�}<�@���<k��<��;�s<�1��&�;�9���<�Q���s�<+5M�<�=��&��[4=̴��!3�;a���l��;kD�����ԝ�H��;� =d�{���Q�"�/=�M�Y��פ�z:�<k;�w�U�߃|<>B�<(�{�a:�<+G�<�Fc��O =����_�$��<\�C=�Y���\>< ��mz<��|��9�:�ya��i1=�2O=?c�5n���<�)��O찼{��,f$�*L_:�&���<�?*=q�\�`*=�ȼ��7��=
����)��h��@���N�a�J��ֻ�=ݧ2==��<Ď����,=4
=k9B<y�;X�J�ֲc<�\1<�����<�]W=���=�t��\K<;���R�J��5=K�A�����;LM�<�sQ=nE=~�0=D�<�8K;�ˋ9�\��?(=��G�<[�).���\�5��T�<�k��q��[�L�\<��<�;�px�<7���*<jH<֗˼�QF=����� <�~=Y �<g�8��s�oPU=b�P=�gj=��=�sf�F��<�r#�#�����<R�A=���<���Fk3����<G�6��RU<�<w臼�b����?�<\'i�v�t=���<�at���X=��w�n=�<�e�:�0=�p�v2���a�<�\J<�h<�=2�R�1�՜-�|��vM=eS$=w!ȼ��=�=~"��?���E����)�=a�¼���<x�;��)�$�˻��U�SW0=��n�tU��Y����)�%g�<����[��P��{5=�0�t\4����;{%׼�x<��̼f�<.��������<76�<}j��vA<.�>��<E컺���:��<:-=��=^�=#Q]=}�=�I?;�<o��xoл*H<�=�v��#?�v�[�:;�1&=JAP���=r�t<ݯR�A4����=w"9��K�Ş@�(M"���;��H�ϕ%���q�pD�M��;$�=eX����P;�=(��lH������<�^=��	��f]��M<-X�.)�;��i<#�޼�s��\�<�7^�ݰ#=�.S=ؓU�������}�=-<��#=P: =�l��<�=�L��� �Hh\��<8B-;K�t<��=����<>��<!e��F��y�<C�� �l=θQ=t�&�C0�<?�ڻ��=��$=L�<+�i=k�o��=�_�:}֞�.V=�ɥ;k���"����'� ���=���B';�<=xc����.��2Q=��a��<4�@=/�C�8�X=� ��m9��qs=h��rx=��<�sU<���ga=����gU�a]8ځP�w�/=��~=ۏ^=�K��־�똁<c�W�F�E=M������0�����;����Df(��x2��*�{=\q������.�<?���TT <G�Y=���HY=f"<��4��ǼL=��5�ǜ=�>`�f�� |��QA;̼<����&=\����R�9N<����;�'�Pv�0���a�u+,=���㷝���c�����6B=� �Ճ<��_=��,=ޗ�k�e��ǖ�W=c�<!"��	���3�u,p�};�<tAu�� =�N����uee<�9d<�e���g<�����$ݼ.���I�=!�����_=	�v�%��'�z=��3=Ē]�6D�<ͅ0���;�fa�>�d�h��<e�F=$16=?�;sq��?dļ��<�:�<�������<��^�#=��0<O�
=�d=��P�(����4=0��<z)U����<yP3=J��?��#�<t1H��`W�D��C(x<��2Lg�.�.���=��0�G=@^V��jP��&P<� "�p��<PP�ϙb=0U���s=��{;���4\=��ɻڵ9=�Ƽ:�d��^<��5<m�=���(6��=}�=(A=�<�C޺1��<dx��ֺ<�e;��S�<I
��
=܉���Ί�߮ü2��k"��T��L�S=�p=wM7�_7�e�<`�i�]U7<�N��@V��t�<*9Ѽ��Q=��,�}"���<K���DLB=��?<���<7:%=�
=�>�<2(�;=���!=�|l�P]@=����c&���:��ssL=9�˼���<�!W<(�N���=��R=�4l=�"d���һ�=(�� &���=y]}���=
��m�p��2=~�=l�.��7'�z�<:-=�=O���U��u�ݼR�4:��s��Y*=1 ��y�R���Z=��==��_T�uK/=��8=���<�Y��6���#�
���@�.0':��<p�p=���<<-=&Rn=oGϼ���<��d�N�1</p<<�jL�IL-=�hG�5u�<
�+�Ɵ�m��<~!=V�<R��h=��<��k�H=\/���ݻaR=O�ܼ���*!=�r=*��<�\�P�<�!��<=�=�@�<�?=v��{�c=�����<~��)��Xq�S}�<0���n��q�a���U=�.�ѽ<ń6=��!���7��9=w߼<~i9�)|Q={ƛ�a�� n�����H=�T=,�=hb=�J<�K���k���<8���W=�uԼ|�����<��=S=7<咩<T�k���>���N� �.=sD����<[m�</��g�/<�f�����w��(Wd���Z�4=�JM=r�	=	��$������r9Ӽ��u<q�y;��<�c]�x�E=(���/��
<�t�mh@=�8=�$�����;�X�&v}=ٹ5=��7<�[�<�����<0ûD�=G��p�;;ca�<W(�<��~�,=��G�
�G�Nf��YT�J/��b=Wm`=?i�<�E�#�<��=�ɼ:Z;��*����<�>�;_D=��T��N<��=~�Y���*�O��MW�<k^��s�c�\��׸����=��<�5=��9����<���%<�eN=��{=�o��.��N�9�B���28�8�<�~�<�������˼��!=�� =SyJ��.�h�º������B�LR���C�:�-_<����y�e=9=�Jk�`����d�Q�<�9
=��û ���(F�!�J�qX���=np<��V��%�
y=&�T���Z=�0l�>붼2�̼T�)����<���<�œ��~<=v�j�����|]=��K�w��%@O�D?=�p�B�4����<����P5��x=����r�=◘�<)���=�ζ�)�U<�*��O=���<�?<��J��R-=��m��~2=� =}=Áܼ���aB<qz�<W�~=Ձ���"5=��S<��<u�>��J�ɔX���4�#�����'�ټKh%=d
 =%?
�	�l=�!��T��*'�iz����<�Q�L���:6�< H'���V�����Iz�ǥ��0�A=�|��cǐ<�D�\�#=��v�k�<��L���=��������j�<��<e�<1V�w�~<m(�<g3=.u ����<�cؼ/� <!
C���]�L�<�2;=�� ��I<��<�HFu�[8�<!f�;4�o�!-��;+� �T%��a,<e���x<�t��j@={�=������&�);e�"=:V�<� A���<߹<u�=�H=�U�6���Z�;��&=~����'��<G�C=c<h��[r=���;!�R=���<,�<�_j���=���<�~���jM=ʽҺ�s��E[<e����Fs��#�<�cQ�CbT�Áּa�-#%<o.>���Z<�5;���g<�?%;
jg�$���F�:=�et<��:0[=�&<J�9��Mu�U[ =H/��)ɼ�g�e�A��	#�oq�<:�h<>r��d�<��W��.�<?�������t'��R���Ld=��E<���qT˼��$;Z��d�=qF=˦����UD=��<Jmn=D���� ��Q�}A=�❼�@�� 4�<�?=I[,���<�1i���Vf)�Ȃ<;4�F<Y/�-	�k����W��E[<a�i�s�<�Y+���b�����e����A=��<��<}>N=�H�:��ļ��;A8�<�~�8�a<o=�֠<�eT��,\���<�I�,�<��<�!�<o�,��K�<�ϸ��V=������^=ۧ�� T=?�=}Qj;�G�|0�b/=g�i<�4�< H���ŵ��y��==��)����g�<�'�-!�TE�;��<����ļ��8�O�=?f"=2!�<)!�:���vڭ<p���{�I������9��᛺����
=�s'<�$���(=�v��)mɼAM��w�;@Y�.��<K�=���=I��:�^��D���*=8�W�Ԣ˼£<D2d;|�g;��μh�<�o��V�<�~�[*H:��+=�D=��v=l9�<מ{=�����<6�ؼ�͏�I	=��3�@+�=7KF=~��<�f�;�Y(=n�#���#=5B��{�<��;A`�l��<Vo+���<wMd<�������u�:�_3=�+=N�=-��<도��)��#��<��%=l�2=�l@��7X�"�<8N��c�2=QE�<T\8�H+~���ټ;��>�.=�W	=��v��P=8b;�ۉ;7�J�8���<r=`s#<�^�:h�����<��?=��I(k=�c�;d�R���;Tg��Ob��*=�aS=�=W=<��=��5�o��:�V���uE�-}�;7Q���=�Jh=y^�|��nt�����<��1=��&����l=3V9�?�s�ZG<Ҷ=x����r;�?�<Ou?=�Q$<��<��5��6�UN�<��-��6n�<��={_�9��1=F�.=c��~�����N;|4��4����p�<4�ƼU��<�7���ռ�9�T��=�|�;W(��k�;	ȫ��Cʼ��=:1��Re��q=�M=|�5=@��<c_d=�u<b_���a:��J}��<=�"=�
ؼ���<zdt=��&=�q=�3D��Z�;j�&�v�/�
IK=b�$<�7F�ې^�^2�<�z�x|�M�J=��5�������n=)Hi�3�o=#� �[Z=�Da=1T�<���;��j��n	�DZ�<<�d=�F��@��3������%=_3H���V��?�<!4�0(�:8A<�.�<��=3�t�j�
K����<x��P>=�~�<:�`���x�{�2=��Q�<k��<�\]��9=��=N	��U�:<�c<>�<.��<V1��,�Ӽ;#w<0 �)�<1�8<��:=I�=o�/=���+��;z��CL=��<�<�y���H*� ���׻�RM��vO���Ɲ�<��<ՠ�<�����;�E3�����+Xr�+l=��=8z��2�K<U'=�����,<˿4=��!�K��<��=:ɣ<*g=��t=$O�x�ۼy��<PB:=꥿��a���_=|	[�"�ͼ�F��7��g*�y�<~��<��+;�_G�j�}`�<0\����Y�Y[�u=�"��<��P�K;���<_S=��K=����܋�<��
���A�6"�)ea�u�Y�/++��F��<�Y�<��{<R�8�*�=� ��l]!=�w��Ǎ3=]h�Pu4��L��,/=S
=�������<��<�7=�:"���E=]��@��O�;�{�:��</���ɫ <5��G��<1A���M����<-��<��=r���_��<�(��!�#�<��+�m
 =7�<򧀼 �M�m-<�� ɹ��t�9X���r=�ؐ�6�<��6< pR�J!<�1b=��<FܼEi�<�O�<�G=_cռ<�J=��^:�g=�B!�buk��==�*;!a�<��
�,�+��g=Q��<�켺

�F�C=�;�e==�ʠ�
��[V)=�sٺe���R�<W�=�j|��{<���p�p��8k��\ټh��<͍�<��=[�<<j��Q^� Bt<"���K=25@��s>=��=P�?=�<�d���K�<��$=�n<�,5=�f���o�:�9��F뙼�H�]��<�3�<5���Ռ<ޑ=]?��F�<XNG�:�=c�%=���<%��䟼��[����;�:��L;˄�����{&<��^<�^�.��<��Q=L�=F���?E�뭡<�,<:�<Q=g�<�};m�.�]eI��o<?j=K�<{�"�M�6=U�7�Ͷ��m5=�i�<ͤؼ�(뼘?m=�����f=5��<�Y�<I��<!���}��)�/���r�Ҹ<��.��[`�.b�=<#�N��&l/=
m�!2�O'��2�;��A(<x�]��JI=�˻;�};=�;k���;1��;�s�6�,{�<��Q=u�p�x�&ȇ=�lQ���=��6��_V���<_�&��qW��@��ͻ�^�O=j=;?�=;=���;u)<=�m3=�ۄ;���<�8��j=b}ּ��X�<b�: "=�yb=7���w=c�Z=��������)	���i>=�	E<Kp#=H�F�Ἕ���E�7=Z����L=��c��'�<���<�� =̨�XO�:MI��Hɼ�|��?�5��,]�H	�<)8��1z<r����@�N��<�<~v�<,D=���<C�׼-�E��e�;����#(=b]1<L_w<F�AF(;�� ��{
=��<�Rb=V��V�j�A=���<�G�0´:�*�<��D���<ݹ2=�=��<���<�vh<3m�x��<�5Z<xO><��S������w]<��=��<3<�ri;s-T�,�k��.9=_�(:#<�=n�E���5-B=_h�+X�<�����L2=k�}�3�<�P��K�����j=O�%<��=U�%��`�;T7= ��<q��;}�\=���;`~�<!����)���ӻE�e��V-��f6=�A���=�4����F=�}�<����Dz�;���<��<��=0�	=����ѳ�cf=uĈ�ǜ�<�V�ci=�B=I��:ħ������J�<�w�<n��l����5;�������<�.�u�-=���<G�'���=�͜<A�Z�\�E=+�;��dn=]O=�&d=�P=�y=n��<E�':�:K�(<N$ �p����<��<ݭ�&̼�<f�<+K�:w�=�a<�hg<���<�i�<cV=�ā�:�����sJR�H����4<K�< �<i!o<�[�<k�»KP��kP=�=���E/<�/�Ȅ�;t��<p�F=�-1=��;�l=e�+����)���߼�=��%��y�=׿�;;��;����Zy=�b���@;='4��u��j�<�q	=���R@:�n6<�'I=k�^;։�<�K�<<�A�~�7~^��<��B���<�~�����<Ѹ<�e��̦滍�<=���:/�a<Q���< s���a���<�L�c���PZ\<��B�f.}<�\��FF��&���U=�L��9=ɔ���T�#�=$�`��`	=o�,��/���|�`[�<��i��w�;.ͼ0�@�Dꉼ�,���.ʼP�˼\#��xQ=r�����=O#�<aa��]����;���<x�#�=��<Aǘ<b�P���$�h\&��&��B�<�'3���T���<��<<7�<^%N=�\A��?�G��kZ���ݼ:����+<�bO�-�;ۨ�<�1�<���<?�,�$2��0�_�h:5<�)���C�ً=�p�� =Qe=C�ݼJ���O�<�%F<ڗػ幺�~�Fp�J�<N������ ��$T�_1U�� =!�(��D;��傻*¯<��=��<��;��'���;�={�4=�'���b=Gb�<X���F`H=1�;<So�qC<M-�|~_=�(s=�ҁ�R�T=��k;�?��7=X�A=��/�,qp���<�`=%���<��X�P&1���M��'<�].��O��*�<v�K=�7=���;�hL�!�h�DQ��&�ݻJ��<gC�<�x���:Ya`�&-���ǆ<�ϼ=�<C����<���<��2=�A�
!�;�w�Z�<�I��< �'=K�M?�;�;��	�O�-=F�<�M$=��k�հ�9{�%;��/<Gl��|������A}H:�H�Y�:;n�T�a[�<N�/=y�L<����/�a<qI�I�h=��ּ��;���;gė��.�<�C<4��5�C=�;��Y��<uL5��]�$�b����<;[�;��<Ωv=c�*��g0��<��ܼ+=C<4;�<�S===��8<s��4�����on<�t=?4M�ؽ=���I0<l	=����$#;�����2�h�?�OJT�D�L�/)ټ��y�A���<S�0�>�=�6<=�mp=.�W=�����׀��I=��f;P:=���T�$;u=)⻖�==>�k��:=W�<�>=�[[=��	�i�H;I�<T��ɝ���C�1��g�t���<{�=�\�I�	g�;�m[�$9�<�
=�X =�细��\͝��O!��� <��X��\Y��m=d���@<�b$=)��<Y���T
=�r?��3��k˼lR�<`Qۼ,��Z�c����<�n<�p=�������<I!<�ƅ=�X`���&;�Ԁ��R=�T]�=��9)����R�V.r=9�l<�\��<�~	=��b��NL��n=;(%���;��1�޴�; 嶼�g���U��<}hm=�\#���<��k�/�x�ɮ��&�
<s<���輂Xa=�!K;toI�H��<�O��׌=O~��E��A�#=�]�5�_<֜i=��߼��<H�W<'S�;^�n���<�X��3ܻr[�:��&��3<��4�sa�;�����F�@�<u�V�W��7�<I9��z@�<W6��B��b}�<K�w���9�B�w��iT<I1�6��s<k#��+��*cԼ,`�;���^��)7=�l"=9�]=��JO=�����M���;[R���J[<N1B�z�����.<v���7iL<1���%��1Y=#�/�x݈����������#��}�)=U�<a��<�q��F�
���cD��T#=ZP=C\=b �<0`C����<���;`P�<N	���Q�����<��=�����&y���wR�༦����]<�;^��<U�=Cj<��<�J�ʂ=���;aX=��������V�)y��qo�ЦY��(ۼ���{�<�<�r+=�[�;Yk���:=�#<X�<Ȏ�<{]=�Iu����@��y=0n�9<�=��~�NkU=�K=[�!<�J�:��<ٷ;�h���-;	�)���<�;���+=?���̼�B༵Հ���<�x�;��=����<��?=�V�Q�H=��'���=w|�}�-�<P鼽o���߇:��λP_���:���ռ��[i;�#���;��6<�[ۼۼ;=2=���=E��ѝK����<��L=���;I1=,��<ӓ!��/Q��#�����|b<�d*<Gd�=�,��(�a��<�f=Y_��㹤9�鋼�	��so=g�H=�)�;>9~���<{���b�Q<��q�f�#<�&���E\�� 7�<r�u����<�\�<e\������X=���=wE7�¢�oM6=E��ٞ6=i���t�
=��;='���/K�H+ ���,�⨻<��,��:Iy��:1�<���<�.O���)���`=�ݮ<�== =K�#l<W=#ʼ�Oͺl���>=�9<�iX��s	=��'�s���ټdN%��^��V�<O���U�n�)�G��;/�p=�a=�d�sO�� 3K=��`�Eg��������[��^<=S�1�^��@D=�l$�%�<���<��X=V����ѼZpt�s;\u;�U�ɻUQ[��.>=�Z=�Hv�h]�;Շ����S�c�ԼT���A=l�<c�^;�C���q˼wzy�a�л�� �ho���? =1�.=޾�<*��<� =9���d�2߻�:�G��P���HaܼI��<�o<��طc�8a�x��m����2���`���x=�=؃��*��ފ���)w�[a�������w�%�D=EϿ<�C�:rc���&0��=l�]格L=ʘ<�ɯ;�ϧ<'�
�>���~�޼��<�,9=L��Bi=����?�<�@�<���9�B=�-�~Wʼ<1�<>T� g$�C$;;;��&��[=k(=�\�<}�<ڙ0<���0�@��f<���:j�[=��`=�����g���;��<߅�<H����G=�,�m���=1�c=�{=F�7=x=A�=�B��.�1=+������<7��A=��<>>�=��<�*=���<���<��]�.�7�}�:IVڼ�5���A�D>�<q�U�"�S=���<�u���S�=<Le={��<��;���<�k��V=� r=��[�N��<9�L��V��T@�H�H=�]�<�[�Яt�e��e� =J��<��ݻ)=^���{=Vk�<��<E�<W�<�웽��a=,�R<�]P=0�{�pTۼ�n
�=,�[6�;�˔��ض<:�<Vt����;<�<��<�v%�K\�<��L=�=?���-L�;U�ѼǩѼ���<�
�l�:��x�)A!=�QJ�Np%<��	=�6'� ��<;�=4��a>/=1�#=�8#����<۳��A�b�<r�Ǽ:��^A=�7�<�r_�O�c=��[<d���|;<����h5<��"��C�;zԎ<Y�;=Qm��L�n�B=f,)��J���c8'�<�����k=�$ڼ��	�y��=��ؼjP�<�5����]�����;��0=W==2�9=Wj����<����k5�o�2��i=^�B=^�軮ɦ<�Oc=��&<��<��q�6!��%"��Fe<�/Ἠ��yCK��8?���
<J�n�Z��R�ZL�<3�)=�"��t*=�6���7<vli�~ۈ�8�B�j�H���>�H�t<p!�<�6�<����e�䊅�7��R헽80A�)ѱ<�ǳ���4��C�<�D<a=���=��:���.�>�j=*�B;&H=Ɩ�<%{a<�K=v�I=��;=-�	=G��xh��ab�G�e��[］�)=v�\�`�ҼB~�q�<��=S[=�Q=0Ә<�=�LL=�(���=g���B<�r�u�a=ߚ�c���Z0<���<9:�<l:����e��U�<0����ѻ��P���X�?h��x�(�5�ӻL2���IT���=�"�<91`�o/�J����O��u��D2��dW�k�ü�<���
m�=K��1��;[F
�}��o<m�=���p=V�,=;���9
c���5��e�����:��d=�i �wPb=����Q7|<�X+��b=C=zq=�8�<fG:=��=
d�<��D=��,=Ջ�<���X��<�h�r�(=C�[<r�=b�i=��<����)�'�9�G�N���
#��H�<�=Mdƻ��|=�$��t� ���x;gH�N=:=S�:=geC=��-��}��Y;��������+<�؈�x��<�8�\\���D"=�A��3=��G=� �<��N�~V=�h�<&$!=gk�<�;3��<^���mz��pt�m��!�<9=Vrż!勼4���t��@-=|M�<�Y<�=I�1<s�8=DT!�'�<��<�&���=��.=뵢�=l�m�Y�W�n=�i=��Q;Ax�O)��tԼد���2��c�<��|<�h9<7s=Ӣ<���<�P=N�D<yK$=\C>�d��J�=QC<v�>=�Ǽ������72b=e�O=�7=T|�<� �<���<�� �&�伢X�<���;c��<��&�Y���N˂=��Q�&����7�=3��<��8���<Y�,�Q�<��x=?F�<
�x<�f\=i[�<��ּ��Z��U=[=����1�<��b(�<�};�(��[��;I�<����<�;K�ֻ�O)������.��㼋�(<�N;�<�T���7<<�x�eT=��i���
<�J����,g<�:�<���<�3��ŋ�����*�=P�N�S9��<�#���;=�#]=�b�<̎t�+��Myռy���J�9==�4�n�(�ԫ-=�j�<*^,=�3���=}>�B�=6��<fǤ��<{7;�h=�֡��wB=<x1=�0=��Z=���<��<��5="��6*)����9�S�����;U��;n*�<�o(=?�+]];�Վ=Kp);ֺg���
=�.:8�Ǽ0k=��M�N�<l[�<{_��a<��+ =��X=�i=�g6�ۄ����8<{�<m/=��t�=�C;h;=�2�9�d��r�2����;��'��[�;�	6=�D7�ԭ�<#6<�����\�9e=���=WR��-���@���<��/�k5)���=�k�#܅�~8g�������<<�qj=�L����<�v�=�����=o㵸�bY=0���<Њ<�7=缅<SGG<H�Լڌe�Mz޼՟)���;|WQ�$:ۼix=Q��<�6]=j�;��=����9��&��x*�m=+��1<M��:���XH<�����Q=��<oy+��`.��	���j�<�A=������;i7= ���Y�<8]E=<������k+=�nV�����ټL("�,+$��"=�����A=�a>���r�$���<}��:���<��d�W�=�S�<�	 =����J�K�(���0��9��3X��ݲ��U^=�<�EL��LA=[/S=�/^=�|w=@)��:����i��䬚���;;k`Y��B%=�><�i<cvV��yP=��J�vK"�ϾH�����2$<W�=cQ=��p=d�;��=�v漑�-=�p�<ᾨ�W0���,����<7�;..=e�0�d��د�<N�\;$�=Oӿ<T!�;IS<v����<W�1=�p�d�<�=���<����v	]�Wf,��]t�4���̦<����4��u='�y�M�H=��=��0�7E?=�Vq��2��*�<��w<K��퉖<�&�Ϸ�<ż����촅�2�<ju�<��<�I=@���q2�`�B<�ٴ<(#=��r�o���W<&�!=���=K��<g�,=��d�`�=W1�������<*<
��<k4�͉&=�j6=7�0�7�к�G�<�|)=Q!����]B��w�c<�/T<��<�@���u�<t0�<ϛ1;y�=�y��*�;���|%��5����<����s4�ca����=�\�}��m =n��<m��p6�<�x5��R=��3=D�ݼeqݼ��0���=�-��UU�<�Ԑ��������<:�i<pro��l=حݼ�x>=�"����G��h�;���G�w=�eD�8����1��T�\�<&:P=3m�<��=�=�<�U�;���<��=;F=�Q;��[�=7;�`�B=�PU=�4���A=�N=��Ѽ���<�,=UN5=� q;}�;-��p�5���;�=����"�<������;~3~=o��<�o	�]��ȃF=����	���/����< `�<l�=��������~��;h�`�#:<�c��|�;�4<��Իb�{�^5��0�Dh-���!<�9��=�7ܼ�k����/<�NB��CQ��l=E-�<�<.ǌ<A�˺H�<�i�o ���i�/������M=p�ؼ_������<���rd��1��<n�;�B=a�k=goi�d$1�w����5=G5=�=uq]=OB�λN=T�;��ǻV^���;+��A߯�
���%�4���>��mi=��I�8������Lh=|t,�k�<��^�OKA�\8�<®��	{����;+���yf���P�kY��Ŏ:Ӏ+=YO�v2�<�N��H�x������/�;�b�\=;�=@��ux=A�:FZ=���;=��<G�'=P<ֻ�_	�����%Y�<6:���X=<<ϼ�_%<��׼Jɲ�G���uW���<V!=�����uI�:n<���<Q����<S1<P����|����<V=�<i9S�3"�;:0����=b��0��<)���G�a<6�=Oh	����<J�Z<$V��xN<�#U� ��!�H����R��<(F9=\nӼ'g���==U4;=��i=��b���<[!W��A��;�V�����<�O�c�W=}�L=L�=�~��1氼��F�>��Z#$�2�`��q%;�L�<X�&=����C�n<=׼�ꐼu:W����~��<<��;��b=�\=&�<�4�<�|�<��C=<C�;��*�)=�=��<T�=�zϼ3~�=?L=_��<k��!p�l�O=,f8�ҳ����<rp����&��8N=%rA���<�$=(
�<1=��t�<���;)�V���ȼ��=�w#=�M�< ~9����UU�U	 ����:�<����f��Y����.;;N �s:<�'<7R�}؎�ԨѼ���<��U;.W2<��Z=no`�A?,=q+H�9>�:��<�m��UB���=g�=�5Źd���a �ݾ*�X�)��kA�N�<�J�NC1=�(<=Ѻ��I��K���<��E<��
lP�%r���2Ǽ��K����<q����zl=2����[�<�I��
�#�<�[��}h���~�M9=��$=�����O=Q.�W��2<y#!=�o�3�=�Z;�;ü� J���L=>5=�?<�<�;Ʈ`��[U���E=i�-�t~ͼ���7�;)>8����6����Z�`=��"=��U���p=�h�<�J�y���H�W�S¼�-�<6=�=Qby=zj"=vbu;d&�.#����BT��>�¤��@9��༼��;�N��$�<��漐TK�� ��"�<{��Z���^�<�����R>����<�a��!=܃�<Xʟ;f"��덼C�1�o�,�=XD=_-=F�ռ^�<�j�����:��8F��?Z�jGc��]�A��<=��7����3=i��<��	=�XQ=.�2;��<��]� <��<�q�<7���;�1�<*[�-�Y��(R��(<ȡ;�M�<�"�U�<�����;�Ig:�B伀�g=K�5��'<=L����m㪼�~<5��	<�Ѧ��iF��{P=�ȴ��o���6��A�c�<_��m�%����<�����c�$�V�]n=�-���K=	"`��'�<� J=¤=u[����J�=�M���=�k�; ���UK��u2��P@�*|R�W*=Հ�
��z���P��=�՛<�k=����5�_*=B"�<�á��)��D���^���5���:��j=wB���"�<����eD=-)μ�DO�&�Y=8�&=ƹ=�m�:���zoU�dun=1/<��� &(��<�{�P!=:�+=T�;�m/�HӼ�e�<�y=�T�/���{�N�����t==�6=�J<Yp=���yF�<�|ڼW�WT�;�d��N<���<R��;&��0�6=.%<Ka0=%N;�S��=  ���&���S�K�#=]�;֖�=�+=V�<��<�H�����a=+�G=Ųz�Jʼ�,=���e�<$��'pj����v����z�;�������Y)w=)�A=�,��Q#;� S<�Q�<���<������<��<�r�����Ba=��ҿ�<K�::a��z�o��Ï�##,=;p��Q׼�k=����hq��PS<g��<�1=r+�}��	�ݼη��ա=����7=(n�3���m�ؗ=l�\�!^7=9�>�-=������<ڴļ5�G=��r;!?��{X�+�2<W��<:���~[����p�9��	����ŻY��l�#<�����K=�䱼B�'���;�m���O=�@��v$;�=���<)B�+v<��<��{����C�3�<��H<_�=9�g=
�r<!�P����;\/�<���<�6�݈8<��;����o-���=ct=��=_�m=�J���0�(�A<�C�2�Ƽlư<�},�;�8=�=d.�<�c��h=�`=!�d�*𝼚N�T;Ġ��(<�������w�Q��μc���`�<�6�.�q�hJ)=��=��<����fe�:��=7$>=�5�<�]1�A<;I�e�����=uἹ�(=v&��n�=�����đ���y�k�3=���;
��ȇ<_�%�i.=Q��<ɔ2���ܼՂ��!<dJ\=��<�[�<,t3=�S�t�$<�1��3A���5(<<m��fk=z�;�`<����~>��xμ;h�{����=��<
�z����<:)<��<�;�"�:��4=�Ɂ<�kg;]@=N�G�覌��X��. Y=Q�=���<�;�T����	�B�0��z�;�2�Nz=2Q%=�`�!GQ=CZL���=�l�;��>��w�;Y��<�F�<V\)=�E==c�;����U��	=�I=)�� �;R�;|��$<1J�<�R�<�	(;c��;�Uܺ���MJ= W4���μL��I��;%��<Q^�� ��<�0@�����ջiC<�C/=<v =�8|����<��u�g�=�dB=��t��^=�D���߼("�������ּ<�\�7��uλ�}ּ)�?�+�=�ģ<\ *=�y6��@O���;�Ʉ�:z;��g<�&=BbV=xqP��$e==�-�Wz��V��5s��U�$F�<�+ʼ{*m�a��KqI=�U�<π���c�K��5�<^.=���=?��>��y=4g�:2�H�ڣl<��(��6�Ĳ�<c�8=,5��=�Q\<�=�0O� ��<sÏ=`�4�
�+����<4R�<�n�=5O�]lQ=�m�$/=�v��޼�f�<�x��Δ��ۊ�v�.;�Ǆ�f�<�2�R�Q�m�f����<��`�'VW�w���7���0�_n�<�b;�h��rWv<����1E�=rM��}�����<3m.=�^� �O�2=hZU���$�Z+F=��@��:�($��w�;A���L=��=ȉ�d+A��'=���9�8�N烼��*:"�ջ�9��]<�囊=��R��kN�
3=���n��<F�=.�#���)=�b�=��<W��5�}��L=�G��I6�[@ͼ���<�<d=�^=��
;�I�: �W;k��<������Z=��t�U��m=;>�=6ʊ��o\��C���pL=b�h<�U �\��<as���j��́������c�<�S��!<��ԼV(�<��`=��M�W�YmD<@�<h�G=������������={N6=��<��D��ռ3�]��J@=�.���,/�Y�:K'�Qv�<���O|c���s=������=��ߕ�q������&=A�g�&qh��3-;5�=���K=�!����i<�[=�1ɼ�I�<.Bd���i=#��cS�;2<M=�^X�j�μbW
�t��<�m»ݳ��7x	=�v~=�J8;4�,<�<���<g=+��p=���<���;��o���[��)|�8�V=���=��<;$�̄�<0%Z=d�<�,����ӻ�>C��L<(�)=�9�t�=�)l=aY<���;��,���\<���;��ϼ.؍�1���ͨw�'�=��Z�\�<UT,<nP<Ty=�/k=�Ƅ�s(�ϛ���NG�y�9g=)T<d<��1�zYK=��*=v��=L)�G�=�'��*=9H�8�e�y�="I���+ʼ������Z=	�Y���0=��M<�@=�>$=�G	��P����<~�<��=��M�v��<���<M�<=~�d��b6<����=o�<��<�")�G��Ph,=�u(=�a=]��<�=��2�M;i�Oc����<�g��d
J=��=W��<>�*=�5s����<d����
<B��<~���%�A�{�����z�f"&��8��h=is~=�W9=�ZP�n�j�{�w;������<	�E��t�<&�X��̼Â�EL0�b�,={^:=܃�<H�ļ��<4��n' <��R=�%`<�I+=q����3;*�c�^�z=5L����p=�>�<-�<@+k�F�@=�� ���;���<��3=���flμ����3� �c�!<�ߊ==%=a,��R�<�Z���R=���F�p=���.�Ӽp=6}=�QǼ�E��D.n�3�<�xX��\=;A=���0=5����|�f���U�<:Y�r�=+��=��oU���{n�v�W=���<ؒ	��:�<�=�K�����V<)�<O�j�7)��CԼ�D�<� L��[y=� �<�F���s;�4<a��<§<g�a�7M��Oq�_8;�0�<0?@�:�>=��H�[9�ҍ��0=H;(=:��< 1U���!����*��Q�<ZkJ��\��:�^�i<�'<�ЄS<�#�5�=����,�����<��/��W<�1'��ҩ�D�m;�2g=L�<��H<zC���j==[=;g��e�{a�<���<b��Ŋ+=��H=��<�,E�G:�[��<�O�<�pS���V=�ü��Q�@	=�ɼ�0<�ut<^�9=s	<��J���x�<��O=�E�rV��a�<���<��;A`*=�)D<�E<=_yP=��`���%=@O=X��Γ=Tm(<�E�ʇ;����V��MZ=���8N���#<���ZS|���=�=s:=�����Fjּ���d=�yA�03=2�����e=0l�3K��*i��_=ڀ��@��U=�J���I=�2&�����:����\=��S<�!ռ��<:R�d	����p�q=l�<gZ=5=ֹ���N=i<;o<߃��!]���r���q��;��;�;�6���;��s��;�䴼�G�c|�<��<�[�@D��>Z�%$\���2�K9��<�6=AoX�Β9���9�����*�6���.=g��<à;�������<w8�Ţ��<y��;=�o�;�LA�S� =(�=�V�<�f=�*`=�*�4pۼP� ���I��<x �<n��;��=�I_������Rk���F=t]=4i�;8�)���9�A�a=#���� ������<u06� �J�I=?/f<qSͼ�;�3�̼��:�9���Q=��	=�%��["��5��D>:,T����<=�����h|.<��`=��|;ǖ�o~;=�]��C���l������d=��<�;���w��Լ��(�9��I���A<�BR���_�<��*��6<��<d3�����<�{=�#�;Q�<^]h��&��F9��L��v��=2��#`=r�s=��<ݤ!=�D@=�s�<���<�=��?=!Sz=6Ƽ�PO<������ͼ�f'=�$�Kg��	)<�W=��ɣ<q=L/����x��X\��v.�0Kּ�5�͸�,芽j�<���]%=r�5=HA=݄���=�Z=3�<�1�#�	=�=@�ỡP�t.�<q�ļ��0=t �:�y�qμB`=�ֶ�L�P=�$�֬J��Yt�ձ�z��<��Y�����=�>0�<����:�<E����xE<}p��Ni�GD��-���U:�L�<����R=��H�P�=�"�y��;��������@��Vw���r�?�=��@;w���W���M=�����&=�0	=�(O�2M=0(;�|�<X��<&zG<��k=������<�=d��=�;чY����<wM<x8�<��I�6��<�+���J=�L�$���;��mQE�c�s=�`��t;o�=uA���I���>=�}�r�<,卺Pb��I��;�[^�	D���T���=��A<+�p��6M�1�-��LԼ��L�����n2<��:�]��kj�E毻�u=~�w��L�������=�d�=^�O=5_=r��<ܘ�<G�ڼ��j=�����}�.���l"�s`ü�O=a�/��M$��/^��c�9:=<�L=D��<�ΐ��6�E5����<�=�~s�����<d=�=����"����v�.�;���i�=�����-��-��N;>q��J�9{���v=�7��x �y�+�S0=�v��b&=���w;�%u=e<����X:�C8�L�h=��S=���_<=�����2���<��`=��P=�M=0j-=c�l���6=7V=A:��M���7��E�\�c�K=
������;��|��T<k#a���<�e�=�<�땼�S3��u1���&=��<��y����[�*�T�����B\=x�����z=�2G=JC[=fVL=:� �D̻1� �-6"�Ii=��@��ػB8=*�a=�:O�Ra9��_�;/-��j����=��2<��<�<{� =1m^�ĝ=�K�����<:��6�<<Dz=�7n�+)�^E4<�Py<��I<i=Y =5e��c���4 =��=4�B�~O=���e<��!������9=���1�ݼ<�';�W<y�<u=��<:���=m"�&�5=4=�<�=K��b:� ��<2O���,��U�;�)��������Y=��=X��<=X�<�4=wS=�v�<����/�"=�9P=n�>=���<JmL� u<�QM��!=
B$��M@;�8�=B'�=�:��;����^�?=�?�<�f���r�d�=(]��<~�}V�<D���n�5|q�� �3�#=<ȼ'':���=�0��� ���wO���;�F&���o$=Q?���<~D�<X;E=������<ݢ��ػ���;F��:]����!�@i �%��,#=ua���S3�rW�9*�C<��<}��N>�hm/:	5<	}�=�KO���6=��<�R�'�/�P=\��;Z�D<�Gż�훺[�Ҽ���<��k<�8�;�nC=>v�:�\ =X���ѷ�<���������!=>=���8Κ���&�ɉ=��=�bp<�6�	���kA�0 =X=����<����<]9)=1�M;��+<a�꼮�=��&�E��Xz=�CQ=T%?;h�<�pW� �m����\�<ckT�/='�<Z3;W�T=��C=�=ļi��<t���9��<$>N=g�2���?��� �/�<)�V�,q�|�	i�t�d�b޼^=����%�?��T������~I�y��<�"P<Pt$<Ea�;<TV=a�M��=ꗻ�3<?�6<�^c=� ��0������'�E��4��x�:\=��<E�!��-��#�%��<y,G=ٖ<�+���(=񀁼�A='��<Cڻȸ�<�'c<��0={�@�#���=�T��cڻ�b�~=� I��u�<Tݏ=����Jd���<��;�zm�<+��V��<Q�<4��@����<�)%=�g��ݣ��H;;�#=$v�;��D�kt:	��;�F�<��L;tW�O�û_��<~�w=3��7���U�V���<�+�;Kh��� �=Z�<W;=�ߺz���Bl����'�!pq=��=CfF��k6�h�^�N�<Zc�D����< �O=J�g�$om��o�<��<b��<��W���{�=�ƶC=3?�Z���+BH;M�*�����7�gI=���!�Ҽd�C�a� =FPл9i=�Ǽ(X=�p�<Q������;K�:�3�;��?�N���ӻ���<�#<��!=��;�W=��g;�K�4�~:ۡ=���<�4A����<,=_%d=;2<�~%<�/!=M&<�^��'2���Y�=��=���f(@={��(e=��T=���;#ZA<�v#=�P�:ǘ���<�u��f6'���4=~�	�,���	X:=�(=.��<1]=
���PM��q<��`�~�6���)<	��<����#�����<�:��^-�<o+<���j����]<fig�L�C��>=ހ�<Y�<���<��=�'N�Ø�<%�=�)���n�&=E<S���<�W�M�R=�����ɼ%��<�L�l�x�-�a=|�*���g;�IS=���<�;y$d�{hʼy{��C߼0�:=��a�5=	�R�jĺN2��dG��K�;�Ѽ�L��]�;V{=OO���c<8[��	�����h=G�L<!ջ��9C�>eS���<���<�6s���Q;4��<y�<�w��⼿J����|�	%���<��5��E�;}p׼\��<��u<o�V=�Ԉ��Q�*�=���=g���=Lv]�� ���9`�t9!��p����¼��3�W>ἇT��[8����}��<Gǐ=�d�����������#<�#C<��޻�z�9�c_��E<��>U=��r���=1R3�Lʷ<�����&���7#���<;�j�Jd��{r=�i���=wֶ<�2<��x<=vY=�_�<�S������ļ�6l����<9}~��p�<�ᘼI=�A	�Q{@<E��6�2=�3��F�<�=�ic<���b�J=�$��u�<<.�Z�xж�h���a;=�쳻)��<��$�<�NV=�.L=�ļ[Q`��i�<sx�A�%�;h-����ڄ��F��Ո<`B�<�4�<�����<1�&=�n;\IC�yNU��O�<j#� <!W;��B���;<�H0�!�q���n=hp%��L�<��<v&W�D=O<�W=R(e���z�	��=� ��Y�<���;'J=�V�lt9;]������:�3(�@L�<#�����7��t���5�\=={����\�����1�<�(�<��=YW��'�3j�<�Լ��<);!=S��#�;=�}7=�3�QbK���<p�6=I�@��z:�t<b���F;�����<晶<Nh;��a��pJ�yk�LH��6��Y��1a<�q7=k/J=�|�<fy�#j.�7�<n�0�����-�Լ.��<T�˼�?�<�U	�g�1��?u�y���c �[�w��Ox���< ��D�<^�^=����K<$��ϼy%<R ��Ny��O��_��w�=��#�\T=�����`^</[�;�j��ц<�w���h=9ٶ�7�)=0�b=ʇY����~�J�{�:򮼜� �U;X=`76���,R�;a��ʍ�<Z/����@懽T,�&"m��m=��A�4�$��q�<B�<�--�Im�<[����<>�n��A�<��/=���ys=��&��(=/CE��r�<Qg�</<f�8�J������t)�;�-j=��z=:m�<��>�D;P7���h��wE��gք<4t�<63=kj�=\8=�3G��S�<]v�� �����=�a1<>�����b=�S<�_h�$7�<���4�=���<o��<j�=�Q
=�����M�C�*<����F���=O�W{�X7=}�W=��8=�iN�$)0��ݱ<�l�w,@��P=� ���n��W=���<���<��=��O�aLȼ����=aa�����;� �:]�<��Ǽ�yQ<]n6=:9=��F<�w�:�\������q����x����
=�^"�@�L��Z＂��<Y���5��C�#Z<b �~��;_[=|�߼�EŻ�8*���_��
w��| �:�<T�?�Z��<�?=�"X����<��i=
�N=���B��}y���:N��Du� �Q����<����
W�}==�툼�Y=�	}=Q�:A>������F
=�7;��;��i�7�=;崼�ѐK�����鄽������<��8��Qp��=S��<���<۵6��E�<�= �<:���=�S;�u1=C5�<�� =wp=x �<q����(Լ�_����-ỹߴ��d�<<��<!)�����U�S�e?=MB���9=m����-��0���=,�L�B�5��<HY�<<�=*�*��QW=xq�=h�<O�
=b�����;6�<濣��l<���|��|�<���)q���Q�<���=D<��a�̜o�{D�2T�N3\=�u(�2�F=IҸ<i��<"�E��+"��z=��<�_�<�U>;9hy<S�==�Vü(�G=>�<>b�<Lz)�������<��H=d5=�/;A�=��<�f����R�����<(=�<��t<q��<��C�0(=�V=p%�<^�b=>T�;.	��˼v	=�b<�x�Umm=��<ձ�=Z���A=6g�<I↻�q�r%�<R-=��+=𾭼���<F�=cJ�<�dԼ��v=H��Ǽ1�	Bn����<.J�p`=�C$=��׼��2=�VV=���E�%�(�2=y��ʛK�e2A=��;D*�̎�<���<̺�<�q�<`�EF<Z9�<��R=�
:��a<�n<i�;zQ�=�M<K4=��7��Ԃ�.B�*k�����_1���f=�n�?5���W	=Rmf=��<�^��6D=_��<S�9���1�z�ἴR<�:e/<�!�X7.���]�������_=4�<�7ϻ���;H"���<���<��e�R��F�<��T�Y�)=�Q4=}ؼ�K =d�=^���Ȍ�,��<�+1=%/�z-%���0�+�>=C٦<4{=��3W-��,�=a8�<6׻<E����<7A�m�1��3��� =�Na<��ՏF����;���<�Ț<v�p�ڭE=)��<��I��. ��i�<���<gcռ>�:ZU��`'<!�T���f��Ƈ���I���?�x4==��=R��Z=�}��I�I���6=z�{��8��)���};��.=�E��>=�j�=}5;�~�<��S�spQ�sL��r�l<.mE��$y<�=�Ͷ=���;Z{�xN����:�"���;=�ΐ< ���u��;�
=��</K=�	����w�M��<�<=rK���]�IK_�:x�<`�==nsT=�:<���<$�<� I�l�:c��_��<�%�<Q��=��r=y
t�Ҟ =ŇJ=M$�<⡼`6?����"b�;���<N �;L4��g|�<�K=���}�5�&=�p%�fe=^@&;�u�<ɪo=�뉽4%��ti=Ý�:�t�<��x<3*=�ES�|�A�Q�׻Ǉ�<��C�	�ȼ�|�<�R=��ż?7�<:Y<�;�<�h#=G઻�z�&�<
�=LR3=�¼/x�<���<�c��7�3�=N`(����<�?G�������<�P3=n�&���V=��Ǽ�� =�8�<Qr�4$����a3=4�&��qF����=D�
���%=�Xh=^�=���<e�<C_�;��R�n�<�#-=67�/�<�'#� Ǆ�9C_=6h=�9�d�<B���m�T�\�0����=rd�<TZ�<I�j<���F[<���{�_4ۼ2��<I���p�ŕ��^� +<t�<��<��<~�$=kve�9u6=J<�hѼ�;�yL=a�v<}�$<�M;�U�ƞ��;��<�YS<�s�;�W�O���R�<%ُ;+�<�\�<�8S<��]�M��<��[:�� <�=,=I��<��B�Y�j��#=>A�����<�կ:�Tq< '��:�ᩔ�r�g<J=�<Y�@�}M�<�<�;5�<%���շ��<\ʼJ�c��⛻]�<e��-�<��G?=����T�;�@=��L��܄�|�&=2��d$b��W�N����%��0_��>�KAK�P� ����<�j�=��������==�h!����<�_
=�v�<��D�I�r:�9=��»$R�H I=	�<"�T��<���<�%=��<�/��0��<�(]���$�v��/p�(HY=E&�<K�����Q��B�<�<�:�fl��\��I�;�d<6=�,ֻP�
=s{�<}�Z=�:��S:<�{=��ռ�$�<V'��}�<nEԼ%n>� ��F���-~�;QII�oO%���I=]L�<=���0�F�<Q�>�o%�6�l=xׯ��8?���m<�씽Z��<�F���-?��ۤ�:^�:F^�<gW=���<bE�[�8����9�!��;��)��4�:��;@�=$����i=D��Gh���=�gR�~�=��T������Ҽzi�<�����t: o=fH=)UX=Ǚ �����<f�"=�虽b�K<��ټW�p� L-<�S�>h�<�2=h��<cS+=��c���#���t=o(��P=OS�;��<#?�jL����O=��{�JE�J��<�=�<}��J�ݼ�
�Vؿ</���T�,�P�j52=�H�<L/Ѽ~<��M��$���{�<�������{=1�"<�y =N�<��=g=��;��Z��Ċ=�,ż���V`�;E�8=�`�=齤� P.�ì�<�����C���)=Bɹ<a������<CC=�(=L���� ��e=}�s�����gN��ټ�4����A�)O����#�f�<����ٟ<�mP<��<��I=^Ƽ�{�<ր��7�:��T��ʕ<��<$�X�Q<�Q��5��J�@�}ü�:��r��O�=N��<�#�<�vлu!λ*g^=�5=Z�.=�%�<�sA�ܖ4<ŋ����<5�#:��=��Z���=��T;��=�Z���6����=<L.���d���;�N9��!I=�m�v�8=u�P<�Z{=�	�;

�K%v�{O�<JB=^���Ws=�c���]ݻ�u=�w<�Z<�^��T<��@=���<FE��W�<�=C�vX=>��� =�輘���V=<��>8���>���]����<�?k�Z����hv=� �<�c�<m�=�\:=ru��(�1�8cK�0i�<G/꼜�'�G��>�M=2<$���5<����sDh=��7�9y�<6��<�b��B�R�{z�<��C=�<&����<x��<kw�;Z'׻�Ϙ��_=r*�ӱL�s��<琽2�<�^1=<�ۺ�\�����<<tS�S5�<����r=}���y'=�f}��
�;�F<&��<���<�)=2�1�E
@����͛�]���%�!P�K 3��s=��%�z�Y=�H�<��<�!������{�q���\=N��"�0=�w��x�<��;��֧�?5j��}L���b*����<��<��J;���9<Q�����{��`���A-<����W���\��u�=�|�:>���AL����Gǵ���;;w�<��=�e�S�]���<��6�!Q��L]!�M��< =�{*����<��=	����z��	=��N��g4�D����=��B���A;�;=� l�%��@rg���*<���<����)?��B��|��;M��^�=�M =>~��_഼
�V�Q�ɹأ��_��<G�e���@=���wi=�x^=�Do=Y��<��5=��9�v!�I�<$��<77=�"=p�V�ݳ�;uC/�f���"0_<�Sܼ���<e�C<���4�<ym�=������8�<��漣��nP3�w;#����Mx�<�/��B���A�~u>=ܖڼz_�T��}�%=�='�\<d�<���<�R���e=��1���}���:���=zK=?� =(Z޼�<��b�,��<7~��?�,%=jA=�=P^=�����0=�P���;<ow"=j|���=��#��==�Ҽٝh��I;������^S=��=V<�����;X�<ԕ<��k=�<lt�;)�6��ɼ-�<�)�=*�
�k e=�1��噞�@��6�'���	�Dc�<��<5��<$iZ=A�!�j�P�g�:<�Q=��/�&K<ޝ<m����Ƽ �4<��6��{=d(ټ���W������<vW�<���T=�W#= �2�D�V=��׼�:<�o�=�|o�=�=B\%<C��<k�仩G���b=u	8�@�����7��<=T�
�-�!�X f��&�<�@=����3�t7�<�k��	�	�9�x�E=+��:{�d��s;�iܻm��<��]=��-<QE
=��G=����;<� ]j=�c�<S	��n����<_��;�R�<���<	ʬ��̃�-�һ�mh���k=)�#<N��<�Y���<e�<2+=�<Y�ü���q�<6Vn<tWF=��<P =-�=�=G=��2��SD=��ɼwK��l��/D=H�]=)�N���B=��j=To_�.dl<��%�9s�;I��::�<�.�<y�
=p>��P�<���<���<6��<":�9�.��yW��rj��PB=�1|<5��|P=8p����<RV=Yv_��d>�x4=��P�L=�O�<�]<����2A�`�Ӽ��M���μ�z�~N�<`R<'U:<+� =+K%=�_�<`{=��l=,��{��<�t��w�;�F}�y�C�M�����< (z��	=��R�#b���NM���?�M�4��S9�1S;�,D=�ہ='��<#
=����������g=G;M=x�<-|�F����d;��0�SW+��nO����<�d=j�<�����e�H=LoR=���o=��t={�'���������wd#=$��Z��,�<@�b=x�Z=w���Ռ=^��<de<w�_��p7<Ը=$��<�0��.ɼ,0�;�*=uA<b��Y�;36����<*
h;q�X=����19=ekX=A\;�_��;+\��ͬX��=�[=�H��e>�<7c$�]�м�v»�h)���o�1�L=��Ӽd���̼�E��Ԓ<<�ɗ �Cg�<.z�<O��0v.�\n=J�鼓��J:���-��!O<��q��X�<|=p�z;��=�j\����[S%���/=�˼�g2������A���<�La��*@��Xp��s������,��.X=j�,�*_�;[��=�h=C-9�VC6=)H0=�s�������R�:=�S�<Y7=\k�/���o�K�<����H��!�����b�$=���<�54=_gV<�������eΏ<���<�"=U"2<���=��=�>b=�do=�*��`I<�׼W��;�t���]� ?"��lǼ�����P��3[�)]�<Y��ne=�l{<C�W��?�<�	O���=��8<�0�v��9��#<���Z:��0=�ay���U��J��-��9j��d:�7��6��<*ծ<������v<W�Ѽ�
=w��<[h=���<���s��<�O �� ���D���8=ܧ�<Kl�;U��FMt�	�ɼ��==+=�=��(�
T�<O`q;���<�*=�+�pyX=�f�<,p�<���:�ٯ;���C<r�@=E(ȼgL��b�<�ܼA�,���q��^5��I�M�<=���<8Q����<�e�<��N��[�����S�<�2�ц��.Ѩ�'�?=[6�f�|�t��R[�<��=�=��H`<fvk��i
:´�<H%@=�8=��c�Jh�:|g��y"=a�;��ڼm˼2E=*=�I_<��)�v��<��D��;�!t������=�@��;b18>��<1d˼t�`��ӼHͺ+AJ�"������-=��;:�q����<�O5�&#=��3����1�;��<`���Ko;�O{�/�9��X<h��lP�<1u�����q=����r�L@0=j���S �;�M����;�9x�)>+�T�<�8�<T0V=b =��ҼV��<��}�Ĝ軳A��2�;MJy�P ����<�5��œ<���<��:=�0���%����<�6�;puq=/S�q�b�YE��C�J:���<z=�<�@���<F�=��=��Z=����$-�;�#X�V`5��;���=O�L�R?=�<=DN�<�t���CV���)�����Ϟ�N��5k=y�<]���e�|���J�;��
�J�B=�|�<�6��3=�J=J�b;&�<�l�;�����Ἅ���ҳ��V�9�w�:���9�%�=�&/=��j<���B�<���d�=xJV���Լ���;r8	�Zxs<�
`�j�%�L�=���<��Q��&:�!b=i���Q'=<�G���7<A��m=v�a=��=��<�K�<�¼�.a�}.��@�і�|�E=nn=���<>!<�������<���<	�����ȯi��p�����������c�6�C�����>?<B�<4y=�1W<��4���<�jἝ�d=�d=��<�	���Y=;�v���A=TEO�&F*�eӼ�q0=���;mw <��,���<����=*V=�)K=����}.=���<G p��̇�����߮M<�pj����#W�=j�\��2�X�^�^<+4F=�!�<� �<�6��)'f��M���_o=z=���!\=Ϻ����<�{=�֟�L2�3W�;��W=L\=W����:=�YǼ�p= !M�1:x���T=���<!&��$�;�^y<1�߻hB
=q-=��1=�} �M/��M�<9�Q�XV1��/=<�(1�6Qi��Q<�k8=��f<��;.D"=�<��*���*�: �<�y�:���v��<��B=bk=xS����@=YBu�]�<����;7��z��M�z�U<��(�c=�3�<(/:=1�A��?o<�SG���$��涼�$N=�!=�Q�K^�}L���Y��덼�����QV=��E<�C��(4=;�=yp��4&�Y��<ah0��
��!�<ܥ=*�<��#<�9=��D������&��mN�͒P����<��.�zUS��lD�3'�<~%=�b���L#=U�:vq=�'�q�Z\��*�=��.�$�W=E�����r=xC�<&i(�ԉ�;\9(=�߭�pvQ:�<��R��4~�7�<%�Q��&���<�0=�	/�t��Oռ���<��D=�%=*��<��C<�8y=����N=ǳ�<;4�;��<����`=��9��2���G�>u==*\=|�=�~�<�f0������*<P�	���B��!w<��=#��<��=�=�C>�Ds�<!V
=w-a<T��eb=�����~;�&�<��T<�F=�ú>�8=�I?=����i;�N��s�;��4��\� PW<� �<��=�'!=+Rz�9�s�b\$��K4�%G���<�����!�E���<BB^� �~<���<\�<m��=u㼬�t�R;<'�)=�~H=,�T=��<j�@�ec��1=$�"�g��<��ݻ��i<�@K<�eٻ�M=z(�<H�<��w�B��;��=����Y��%=��� �*=,#a�҄�;�
%=��<�e��}�<b2F=XJ<;.�b�� =���Kk=X�R�ѐ���<<���<t����F���j=���<m�����5�H=p����=XSq����>�=�>�<7-��\���U?=�c<���`�-5V�8#ݼ�6��=l�2=3=�<s됻�8����9<��t=����c=b�X�<j�B��\�=��=�|<��K=O���=X\-�$7�kj=�P2��l�6V�zM���I�����<T���=�<���zh�<GV)���<�s5=�� ��sa=X�Q=����[<�g���I1=��C<��O���p=�j�/<��d�;���=��<��%�7��<�����᫼1'5=-_�WD:=&<�ļ�j=��P=�4=�2�;����nz���zj�<�^�<�#�+c����=��Z���<�GJ9Nv��#����)����<�qx<s�<#佼�/����_!�2 ���h�J�S��4F=�jy<��o���W�9W�d�= ��"tB=�&'<GtV:wN������:=T	z���Q�=�B:=;�P;8O=t>%=�I�<��B<d=J�=0�����;��<,���=Y	=�%��Ⱥ��؟+=��g��E<ZS�6W�<��P�����eu=5w�<z�<I(t�s"��.����*2���<!66=�������?ua��\�;��;�j�>m�To.=:
<vJ�;��R�NVټJ�"���<��4��W���c��\�<n�9=Щ3�ܒ˻3$=]����;�<,5��[�=��9�C� =(�_;����O=�;�9��\=׹�Q�׻7Լ'���H�:�쮼>Ȳ�����GRw���r<"�5<Ś�DLq�
�k�g0g<�C=�[���ט<~�<��s�>�8��e���hP��B�^ǟ�s�;���<��
�R�$=��n=��黰
2=��l��	=ʉ^�}�@�H5뼸��<�ۏ:�*{=|�\�v���:�;=_)��<�~	�ҕ�<p t=6vo=�9�->`<�w;d6��5����cRn<����Y׼S<�<�F<��ͺ�Rj=�Qv��(9=��6=�G@=�$ =	C�;�*<�%V=�Pػ���ޝ@�C�$�p��<�[*= �I=(ٝ<�o<�F.�.�<~���CU�iu*���4=�1d<R�̈�s���eѹ�z=ؒo�K��<阮=�^3=�Ii�^+��eld=ì�<ݿ����e<��<�;U<�y=W-=�y+=��y�����C>���=��<�^F����
n?=<51=�p=�qb���:*0H���Ӽ@H��5߬�U�&��.��I�$�	�m:=�K<�"���t!=:T�<��=<���;^�e��+<<�P=��.<�.�<���9��L��==+=�F�>tȼ}-���>��qQ�-TT<�hS<z�<�g;D(!���H�΂=4��<��;�:�<S�#��"ۻ2���*=Z���(�q<�i=h��H<%����>c��)V=����z��bP=)�=A0=߿
=���f=;=-\����:��e=�@={׸<!J<;�>_;!aμ[*����:p��<Ul�s�b=#v���<�((�5=��O<��w=�[�=�,���2�o���Y=`��;C��;9�:�`�k<Y��=M���ϼ�� =(g.���Q�%�Q<��l<b_���0�|Е������%=6�G��}�<��#=p�;&�=�M��1�^��{�;锹��~����O=��@=�ZͻN֦���Ż&8�m�<�1��=��_�����^^�#t�<\�V=��م=��A��:��[BV=\T;=����D�<I*�<®=
��<O6�;��F=�+<��g�i��<T4E=�2L��x�;ʫk�2?<_(�54 ��Q=C�=-\J=����!v�Zi-=�����4���U=�/�<C�����<c�s=�m�=|4�"@�<���;gr:�{v���2�>���E=@��̛1=iVE�3� <�5��4�;�a$��>#=�mb=L�?��pu:4�<m��<��R�b�>�o�:�Mڊ<�K=�Z�;Z��=[���=8=9�=<�#<������)=�f�EY����;��ȼ��<$�B<`[<Z"���պO�J���=�Cd=҈S=�i��bq��� =M}P����V0�:�ֿ<�i�x-=�`�<��>���/=o��<�w�<�F==���%=��	��7=쮜��J=�����X��=JKX�s0���V�=�V=�'&<F�h=/]�1�=����Ь:A�Q=�HX=0D='��<�>^=��n<��e����%���g�=e�;nBb��;k�)�ě�<|<��ޑǼ��_<Y���x��<�5м��Z�`��]��<5W0���N�7 �=�=�=���X=��=�ࢼb��:�R%=R�=��<�[R�׫:=k	�=���<�4+� ~|=�-��A8���G=&*<z��QZ�/˻�=�"���A=�ؼi�=MV={� ��{2�۳@�:5�;J�<���<gfP=��ʼz�F�<3*0<��<_������L�)]�<K����k=�b�<A��;�X6�*g <]g=X�߻TB�=m�ڼ��-<�:=��;��f�*wn=5�һ�o �Td<ip�=�/=u��<o]Ϻ��3=�t���x��O/=�w&=�e�<�f$=��<�0���,�<i����g<H�D=c�{���j�)<8<h�⼐��;��Y�Z�&=My�'�b�f<�=���<	��<�u�V�K<�"=��<�G/=en=x��<��e�֯L�M�3=UJ�;��B=��_��=*�i�����tջM�J��<�63=�%!:፻b�v=ҿ=pLg���<�bz<�żĽ"��(=�r;s��u)E��I� 1�<�%���\�[5=�����;�<=����b�<ծU<��\<�fW��qɼ�p_��_�sZH�Xf�<�P�X�>=�8�9�];�e�<�!�<�%���=tf���e���=?�1=C!b��%�p<�(�<���jX=��O�@8w�Dj�dJ�<3�����7<,��@����&�;W`� Z=��˼�s+����<�w�ZLN��ԍ�~�����6<�}�'�����d=��)�󛃼�=.s�AgǻwӼ�"F=]ʼ�0��ቼ#�6<��j��7s;IK;���=�Q�Q|�;�2�<~"Ҽ��O<],��W���g?��?=�o�<m�:R�U��>|�AR}7#�_=ڃ�<]J={g�;;٬��W�qs�+in<9��<l�h=_� =����ȇ=�'=Eˢ����<���<H-\���>=��
;-9=A��;�E��I=�����<Ev���T=�3�Ek��ׯS=��'����j� ��zs�_�%��Hq<A�	==a� �����:ڔ���Ӻq ��f¼2 8=RI�<Ԍ��p���A�L=����z<Q�<��I5�p������b��;f��<�J=��<-<������I�oz\=�p=0�&���;d?=�$/=��'=���M=l�$��<u����rf<�u=�#=��</S	=�f�iR�����O���W��[��$l��2O��|�c��m�0풻�(�v�=I�缶�U=�K�:QSy=3,�<2l:��7=[=g�<#��<߻��˼mX=d��b�C��-?��;:�����`㼝7�(61����;�Pn<I�:ՄI=�+=W'�Ä�<��><�����Q�Apr=N¼21��&�<W��<lhr<���$KƼ�Ls=݇&=(�O=��F=��� $м�>=�Rc��9!�D�ú�2�<��D=�,=�:�dYU�r�H���Y=
$Ҽ�/����:��6����F��y�R�Y1q��z�<[¤9X�<t�=r�<Kk�=[S-=���<ܑ=.�Q=찒;�)���;7�<�7;6����;1�G�?�I���P�5��*�����\=lp�@�����,����.����J=*J<'���bP=˽=�I�<"�7=Y��͔:=�쯻�d�5��:�}j;�~M=Fe�<A��������e�;� 
=�8=��ϼn��<��p=�D#��!=��5�J���a;�U�[���U��!=�V���j;����]Y_��V���k�ku���p�;��*���Y=gq�<���<P�3��>�<�f�<g�<��@��,A=ww�<��a�M��;��=h��<���:<��<�{�<�1�<X2Z<��Ǉ��를�{=I�=�=�5@<���;S]��Z�	=�t�<%=�� �-���s�=�pt�I�t�(������_:�S:]<��$���1�z<P]�/Q	=��W=X��;Al#=��=7�;=s��Ƌ�<mu[=K�E�T�&=�%@�����8�A����*��������f�ϻ�:��nF=����p:���<2�G�鄍�2��;%-�H��<J{q='UV=yſ<9��:�n=WjM=��弙Od=kz�3��<�:L������̢�-��ͦu�Ǥ�<�Q=Wߺr(�@8T=�E=��*=�>k<4�;Y�<��漢�k;j�I=DWz=#rR:�_�;.%�<"�t=���ju3=��#��p�;��<T��=�7R<���շ��9:¼PsO�o�g��ED=�8�� ��[���E<�Z7�a^a����#1�9�P=�/=�0���=$;���h=y��;�W�<C�S=_�<���<s*$��d�<��l�@=ٚ	�="�<�޴�T{G<$�Ի4F�<ݮ�W=)��oa=Ċ�pW�<,���oZ=�,���qһ�,=JS=�+���%��9��lI7����'�=<�Ȗ�Y��<z:s<� <㞉�oH7=��I=SP=�+�0�¼T���(�X�y/�;c*�<�d�h�d<<�:�.Y�<6\=��H��.<��I=��<��<"��<�1��ڷ<�C<=7�:=��<�<�<�ً��C��`χ��tX��f�Y.,�!�&;�J,=9�;�6L= �`=8~S�gE)��{V�y=�
$=�<j3�v�:=^\c�us�Aq�;��A;!�$�t<[������<��g=P%6��!���z�uՁ��8�<�!z=�G�<ث]=������ͼ�1��p���K�F<��b��r
=0o=��<�L�\���x�<�.P=�?� ���9�3
��rR< �����6<�|`�4Ua�Lz$�*�=����V =��7=Z��<uRt=�����-<CA��x^����<�MP�k3G��H�<�4=�A��m&�e=;+�;w;k����څ<�{�T�=K�\�O�;�E|<�P�<5I\�&�^���3=K�=��C��Y�T,<�m$=�r=[�����==f��EO|=���<b��;bTӻ*��<G.�u�<k! �[1�;c�<�k��6g��	�<��(=�߄�&���Q �9~L=����BG������;�Bt��"/=|��:��=	�9�� <�����#*��pp��	�� s=��g�S�U�V�4=AB������<\�����<��!��>=��T��3E=+�<�	8�A�\=�ػ8+<�-�]�<�Qݹ�');�ʾ��9=�@�<� ��{ּ��<=v*4�&�W=����u>��-A<�CP�1e�k���仼x��W��a��;mt ��x=���fD�<k�=�q���m&=r)v=.M~�q|�<֣P����<H
&="h��嗼"����	��v*�Ǌ�<��=�W���}8��q�[�%:������0=D��<�-�<��=0�$<]�;�#Lu��E���H<��<p4g:�7c����<�H&=�]T�P_��9<�ё���/<J!��[-=0d=�=����<n!=j��<M7������W;��T����;g]<dR_=y��<��f��-%=s�1�A4s���{��3g=����f�0M�nD=]=�;�=k=�"�l�������쳻��9<Sf!=��˻��;�t)�6��eV�C�J��B�<���UG";N�b���*<�6?<�ּJ&�[T�<�Q=���<�B������}���#X�c��"g�j&=&L):σ$=j��;�=%A=<K�9����<?�4=,<n^���-=� .=��<��$=�Z1�uH�<bs�<��=�;=�%���=|y$=
8��z;ۊ�<��E��QN<�zټ��d<D��ϗT=D6&=��<�^<d��m+=R�<�� =��A��9�)�=�"�=q<�5���.�|,(��3�<�DO=�gJ�w�� �_=��[��y=ϦǼ��OH=\�P<�_;�O<~i��#b�<�8<-tA�(&���<ĶR�����,'���d=a�߼�	�<���� �e��䃼�.E��9x<��<��2�	��<�A�qn�<٨�����<^��<�%�����<��<&��<)佼��r<Z��<�f*��(C=��;Y�$=��=�߼:��;���ݙ#=t˜�;Z'=��Ի�� ���5_=��K�V<�\<�z{L��?ϼ��F��%2=`)g;�=���<�*<����</M�;�+ع������o��P��<OuO�d+�<�;I�d�2�'��輜,\�G��ߋ��t �����k�;��j@����P�؍�[����z�l9�<�@�<�Z���+�������<\��"[G9
l��!�:Q�l;�(:dK=����,�<q�D�#���utۼ�;==X�D=��=bO^8��'=�)J=l%K=���yƼ��㻍j�;�"=p"��%��<��Lt�Q9v�����q>��f:�(�(�P��<�=A?a�``<�M�<�0<=�������WA=��);���<�t.�7��<L�R��G���+�N&����s<(�f���=V%�<%�Ȼ
,=|�
=�<.?�=A{x��1};�lQ�ڍ�<��传ȝ�=D=��@�f'�;�#='�ϼ�G�i~��>C=M{�v���<V�*�9<��E4&<Cm|=F�J=}u��&��E�<`�t
'��j���=+ؘ<R��<�ۖ�w��<k����f��8V��։<�DV=*�<�/�� ռ�J��=�5G=R�F�P�UȮ<$En���j; ���3�C��l���<��E����:s�?=Co�)E޼~Q=�h�<�ç<u};�1 ���=��8<���u��;r�ܼ���<��N=���J+=�r<9sȺ��#=WU4<���;}�H�l��<��`=���;<�=`c3<#�����u��f\����<�7��C�)�Y�S=v}_=k�缀�\=h�]=�tl��h&�Rl4=�� =�tS=�>-=xL��Ъ[�TL\��T=ݶ#�BX
��3�:�p�+�\x�;3	_=�=w��<;W:���%=�BD�^=�������G��;F�z�kƆ��Cz���6<X�Z���<w�(<�]\���=�ܼ����_��Ǹ��x�;&�<Ar@=��<|��<J��	�<�P`=��<���=�%�]�a�/�>���o���Q;I���<mޯ���1=�����=�*=��<�"=��;-(D��
�:��V�XZ���V�	_���t9<f�v;(6�<q)�����<��=��+��a=��m��!׼�*�����Ճ&��(=}.��)&��$��tR=΋���׻`�a={��9� H;�i�<o��mrԻq�;g��;�{�Ɇ��ռJ�#<��E=�`�����Ԁ¼wI;����9=H:�pg�|��Q�n<�S;t�<�滼�V ��n�<��N=���:�{��Zn<\<ݼ�t3�uü�^%��L�*�N���=�瘻��Ӽɹe�O��<;�v���5��s�r�X=;3=���<��;�� =���M=��3=BR=>H<�wo=��=!#-=���=dt����@�6=���$�Z=�ur<����v(���G�p ���8=�c;�xN=5x/�X����<
�U=��=��D=tOI=���Y��[�<g�=�m��(�<��j=|��<�[!;\�<���=�/�<�ʈ<�rH���I�(/�<�#=0@=q��;�<}�q���z�"kV�^Q �w=L�&=-|�<��ۼ
��<2�E�m����4<}�μ�d=��%=�̇;T����X��zm�d9@=l�M<7�[�'���w�;��0���G=B�3��9i=!�D���l��ȶ����K����ּEQr�;r�<��=z�j��r��9��j3���3=-G=+]C�Ԝ�|�=��%��v=Q��<����p���޺3��[�:�<䨡��AO�1��;�$���R��Ǽ�{=#�}=��<h�0=%�U=�9]�`FH��4=$�<�D';t�1<��.<⚼ø;=�\�;�
����%=��a: [:�/=�e0=�WT��k���';^�<u�`=�q�����<6F��{�%��X<l��<޼EU����:L]B=<�< MP=��U���<q��=V^==+0i<�d ;�,Ż�M<
VҼ�3ٻ�D��HN=�c==��8=�K�����D0q���º���<���<����$�==��L=�r�=䡼}��<E�K�bC��� �}��:;�<�f(=��;�ۼ($$=�2�<��<!�ػ�� �3X�;y��<��¼P3ػ��<KX8<0!�Mm=��1�&�$��%i<�$K�"��<����Lz�6��<�-y<�xW=��<�U�I��W἗�Z��b?�+5鼗�<��<�kI���x���M�WbL��i�7f =f����ʼ�f'=8�;.���ʎ����:".4�2�	=�={��.�{���IE����n���p=j6=�\�R�<��<)������;�m�<ک��χ��{o=/�e<Yغ���8���S<(C=�u��`=D�M�-ғ<n�*�V,�=��=�a=�	F�5�;=�B�Ʒ�2�$=�л�J�'���24=�F���c@�_;=iI��[���1�C��;�=a��<����]�)�b"=�V�l����v��:=��;<<_|<M@=�>=�;���u���+=]1=�6�'ꂼeлl̾<���[��g�ּ�nD=�2I<Nq=��0=b�G��?e=��o<-�N=�MD�;�FK��)(�����2��=	�p:�b=��(<�}ἂ;C==���n"=3S.<�d�=eٟ����c�<ƙ��=)=ޯ��=D�<�#��;l㒻�a�����w=�}%�T�S�j�=[Zi<M�<jS�<Y}�<��j=�\�<3�;��?�(H��{��2<��-=��������1�)
=g��<�Yo��譼?9<�m>=�������;���<�q�<XL`�DYc<�+����f0���<�5�<4cI��|�(��d�(�UR�= G+<�C=���t�<��V<�̿���ۼ�P<()���y��h1=s=<�$��<?�c<k���0<�f9=���0S�<e�;<Q�<a:E��<2ՠ��^�<e���;��<B)=<��N�-�R=$�=�ؼ��T=��==zO<W,�<a;�tu!=�rm�V�<jU:q'�r���V;�54=��v<eh�<�r˼��T���<��伍����~�=Nܻ<*̽;"x\=J&r�	<:;JGϼY��<H=��=s�;�q:=�!4=�+�<5�)=�&�=�F��E$.�����#��ڻ�=?�q=�fO=?���Ed���|��20=�@9�EA=���<�J�� �<^�h=(t�<U�<ß<��޼�&:SrY�J_���G�<����E<a�=�O2;���<�s,��%�H<��<Hg<pj<v"=R��Q�;٬��:&�q����N=lʻ�V =,�<B�ӻ��'��y�<�i��¡ػY��<�=������Z+�����au<��<�\=ZQ����4<Tr�_�e������13�ݓ=��8=@. <�c���<�x.<�����;Ge<Dl=��<O)��bs=�&=<�>S=?�e=w ��ݬ�<ek��P�����}.y����9.d%=��&=b�a<K=C	���"":ŝ<�=s�=������<K'�	Ŕ:�W���={i=v��<��<w�4=I���{
�s��<l�\�/<̩��p#L��S+�N�;��='��ѡ<��㼪�U��=	뺼��=x^<p�B�l ��(=���<sq:7݇<z� ���#=Y�m�3�<�ay=�6�?M��n=�\$�,���b=������!�M<k$ּv���,A�U˝<ݦ-=�uм^�<��C���A���~:D�]<ۥ=�ֺ<�bL=i:l= Y1=K ��%�w��[q����<�ß<H�0=�iE�G�=Q L=M��<��*==#k�1�<'mK<��������<�Pe=<`�=�[�b�i�-�D�����8A=N�j<Y���=�ZX��y;�V(=1%i=��p=�2=��a<5��<�y =ׅ�<ȭT�u崼�\=I2<Lz��HZ�q��<[��<��=g���R<��J�S{��vݻ0����W<1t��&z���|���i=��K�A�
=p+껕f�=��ۻ�k=�Yܼc�=[Q�<ٳ@=��0�'�9��H�;��V<*�b;�
���=�Sd��b���u=P����;�BQ���K�|�&�mN<N �uX=��=3|��H��=����:C�Ӽ&X<��WV���Y� E=$�޼�~6�&�f�b��a���ƻ��u��}=�Sμ�=͑=:v-�v:�<7�ռY�<�.���ۻ�.���*���S���d;�����G=y'ռ(=�y�<w�.=	�,�Ǘ�<䂽<�C==}����BLT=�� =ǟ>�ˌ =y�;=jΊ=;=�$���+�<N!L�<��Ӽ)=��/<f_ʼ8e<�X�~�;��.8Ynm�����@�9�@L�+�a�d}P=����<9:���	<��<�G�;*���W=��'<��X;���q��4J=܈O<mR=Ρ��W�ޙ)=~w�z?=tx����'����<C�@���,t����}�9=י�<
�<'�4��Q=orp��p��qLc;��.��T��}=�?Ƽ�Ѽ�y�<�F�$��<��;�⯻�k=�׊�� �<���<�<E/+�$��n��9��<`��<�
Z=���cA����ͼ=m� �K=�C�I)�<�#�$=U�k�0Z�<#��d���?NB���<B�=�嬼╊<x�ϼ]�=�F <�X<�<~� �F��<W�!�ORG���K��2;
�
�N`����<��=�pt=j���k@<�<wR�;CV����<��;. =��=�@� ��=5o-�I�<D����=<&�f
��|=\�ʼ��,��+�v�8>B�UNI�u�/��ݺ� O��JмLK=�X��[dZ���=�Gx<��9���5��h�<��.��������ߺe�<��<�sS���)���Sj<�2Ҽ�����;=�d4<�d���B�^w�=�
����;�Y��`=P=��
<޷��"=3�<�t�<ŊJ�Z<Q4�Hj���)��$�;�-~�U+�<˄e����:A�=~��<��ٻ����x�=]=� ;�"�:6��̪���X��B��k�(���dkF;�>��	����f�����9��=d��Ȱ�<�ݺ���<q�=O�9�׺V�'�#=^g�eh�a�>��@�<E�E�#X=N�8=�X-<h�=�p<<���
8˼%h�up �t����y�<��(�?�p�ݮ�yJ6<�,<�N!f=z
�{^Ѽ��K=U��<C�e�ز<i1= �*��*�;��a=�d=q�=��by�<��
=g9=��_��M���������E%=��=��k���e���A<��Q�	]=q�N<�!)=3z�<�C=���<Ǵ��]�<=
�w=k.=�W9=���gi1;?Iq=�>a�U�4=����4��q�G!u=:�;�b=%�=�57<���h#<���y�?��<�<�<6�F�=��
�`�$�<#�<�U<���Z=5�{�z��<��� �뼍O�<r�һ<��<��Y=�GT��4*�S�j��_�<�"��k�9�_�K�=���;��n=8���&$�<o�<��<0=��.<�	#��OA=(�¼U�ϼt ��ԁu=n\��;D�,J����<��<�|��8=n��5<Y	��<Lw�:�f�����}�g=�ht<�8�<G~<��̏<��s��m����5=�r�J�= _���\u�^�<mXz<��%��� =Qż<�jd=D{`��r�<:]@���q���C�^T ��/[���<��b==�r��mI=�������鹋���:=��=�@=S%�=G��=�8�=�����H=�⾻�غ�W=ROh�<<��? ����<�9E������w����<��H��<�.=^��g�Cޜ;��{�}�G�8f�<uwһ��<��^�OI<G�5=N�����݊�<T+=C=N�=$�ؼ@�<� �{�<6��;l�=:q��1�=5<�;�`,��`��'���d�R��=P50��z� �=ÎT=��e����!�:�y<S���Ҋ=���<����CW�/�L=u�����<�=<�'������,P=׷���h�<ɠ�<c�;���<�I$���s<�z#�s��<������_����p:b���xu��J��<�ż���\��V.@=�U�<�Y��a�D��>�;�r�<�6W<��&=m�"=���<)�={�>=�J<J�u�s*��$�;�t�ɨ>;ت�<��μ�'���=a�.�\
=�.$?=l܃�]�<A\=H��V�<���;ocX�ۿ������d=+N�<=� =��ϼQa<�&�7�%���Ip=����J¼��>=�d�����;V���he�q®�� ����
=�o���p:t ���=ʻ��W�<	O5�"3L��$=���<�R���=�Ů��1v�|\�a<�<���9$�4E�<�J�[ʳ��X�<p�I=���(�t5�@�4��}���h����� �0�.�_��tX�1�ؼv`=��A�J�K�d��<�lH='i�< #^=(p���	����<MU@�>�\���(<�C�r"�CC��+HJ9��ݻ�r=C�>= j�����<hS=$T:pF�=:7n��C��;�E?<;�ټ�=�<�<�;�^=��ܼ�OżE=G�]���H<7( =�_��Pd<z��<�
;6�=tcS���b<��Լ��;�,j���㆚�NW=�38�ݑ=-y<7���G�Z��X�˼[E=�h:���&%="e��~Լ��<?c�4ȳ;²%=�+ºL�o=�:=Fn�<��j�\�X�w�<^=��A=4�<���"]��S��S�;����,���V=$�"��sK�6�༡�,<>�m����<F������F'=��;��>=��|=�>��)��<⡈=b.������o޼�	/�`zi���N<6�:���=��<�X����<���c=MT��� =<�<�l�����;��<ˎ< +��V�8eW�����<J�<0��<\�;[2q=�5���X���H9��c��=��<��+���;��r���B���;`т��`=%+��)�<��W�BŤ�R���Y,=�/<�TwK���<Q}Ǽ=�=���<�B�;��<�~�rS�Ĝ�<nP8=H��:�����/μ��=�%1�J��<���<=:9<@>�'l̺8tB=�`<�_�kZ�0�<��-�ZR=��;'T=�CA���q<���;M���dD===n�.<���<SF;���<�D<3ݝ;>�<����+�R��ױ�
n��od�aC�M�����,����� �;�=(�C���W�N6?;���7<@���V<��<4�:��;](<�=K�=h�G�\�"��z�<`F��=E4O�p@=_x����9��=æ�#;=��<��.�ۮ�<�Vg��(=�5�</��<�oE�M�T�[�V=X����)=��G=�V>=��<k=`�9��N];��$=�<`퉼!��<�
��G�<�|O=K��<F0=�}:�[�@=�H�7��`�<Q S=��m=�=��&�:��<�P�w�����;%�����<���SS�<���<�y7�(�`==� �^��s뼖�:��<N��<���'�E=�$=��ټ�NQ;�<��#��M{��D�;�-���*�<��¼�H�'�D���8<��ػ;s�<�ҿ�kZ=9���;�G=��c=fY4�s_=�N.=�D=�yQ=,�=�2��A�T��|��<��F������<�?˼�+������=�6;��z=L�_=�-̻ )^=B���9���;=��u�������0��-��g
<sC��+y*=�e�;Ȋ�<�K�<%ܲ<8+j=��<8d�v���uHW=*H=
z3�t���;-����_�'�n<ET���R=�<�x7=��������F���@�.=����Dڶ�Eu9�w%=��(E<�)l<3��<�e<��?=�ü���<P��<k'x�g�0<��ػ�y��K�<ɺ��K-<
CJ=�P<@Y�Uڻ�&=�3=��;ŕܼ�`f��em=\ ��M��ȼ��q�V�+=�Ĩ<�p>��P:��XV�*7���Y����o?=={��3�<� S�6ʟ:
/=�,+���<i��;��<S��b&�|�<��e=T�\=e�K=ϐC����:c
h����<B�n="��xOƼ|�(=]�<�E<�8�<Ǹ`=�f��O*=��!���I=�ʒ�CR��aC�r�=����t2򼃙9��{u<�c�<�(�<�r��> �E=���G?G=Q�<[J�;��S=�:G=;�<����Z�\5=ʔ,=R��� N���;�T�g�v�c=A]g�	1��Oף�[�ٻ� H<�[����<�;�c���� ��X=_E���.=N;= b.�Q=��(=R쌽qn����5zj=17T��V`��%"=i\���6::�7��qg=w��; tD��zS����)�<:xO���2���7�b�_<�[��؈��G��ď`<H�;V��<����R^９=����<=G���M��I�� ��<��<�ω��Y/=��<��;=�=�S*��D ��x=t��;���O��@��q����^�Lܩ�qJ&<��=.��<��ǻ�u:��[m=�1���Տ�%c=��V�MUݼ[eB��k�����(�ݢ=7�<٘�<�����(=�»ҳU��#��;��<"G�<��n=������ż�O���#�3�<��Լ���<vw =C���~c�O�S�$[g�2�<�5<n��:��T<��r=p`��$=v
='���!�<`��<�};G����#<V=Q��<Q������h+ ���2=�������<>�Q��a|<=�<�@=�v�6��<4X6�.�����=]_2��R,=/�{:`1=%0�(X���1=��Z��@&��j4����<�i>=�n2=��"=ëR=��&<^��K�<��:�07�<h�6=�_=��,=�޼L�b<j�=/����<� �	H�/2h<����=O�2�.��r|�<�c< ����_�<YX�<�G=�gZ=�%h=��S��续Py=�r��!!�<v}�;�޺j};aw�;��{<��ջ�ws=��Z��J�;�\�ѹ��.��]q�:�lF=򉷼�sw;U�=u>�h�'�,=�s<��=w�<c��;��<�zH��4�<͗���=k E�n s��e*<��=*��<oot���?=K��S�=r$;���<�
<*��<��^��ի;5D�N�5=G/l��_��{��*Y!�f��;pZ�7@�F�=�/;�����#�F�[=4�'���2�{=�D!��3�H�*�#������E��E� !=�KW��H�<�)��2r=���;AzԻp55�m�j�ڥ���-=萭���%=��|<��޼;���_��?�R���<��1<��"��
=h$��5V�=��=�f=�C׹[�:�(��~:c=�.�;-7� �	=ga�{���A=�붼ɻ�<�B�<JnE=�Zx<Q\!=A߼�>;��t=���<��N��ғ<z=��I1\;Q=$--�I��<�1��T0�<1��;Ac���b�<��2=&�����<e��<��#=�����B����<�r��	YR=��
�����\?�R	�7d�&YN�<�_=�)o�?��;��~ei��R�<]��:��:��ꃽPnh�ߘ=�f=�
��!�<�K<{3�n^C<�<=7�<��=���vm=��F��Z����_=lY�<K���<<��q����<d�t��Y;�qV=�2;�3��j�{j�������-=�f�<�!���;f���K=3�Y=���@�=�ꈽ�;}���d=W���R�S=�7��'b<(�(<D�:=U�<{Bc=��4�c�`���'=d�Y�Q=�[D=	6s�MLP=�����<W1=O�6�/��-���_��3���r<�U+��5�D���</=C�G��g��Rz=���L�	=	ש<���<��*��H�<!FO� �9M�c=�+�<��;b�l�xX1����=G�`���s�P�9<�Ѹ<]M1�c�<���}�:��2=(^/=�	$<J���e��/'	=d�/=wLM=Ʋ9=�F¼5�;C�j����<4�+��m@='�	�e��,(<��-=I��[���pI<�Bj;\XC=d+?=�7h=�6�=�;c<�g=A�f<�|F<��O�#�x��T��Q0����<f�J���<=!�>Pw=�=%H��������������@���n�c�9��zV���<��;<1]�<�JT=������><	�=�Z=
��Xy$=Z;8S�<ŏj�s>�;b\<&�U=#��;o>=߀u=.��;;�H����B�<�r<��缢e��^G#=�=�7<@C���A�T��$!��=BB�;�ji�6[�<o8�;	II==j�<F�=��=b��=T�
���D��[���2�<��<�0��j�<>j��H5=� 5=���<��=6P�<se=T+ۼ�#S��u6�`AA<��
�+��Mw�<xP�;�01��%^�!|=��<,�=3�ͼ@n����<uO�It輚�h�U�"��0w�$�[=�P�#�F��E}<0�<�7-=m�2�T�A���;#eU��;�[(<�Q)=1�ǼW��<`�T=C�G<��Q;������^��Ծ;X�C�����U=L��&�9;K��<8�W��ļHٕ<�����8���y)�lxz<�?��c������<�c/���<�1=$=5��<'KA=��-��<�v=O\�x���[�<���r��<�/<^��:�qG=�  �G�=ni�<(�*<e�B���=��1���"=,0���K<�
J�X�A=ɑ�;��m�ُ��0�E�q���2��<6��q]�<Bh�~X�$[�<ƕi�N��<yu���$����U���-�L��(!���;�l�=�l��L<�HL=�����3��]��Y8w��ƛ<��<��	3�<�<-� =�M��:�3�Ǽ�<�;%L���ȼh�c�[V�<�.�<�S�Sj���r��z<��T�;?�W<�ӎ�-;
=��F= �κ	>%�g,�;��0=�Qm<�>�a�L;��3����<��;�u�;v�o=Ǩ�����2=�bD�
�=�c�	=Ȕ;�k�׻���=O_��=A5��sP���<2@��RcI=�0ٻDo|=G%ռ�9+=&<:�aΊ�h�����<8��8 3=�ȼ�]��!k�L�׸�� Xp�_�'��+=�X����%:"�,?J�&�@�~���[g��<j�<(��uOԼ��H=��e�!=�B�<@U��z=����,=! �x����:<��!��5Ѽ� ���(=��&<�E=�I�ƣ�<���<&2;nQ��W,e��Z;�;�<�A�<B�X:�{g=�mD�S��=ΰ:=� =P�=�0����U=�B)=��=�8B�_?��6�;b�h��gż�S�n|�  <��C���Z=��;c����a=G������]�<��0=��>=�W��Y��[�<f��;�$p�/]���x�<� =O^�<�@)=-�s�"��<�$5�)��;Q��<�+6��ڃ�Q�%��[p��D��92=DZ=M�Ǽ��p�)U�~[����»��2=�&����Ļ����G�\�;=��q�o�P����:$��8��SO;y=���<�<˼8`R=�&G�|��u$=Jmu�hV=C�����}�$��=L�{6�h�#���u�yR���<�7����ջu��<�`��p<�CO<��!<F!�<��9���K��^s=�u�+�����i<� �/� �E끼/L=W���S��<P�V�9�5��*��U��-兼��<���������<ӊ=yb�<��޼��o=��T�z �<�Zۼ�u<�b7=>]\=������|�\	=R����=�,`:����>�b��e<nҾ��8�<�g<�;>E=�}�<�ڣ<V��N�=�#9��Q=����D�מ$=&U<�p= V;vs;��\��R��<v�v�ž(�yy�=cap<��b��K�<�b�R<�;N�o��.5l<#l�<�A�]�<�L��� ]���/=�N=���
�Z=s��;�n��O=�===�_�<��=�˒�܆�;�$=�� �����*��K��}��M&�&p����<N�~��H<;X��/=�&e<�hi=
'<��Ϻt:P���<�>��.�N�<R��:)y��7F��r�<RK='*���_<�6z�pB+=��8�$q7���T='�
���z�h�==G<61=l��<��R<�5=i��<R�W}�<^W=����A�<mc����z<@{�!�ż;-{=�
R���`;nh1<��=��L=�4�1"�<����h�h�6����q:=��9��`m=���<k-��)=� @����<2�ռ��N�s=��ļ^<=�=����=�;�-"����:��:�YL�]IM���<Vy�:1��<����m�㸴�v=� ��^�<\vټ�@��H��YDj<��
=�C;=��J=YL���IA=¼����>tR�чٸ��7;c=�����[=���D��ɧ�<�2F��Ӛ<��@�
�=y�5��4����ݭ4��`+=�ʼ�{=�L�����b{м�2v�ʖ�<�Z�<�Q=n�M<><�<rWû5`���28=账��4����<��<�"�MB�<����4���;�9��:C��1h�:�~M�:P!�����v=�>�<KN=�;p<B�*;<�����Z>�:9�7�`T�<c�=���y��<}B=��}����<ȼ<r�<F�4; �i<x8����=Õt�?��o$�:!����e��tK�;|<F��V�o���=O�<8�=�8�=G\=W�M�g�_��;=�匼_�<��=��*T<��b=���;kuf��Up��[�;C�M=���<��m:����?��
�޼$]�;��=��<Y�;0���a3=�膻�zn����<��<�c=1A:=Gcd�w�A�6�?�`1�<�pv=r�=Z��-x=7A]�/}e=��;[bv=�"�W�Y�2��[QG��/:=��<O�=u�2�hbA=�̼��"�Vu8<[�;��	��I=�w�3&��	=�(��R��<���<�V=[��<b�<=�h���ռ!�=��<*C^��=q/D����<ؗ�;�M��B�<0):��6�<�N��l%= T ��<���y�D�C����=�����?�w���y�}<P�e�x�I<�M=j==�8=�Q�<X�^�I|�ͪg9MV��K���k+=!��׸��hH=�.=�=D�P�-=�t����<%|=���±���ռ%;�X�{<���<�'�H�e� 2�ׂ��j0�i�7���˼�E|=�}�=F�z��<�=��һ{�7=�3=�Vk�%��Ѽ�.P=�4=��;y�1;	G��;��Z=�K���9q�<�
v;�����T;��<Ò���Zw;�ň<x��=�xz<@����!��F�9/";��<4�<��=mK��2�:/��1�=��7������
�H=��.��_�Po�<Y�=MD=+�&�,ւ=(a�:\�m�Ľɺ����[:=J@C�!��<�0e=� <]��<��k��Ի��<��<mZ�uť�]�X���D�A»Do<�jn�:�;�E�<�������H�:�7ߤ<�����<�]q�Lb�<9�ؼk'~<�T_��m=Lf���R��Y�="�,���<� =�\U��b�� <!w=�[F����;ב<Ju=RQ�*�F�Ȯ<E�A=AՈ��AS<V�0;%�3��xϻqJ==�`� ��y�3��<[�V=��q=��\�l<�p���ۼ
�=F�;�
0<ी=mS=��h=OU��])=A�$=|J��� ��P�໙<
��<�����U; �<;5_ <Z���ze�;F�<�D=��O=��8������]�<�S�]8�;���<��ѼN2E�Dv�<�t<+/S=��n=;3�[�'�����=���<O�μS$�WD���6���ڼ�N�<��*����;��X��:��u�Ϻø.=%~\�H�m��<�[�<.E`=�:y��I�� !�z&=�4�;L{�ګ漸=��|=�=hd��u�?=ut=���W=�/m�~$��m� ���<!R	=���@J"=��M�� 7=�/k�jＮ�Q���n�a� =!�[;�b=F��/=',��8�5 �<�gԺ�3=�-��h��tw�����}�<g0=/�;o�=_���́���t=㼠�ϻ��'\��A������?��<����Պ���G=���<2�<;4�	�A`=4f<mFG��>=�7�9��<89<�m�<їU<��<�Ż`P���9=8k=�� =�0F=��f=��<�Cr<?o+=�'��.�<�<� ��N=z����D,�����!(==���x?O<�::=}FP���5=�-9=�W=�[=�\�;۸S<��Q��m<��:����H�{lv=��5=t[<n����=����k��=����C=�I<��c��]=HJ�$�1<1�;v�<��޻�9�<�\�����[��1��I=�Z=� 	���r=������<��@��ἒЖ:�$.=Q(�k[X;P'f�|�M=C�O�~���ϔt�n弱v�=���$;W�@���<�_����7�v�<�¼;�=�(̼H�G<t�l=��_=a �ª|�����}ǹ���=�lD�Ȟ�<D�����X=�P�<�P�<2_X<3�<�Q�wE�:*!:���@=�Ll=s�R=�o�<�-=�G=��;��v�����:9����Լ�8�<��=�F�]��^��i�Q���J;#� ���<��U=�o{��+����<�C�<��>��ی��⁼󻔺A�=sx�E��;��P=}ܩ���=�#�<�|һ���p�h=��$=�s�<t�b�) ;���G=��7=7���5<��м��<�L)=>P���� �"�W�1������a��w|=�5=�;�<N*�.P]����<ݵ=�q�<�bi=:�e=�=;ؤ�mR	�1^�<�A1< 7d<W;D=&�:<|g���7��2�<d��<��<V����=�uM<�:���<W>!�2�ʼ��e��=l��$���a=%+�<�4	950K=�I�/�A��(!=�<b<H�=?<��O����<��=tMü��B��Bo=�����<lQ:�Li�@k7�-�ݼ��U�@�3�������i=�F���2�\G��0�<;�-=�,�<XIG���<�����j@=/�L���i�V���d�c��;�Lg�4����b<;�'=����3%<�h�嫼7߹���"�r��=�C���̼I�\����������,F��q=z�K�u�&��ީ<y�Q��c=�5E=ex�C���M�=�����o=��J���b=o��<A��o)=.�k=?��<��2=Z��<Ip�<����=1��t�j=��h<��<r#Ӽ���;N�-�L�<9üV�~�P3�A�B<��3<H�˼dt��yd�!+�;lsc=fY����5C=��<��=�y�;�\��X�j<,U3�u�6�\���Y=LV���U=�I�:�t�N*�o�);%ؼ;f=HP���8���/�,I���ʻ�<��G<C�=��c�A/ƼB~p���Z��=E,	�ן8����AC�<>�(S5=wR�^㍼t�{=�Ej=�T�،d=>�6=�gi=�<�=��[��\���;��=|��<�ۼ�K=>�<��O�h�� W�S�g<k|y<8�<k�#���&=r1��*[$��7�QpF��˅=��X��T(=��<��
=��=SE=HD=�n#<� A=�ы���=��D=-^=6Nx<s����<^g��W�=�EZ���%=��<F��<�Q�Ӕ���,=C��D=D�L���L=X`��D̳��
��2k�%�<A��d-�<��`<7y==�	�F�=�"<Gt�.>I����;�]�<�-�Xs1=t8X��	n�ն��s0ڼ}���vU��Rc������+=պ<�e�yf�<]�'=ui�l��Ȱ�<U�W=��C�A�ȼ��<��J=�P�<�t���:Y�nK=H8���i�@wh�<�=W��j��'Tn���h�Ϝ�H�</�e=Y�vM=;�(�<&��z=.�P=���8;<��Y<�������5=WM�}��=J3	����;{�_�e_7���6=�W���E��Sμ�K(<��W='���:�<D�h/�(a;;f\<qμ�z��>=#�[=��<υ&��~�ߜ
�^�e;AG�W`�<1��G<��<=�Q=D!��]ȼBE;M�:�'�g=.Lt���!=�<2v���2=M����<�w�����]M<֏j=��}<#=��'=��1=n6��e�c>N��tM=�mg=��=;�B�
ʳ�@�*<!3�<�k�"�w< 6a�l�N�.ݎ�I�=�N��X��+��=st�<ys����=^��;�#��!<�g߼R�P�&���<s$�\R߼u�=�E[���J�Jj7���=��<�S����#<�e�Κݼ���<���;bԏ�з��u=�́���<��=����)�<O�ݼ`���^���Zd���L�m='��MY�;��
<���2u�(�N��9��t��Ë����&��;CP=�˻���=�i=�p�:O+A=D!5�3�n�_J=a��<�ِ���{�c�=V�L=����������L��ހ;�Ǡ���=��6�/B4=�����P=N=(�P��"�<�I�<��U=/��:#(!�*?=T��<Ϥ�;��4�!�<c�r<��=}��:����h:=�z=�J=K��c&-�Y�9�Re�<$�*=�=�=d���𼍒�<�s�<��"=����ˣϼN����"���
����u�߻���GX=�ò<���>�m=�Gż}��;�����4=Q8�;���;��C=O���`�R0=��=Z�n=k�:<2��@9�<}n�t��<��p����<�"��R��&<��=F���>5���:����-?�<��=�e=�����_�7�[�Q=�<@�E�2�+��z��(���=�7@=���<��$=��;6�=̯=x=�G��@�i2n=г9�L���j�<�H�<��X�9�^�j������z�M��<)8�+0���`=^�M��>��P_�,1B��[=C�/�J=n�R�9rn�m
���b�<�7����.�;V�����GE=�G<<\^�T=<_Ձ<�^a�h�=#wǼ��B�==�[R;ҋ�<>�;<=C��<��F�܄��\`=(�!�2hS=(�¼@ �F�=R4Z=���<��a=��_<<."�<)�*=B?1<�x�w�鼫��<#K=p��<t&U�r�#=�8]��C�;:��<��C��kq����� Z=�$2<pB=q;i�0�m!<��=�
=}���8���ԧ��(���f=���=��F�ss�}I=Ld�:��<nx�Z�G��Y��b�<�a-=k?<�`>��f	��i"�#}`���:=v 	��$ܼ��ü��Q=�SN=�6N=�ƫ<�J�5i=7{=���J>{�| =d7�<~�x����<y@1=|�=��%=�F;���6l��B=����t<��	;���P�+�T��]�<+S`�O����5=H����0=�ӧ<Ȕ���9=�'U<�g��r�o;�R����#�=g�=�h>=I���0�K=���~ƅ��~F!=�6F=Ja���V=�I���t\��S���h<~2�<r�m<]?��C�;i~��e�T�X��.g<Xz<��ϼl",=�&����;*	�J�<W�<�ż�#^<�J��U*h���;g���A<��ٺ!P=崳<.�;	�<�+�<�����=���<�ܻ��4=5��;_ d�񹖼�p�9�"��=�q�������<��<�5[=�B_��!�W�M=��t=�
ػPP=�W�RV�<0^f�zd/�#�;=+W�<fr=��-<u��<��<0W�<IƉ=&o�%��<7���O��*I��O=eq=)�%=���мM��F�=p	=��;؎=�E/�Z�<_������<��=��/,<�+=��=>�컉 d���;��<�<-�p ��� =���I��֎��#��ɼ�̪=Z��]|���m<��л�%=#��YU<<�dZ= MO�z��<�Y[=�	�;M��\��1�V=(7�<*���~S��ٮ���!d<�>=����d=�F�<���<�b/�l-a=8��<�?n�1�q������=�Պ�p/;�3�
XL<W�ˁ�d|�Rn��(���뼫m�<��=8_-=G%B���I<[�n=1�\=t�P�A-=��-�,�����C��;ک;ī�� 7�<62@=��l<
�*�n:��%�^��y���?���
x���Ԃ9<���<��{�����:U<Z��r�l!(��U�;�*��Y�:�fd=�SJ<����t�<ܗc:��F�}E;iv=�!:�o��;��*��T<=�<��=���|������vc:s�5)�;83<"6�<��r�\��<�w=�JU=�IT=r��<K�J<6bϻc�N�u�=_�=��W�Z&�6)�R����:�Ak�pr\��@=��Lx�<b y����Z#��h8<�ǁ<��;��*=���<(��<OMK��G\=6֤���=�=��=11�<p��(�μ�豼��$;(�=��]=9Ys<��<��h����;��T�8=Z
;�U2��`c�Q�a�?�C<6(�<`�F�1�fD�<a=F� =�j㼣!������×ɻ�üq����'<�,=3T�}�����J=�>���GK��c�<��!��R=h�`=��̸>�S=M�*�g�u;�j2�=M]���f��薼eݺNZZ=.�V=^v=�����O�G�m<��Q=�h"=f8�I 	<�=�(��^�Qw�<�'=�yY<��ż�����{4u��Gֺ9�)=ܥ��:8=�A
=��<�j�<V\O���<je=U&��5�;�h8���<��(X�sHļ�=[BF�sOT��=���"a�<�R��=�O=��\=30ܼ�X�=ܟn�b�F=V�>���<�\.=b��F�v�9=$>��z���1=+�<ڦ(=q�4��d�<A&=w�G<�'�<�H��z<�=w:"�]��;�@���U;�2S�$�<�%%�WT=��S][=��b�1��;V�@=�D��rG�%�	=O&;��6-���P�<}�=��$�����Ѕ��`=+�;W��<O.=�w~�`O/=�L3�T'I=M�.����;Y�p�8�D=ɼ�Z=����U==��}���=Ѕ��.�<;�Y�֊a=~ܲ��������۾=h>˼0Is�o��i�@�F0<�F��j-�9KN<@�O�3J��W�������1�lJ<��Ӛ�+6�e�
��s��`=5�M=)e�D���=��+3`��#�KhK��dM��0��VY�<�z𼴴=�O:�.EW=�o=���;/�#=�c[�I�g=ӝM���:R]�<���!83�<��HM�<}�f����ݚ�<%RѼ�#-=�g��/5��7�<���P/��]G�D}=���R���G�ټ��<�/�]�V:=E �;~�<��%�2��<��<g�f<�=9��<}�b=iU�/���<q;�md�<��6�@�VD�<�6/<�7�V���m��~/"���<����`*:K[=w_7�Oۏ:���<l�3��̼�b=#��!�<ⱌ<�'��b3�<�VK�P��;�E�4;,�b�Y�D���E��<y�,=*�/�*�*��_tq�aP�=��9<M�-�3�-��>���#=	=[=G�u=�4�<�H=ڽ �r�<j�<oZa=��:��:=����x��!=��q<�_6<ۦ��z0:=�W�
�8=�S� �A�[6�<f�=�Q8=�W=fz��I=�;=KH�<�H�X6=�$����=9�=1.p���#�9��8����ֻ���<a�<Z>N�8���\���1�O��<A���0=h�b����<1[;���;�0^<�g��z8=�."�I�[=��<t�˼�b���G����=��<�׹�1;���<���:�_*=��Z�:�m<Q��=��=�[a�s~�<a�U*Ҽ��l=��m�)4���k_��\C����< 4C=7޽<L�^<9>�&��<�d?�A)(=�t&����}83�s�B=y�<g���G=��C���c=#w��V����<n�.�	W_�t`�)q��]0<t	8��=(�9=��=�N�<͎��(<馨�� ��@hV�����[=:���V;�}?�YM�;�����1�!�����	G��p#�h��<��<*}��1��<ߑ[��ݳ��:;��;�I�����V�۽�8��+�R�%=��l=p���8=�]<hI<���<�_����<���̜'=#)X��ǰ�-�< B=�9�<��=ҩo;D�b=�ڱ< �<���<ft��AG���h<>���	=���Hv=,�E=�
\�`��;	�=�<JX��/!G�"=E��,
0=�Q&��=Ӽ�(��q2�C$!=5Z���A���@<k����,�U�x=��G<4��<k=8cS<�����ɼM+<'�<
�!=�랼�)&�֞=�͐<�'�<BM�<��0���Y��P�;\L+�W��sX�̟;t��<9њ<�=E����b������1�ڢ:�S7���a=+D=�N'=�A=�h��ײk�63=�{�^%��CH<��;%=�",=�1d�W�M=�<�;d��h�r	=�@<=�K=�덽��Լ�6<�����= ``=�b\�dOx�]���JAǼ�m.�	�=��
=Hʬ;�p�Z<���(��h߼U<c�ߠ�<��|=�6�?jF���������G����Q�"v}�3O�<*�R=W����^*=z=o�`=��J�F�ͼ��ؼ-�>��s�������;�l���=�o�:#��=����BX�#m=�A@=Z����r=��"���&=�j4=��ѹ��*?&<��f�@�<�.�<�`�:H�^��R�;/��<ⷻ�rE=�2<���<���'鼴~=�*=�]���ۼ����b�,;�2c;�m&=���<}=��A=R	�<���=l����=Ln9=�폻@A����;��)�82���o�=��U=�E����� ?�?������R�<�e���E<T�T�?�+=N,}<d�r�<[�O��%���<��<PT�<�i<�`h=�u���=i�/��^���=.�0��wR��()��3=���<��k:�ᴼBz|=�?=�)r=�W*=7-J=I~�<��!�6J3�g�d�������J��<��e��o����:<��ּ�Ld<e$%=�O��	5�ƽ��Q+޼{��(�7=�"�]0�<b�:g��;�ǣ�8ļ|�G=K;V<�<����; "= A=�c��'~������<&��<��������-�<���;NTI=�ZV�5��<%�	=}�z<�������QY=���=6��WD�`SW<Z�ּfu�<im=�d��מ<t�%=�=DҼ�n==��;�'>�;O<�	�u����̼��:���<�h���<-4 =\?=w�@�ż����Z�!�7;T!��)��;��X��F�H�g<�Q�;��L=�<k*�z�D�b�<���1�K�H�l�<�+μ�!�N&�;��i<�>�<����!���\<e5�:��T�ݼ���/\=�2 �)��;��-=��λ𱳼}��Մ[='�üm�=�~���M*=�I=1�<>G\=����~��<KD��5�=�j;-�j<�A�<�P��sL��Ǆ���U=�@<��:�Ő<r�ꓼhP<�� �X�����G=#:�<W�ϼB=;˻�/i="��<��<*Y@=��˼�y
=Ǯ(=T�����<�6<<-��/�<�`�rܪ�n���-4=�T8<�O��y��<Q)F=�u= ��:�B���;�$==�� =����KB=�==��;=�
ʻ`������;1=t�K=M�:�<�W���=���������O��(_�R=Su�;�XM=͉=@:(��n<�钽31�Ι�����<䢏�hx.���:��� �?�<#�<[�+��!� x<�і<���8���������:;�m.�=��H=��=J;{�A=~)���{�<�=ԁ�;��N=�͒���U=>.��� <@��=ri��Z�?=!0=�(=U�9��"����<���=$Ꞽ�.+�M'�<�i��A缄�l<�U�R%<=�T<=3����s<�/E��o&�D�<���;�/�s@ݼHcL=܃�������f�'���M<>C�<�8$=��	��FK��U��^=�����{�<	�.=�=Լ��<��;�F�;�=�!h���;,��=1۩;M	h=�K�<D{�����
;8?�<j�<�F��ݲ+=�ټ�:#=�7黽k��ޜ<��ټ�p�Wg<�?1���k=���<G=�K�<U1黈.=�l=X�L�Zg��rTD=
�<*�1=k�9����:�qZ<�*��$���)H<�C�*[�oX
<U`=��.��O�����1�#���'=Bሽ�J�<�:�<�j���*���-<��=�x��4a�b�<���<f�<p=�3=2�<�<,�<mLԼZ�;��W�V)�<�n=�\q=i�=<��=��;%E,=��<%�=��$=�e1^���<� W=�;�<���<$�����=��|;����
=s�q=���<��4=㟁=|2=�+�n;��</=8Y=�޼��o��Z=y4u=�<��<m'(�z}<^��x�=�U���B�<�S=��:��;��q�<��<	�r�����l���$�� �7=��U=�����<k!�A$�;�ޕ��ټ7�1�8�<.�Y=�J�;k�z;��=���<���=Ϫ�1�ȼ��A=+��T匼t%<�%�9��<��ռ�(=�1�<~/S<:��<�u�=�n�<3�=� =�0<�D�����F4˻y�e��+�<���s;���b=�)=��=ν:=�ļ ��PEe��F���<���<# ��4�Ð0�携=�=]�P���1<�_>�K�m<�R�=P�=�۞��8_�'<=�.<�"���[=�;�<��4��@9����<����`�<\R���{�<b��<Q�U=n�?�=޺@�$"N�N�B;Y=h���dj:l�T<�56�v�Q����5�；���#=\�#��^�<Dػ�*��<�<�[<,�B=�>�BL���E<#WW��O<k�'=�<D\�� ������M�!=��
=S�����<� л�1h��!o�4�V<q�������>ż�Ӻ�=~,b='O���/�P��<��O��;b��<$����<��[�N'����w@-�M�<)Z=ɢ<9�:���� 3=4��O���w�<%A=�==��J==p=2>V=�={9<�� �X�<v�=Y֒���V=�B��'.=�c�<��n=z5��=	�^��=J�@�3�1��gA=����	ż�����S#���;�ɂ���m��SW��"E=J�&�2O%�lQ=��<�5��w&��=�^?=� t=���<����h�k�Tf��}�<����rD=b:ӻ[(���,��WD=�I�<��D�'8~=������U��}.���5=��>=;�$����9,��:x�终h���-�<.q ��"������V=	YJ<��(�ӿ�kku�A�E���o<��I����;r�� ;�)(=%^�<~�n<:^</Ӽ4}��:=ߵ�<g)�A�t;p��Tl�<��=���<�W��� =�5C��F\�.�(<�]�<!�H= @�<�	=��q:و������<�40�kN=qQ5=�T�+��<� A��1~=�_>��G����;
��;{/��RN=��4��˅�D�Q�����/�6���@���/�L�=�W�<��O�<�.�������<#�+=o	< $=�t�<��=���S�컩�� �2=��'�J�<y�q=CF��U����<)�?=
�<������-��<k�<?��<�VZ=���$�	���V��9��
;��<t/��xm=�J<d�>��A`=)0 ����;�BL�	��?�V<)8b=i�-=S���%|<��=G����H[<�� ���k�6E�:�;��|�'="r���)=kҼE�Y=��<b;�5>�"�e=QHJ<��8�Qj=�X*=�WN���p��1�<<0���d�9Y�u�b=����4��kE=��V=�� ;G��r��]��;�S=�G��v#��<j=������q=c����d�2�$�]��t�5�^rN����v�w=�;K=/�����.���>=�i������q����(sd;��n��5�ç�=��=X�Z=��=�M=�A���
<��=�"=�L=�dQ=���"����<pN����x�L��(���������p;qc�;I$=�|=��;]���n;���mP�� ��<JO6��;��I=
��9�����tY�<1LV=����c̼��P��J=�<׼�+<���<�|=���"G�<Hs���z�<M��<߹�n�O=�C<i<������<�<�~=GF��(<��;#�<K���=��4=�(�<��%�u=�9�d��<�JI�@��<�+�<���:�`�<���<��<��<�an�V�8=�����/<vd���ݏ<����4��Mj�)���<.�-�ʯ�;`_I;FU�V��<�hr=��d=r��:�V2���C�K.���E��o�:�l=@,b�0�=�ur=qݹ<��<Ne�;>��4m/=�=�6�����;5�=P�<���<)��z�B���<cY=�.A� ��<�I�#�9��8��0=fv�����M���|����G���!�_vA���	�W�u�9�4�S=��;(j�;�f�O�<a��<��6���<~�8�)��Z� ��7��j�!2=c�]=,�VZ8=���7Y��<�;8=�������<�:��ny=�J������^+=xt(< *�t��<�x&��r2=�a�|�r]=��;��$=�b��_<��l6��_�<HE��,�%7)=пA�C_O�VM ��Н�T?�3�=ȹf�������<Kx=K;�>웼�<���:���<�ZG=��:՞����<^�D=�$^=}�:|y=��8���Ǽ�x=���<��<�X�ƪ�<��h=��<��=`6�<��h�q
�<c���" ���r=;=���<���>N=xK�<u.���� �~;�=� %=݁׺�򝼥Xu=w�a;D���=Y���v�����=����.�F�`�����'�m<7H=����&o;<���;��=eW�<�W����;��	�.�5=<4�<��y��f�<��B�d�RU�\���.?K=�ޜ�)9=�n;� �D���<��,=�d=GL^=?5D=Z�)���=s��:�6��7��;�L<�밻Z��;i2�<��<�d#=��Q������C=Y�O�qA~���`=�R�:�@=�&=3#5;7�=�Y����<�t;:��;�5<��<��7�q4���Z;<��M='69=��=/<��6�L=�=*�="��� �;=�=� �w�2�O �<�N�)�!�	�P�<e��R�;�{t=���<S>m=R��<cH�<	;=�B=�-�h0�<�*3=� �<�����@�>V���z����.�#��VL=�4L=�u<�.��N̼�Z
=" ��3"�o=�;/&����<��Ƽa�<YOw=��9= d<څ»/����ֻ�ێ�]���̟<k�Z�m�J��D���O=��ͼ�S�:�!�<sI=KQ����2����<�� =�i6��3C���뼂Aڼ�f:�N��G�7G1=�<qR��a=2�=J�3�ue�<�a���<�V� �ڼ���;��ټ71;�=�d�L�^<z��<��-�ǸZ��N�:FI�<)KQ��5��A=�2�)=z�<N=2��<H=&:T=��<H��<�0t=7�ƻc�"����*^8���<er�;��}2=���<z�'=?GH=�����R=���:�
���J=�d����<i��<�#����<h�^�?� =$d.=̯;=Eh�d=V����^=#쿻����W'�sl	<Ƌ<�뉧�2=m�^�y��;�X��>�<�W�p�����|0�S6K���H<�9=hB2�xѼ,9����D�&=��<1�$�vd�Y�I=]��<�v���A=b�F=����=�I='ۿ<<eW<�����X�00��x��<�&��<J�f)���<�Ο�F�m��'滵C�<�j2;�D��j�/(�����;`�=�E��N[��%�6���������B��'�ͼ?y2�u�^;���<�2[�FK=x8�;q1��=�=@�0=L(<��2=�צ;�B���*E=Xh)�I�H)=7䓼���]�V�����vм�-;E[%�,�M�@��ɒ<��a=pu�j匼:$=k� ��X�PF��	�><R"�<n�6=fy�<ӌ�<$p��%˻�M�<^�8�#rW�b�=�O�<Z�@�%䅼���N=-�W�Q���(=	�<�6Z���<�Y=�>�<�s
�mU4<�bA�q_=��A=�=�;�4�<���pޣ<�� <"�&=f�A=9�]=��;)>���A=^���_k5=��z;���<n�C���;���<�>�w^V�	8<qX�<��<�KE��z�<|�<�O��==��W<�?'��$�Tm=��=�]=H2r=� =IYż�� ���=���<2�=%�<�ܼ��!<T*<���<���<�I;�g�EV�<'�p=Xu{=!�!�>�@<��
���[<�aȼ΁Y����a,�<2��<�,��z���弃�W<S`����@=��X�94=�ֿ;~�=bǁ� 9=����$�H=w%Q�	=~�ѓ�;䉸<�퉼'=a8?=!�F=-G��
��<w�g��(o�p
��-�����<<�o=�	;p���:�E=<��<n�I=�B=�Ψ<���e�q��ݻ.��=ˈW��5<T��2��T����?=�!=��8�>I6=ʰ2=�$��~�;��<�ƨ��m4=@�=���ҷ�#�<���;�}M��y:�$~�8ݛ<�yQ=PJ:�M�;cy�<r�*=[��[��Vu=�>};��=v%4<�:�A/��ʱ��Ӷ����;����j8=j��D+=H��u���9��G�=�Y2=����/D=c����<$ 
=5�ی��`@=�p���<z�:�Z=<�<��@�Z1z=��S=��:9�4=�ro��@=YR7=3��<�@O���?=k�v���/���g�'=��
=��><�!��z�� u ��(��V^=�y[�����Pu��i���Z���/��V�
4�; �\~*���A��܀;7C]�X
��Z�2����F�Q=�\w��9g=�J=�kN�/�#�Q�y�=|�d�w�S=��?�m�� �����t=d`%�$��<�u�=�@����,<�x��#%���:�<	�`����.�D�9�}=E����.=!>���F=���L��<5����e���Y="�t�1H�Z���:>���<���f-
=kI��A��0����<��<忞<�,�(=�=�Z==�ܻhaw���i=�j�<�P==�xE;��<=�,�C�d=��3���<;ʯ ��굼Y#�j�=��3O���=���<Y"��=v��<o��<��Ӽ�RW=Ud =lb��#<���%=ܘ�H����6���ӼL�d=�E��̓���<L�O=�d���B&=�� <�28�A11=W�C�ЦY�����*=ȡh=��:��-�>��H̼�_�<:,=F��<�H=w�p�4�<�C�;�s<0EM�ǈM<�]Z=�5>=.�����|=b�6�c-�h�>��Ҫ;��������n�<��ü֟��OT=��a�.MZ;V�^<DXk=j�=�j�<���;�� <���L�<�}<V�oBT=y$;m�<`q��������7`d'��4=�==x��<4Z^=W=��5=����Q�o�Ҽ�&=8(�=��
�<���s�v��4b�Z1�����x�<+p2=�P*=��<��<�$N�K�<�b�;�(,��p��%��<�Ϛ<� ��J����<�f�<�(�;V$r=�!���V=�/�~M�y)=�:�b=gVC=ݵ�<h�c�=��\K=�"���b�=���2�<�`�<# �<����.1=݌-�����S�=�TX=r6����
�8b�W�b�V�<v���A`p=�*��u4=�R�<K�?�Ab���0��(<3I�<^�<� S<�	8=_n]=�+$<l�$���;90&=���1;5=�\=�{�<<�=~�6<K�¼]穼#B���=�7#�YS	=�;�=L/x�8����%=�	�dE=���<9�K�[��p�L��ZZ�a(� ���9{L=�^;=�5�<$[�<dڂ=��=񜔼��i���k<��	<�2�<I��;�F <p��<R�y=z�7����8;<����1F=�����h:���<��b����Nb=��K�ܘ�In���?4��>E=�C=Sic=eͺ�N���T�،=��<� =B�U<~?��7fy=�!�kn�������,�@�F=�E=�(=�;�L��5��<�K�U���rY=Wj
=�Ψ;��;	5;��F��;�<�d�<72C=����v��=-D=�"D��<���S�<�'=X�s=x4�<m6=D&�<�-=�N=�bg��H�:���;7=��=��g=�¼M�4=�H=���<H8��=�`��3l=6'ĻM�=��@�F�z��]=�Zʼ� ��x���N;{>��d�����D�=��Sʖ;ו+=#ڼy@x�\��<4�;UV�<��k���=�����?<3R=���"=��\=��<��;��:�Ƅ�<隂=�=�*T�_�h��}���<���W�)=��;	0<A�=;�N����Z�<�E�$�^�i1<^�Y�o�Y���I={%���B_���;j�����küԚ�<�Ů:g�a�u~;Q=K=㨠��	=ǟ�:���UG�<�鑼�w=2D<�H0��K�9p7��2���m=O�\=�S5=�&<@�e�����~H�<�z<�>X�;P==kF��<�~6�C��s�j=�Y= ��<��:R�<=ߧR��0�t�<	C��T|�(z��3Q=C�<]5;��-�/�ּv�,���H�D�<����0�Eդ�nʨ�GA�<�tV�<�,�z|=�E����<�t/��b�_��;2��<���C�=�[;y�Y= N��+m;n�u;7:�]=���<��i�)�:�� ���.=�l����7�o�.�l�F=.Dڼ��¼\����o;P2S<)�����<�=F�U<�';=�I<�n����K�N���=����2��:�S`��#i��f<�a<<aQ�2��<�Nd��A =�q= ܼN�;��u<������<�"N;�Ƽ�z=`i�_^^=�C�<��=n9��(�0=��=2\+;i= =��~�eP���;�ty+�_z	;һ<.zZ=z-���"7=46�����G׼�3;M5<�ac���c�3�Լ���<RL��h�x���G����<�9��A*���[��5==h�H<���Hp`=%&0=jp5�¼,��9#=
��<3�I���.=��=�gK��!=�}�i~�;e��=<
;���;��p���<$�={[I=�53��p��Z�A=��-=l�Z=l�	s$��-=K �<g��<�W!=���K�Q=�¥�~�ݻv��W;��
�:S�<�/�<�˼�Լ��/�jh:��.=
���Z� =ݖ߼��=�����c3�M�� ���򒽡������<��(<�@�ý��1Y��ת�i�<<p��嗙�n�1��Ә;2��=
�s=qʼ�c�<C����(=��V=�h=d�Y=-+=�Jf����m��<�����;`������1��zEa���{=�����E�[	m�� ��P�5��F��^��91�i�*A:�l�&����l�=�x=�o�g:?=;����A���׺;&���<~����>=|Z���`6�{��<�T=��d�1�<ɪI�/x�;̦G���	�c���e�=�>�<{D=�'���<<��L=o�#�i8T�: ��1=B��YZ���B�FS\��ʨ;Y⻤���.�<�W ���X��]A��FZ=��J=g�j�7��X',<��Z=փ=o2>���;=�<��8���;x�K1=�R��$��ؿ��
qN<��_����A��<VY�i���<��<�����bR���;���;ϭV�E�}��g��8=�
<tg0�&�\�!�/�wui9l� <S�g=��<��<\�R=`E_=�jj=���<{k�<��
=���`���6a���A��.�)ن;ku{����:����Ѣd=��M�A��<��$�%�T�=�S�<0(���=���0�f?���B���f��u=D���5�<��6+=0�.=��=LX�;��<th=t/:<�
`=���vY�<�	}��5=�=4�=�������<�k��f) ��:ȼ�S[=��<ӝS=F�<n7��AZ���*=�#�<5���N<Y;��T=�w�(ͳ���j=K$=�ʇ���<�@2�� B�.�U=t��dL��p���Y�tA=�$=&�\=�׼w�q<�u��W=�-�<!.��d���ԛ��36�q�[�J��k<X��<=��<�r�I�<���<<u=I=s���:�#=;8/�<G.�o=��"=L�p;�K��6���;U����q�<�^����<��7=�뫼�巼�8�Ż��~��<�NM���;�^�;<�<�;�;3|F=l����伦P=:[�<�@<-��<DT;;_g�HQ�L�<"��;�S7<�t��XU��e}=�ջ�1j=�Z�`U�<U=�S_��?��W��������Y%�(.�=Z�(=7�Z��z��hl��&=㣼<+TW=Lh;=��p=�I��H
=i�¼�2/=�{=�sd<�Sۼ6�0=t�q�� =u?u�15�<-���}M
=~�l=R_�dSۼ	�;�}'�u]!=Z�B=Mq=B	��<~�I��QR9���<~^�<��;��<�F6<�ԫ���Y�.�"<�.�<wʅ;�8ü�=�<�<g�ӏ\<�����s&=�;=�X�<�r��=���m^���w��a�P=Z�;��FA<n�Q�0G��I��<^
�<A�Z��7Ӽ�	w=�I<�Ҙ���;5��<?�<g���eu^<�,�=�:=��f$<[w�= =��><�*I=��ya=l�>��᝻rA�O`$�o� ���J<jE=(�y�d�*��&�=+h��A�]kU�Ť�<n�%1#;�<(+����==ܟ��^s���&�;<1��gJ=��P�2\w��ܲ<��˼?��=X�E�eB ���ݼ���<�w=�1�<Ĉy=ү���l���p(��ݼ����R5�s�E77=>̼�q����=�/Y�~��Vo�;�އ<�e;'ܼ��z��~=��U=�E0����;ý��Ј�<HD�"�<�^��z���D� Bѻ8а<Um�<�����U(=�2�w�<����;�BR�<�I=�.Y�+/	�l�=�=�=�# =��=z��:�j=%䅼��R�ԟ���c=c����L<�d:���<R��(�oe>=���F�<����I�}���=�}�;�(=�Rr��~|=y�<�<=���=&1�<	"~��M��du�ǖ7�\�7��-�����=�Ë���ټ��v�>��`��X\�Wy���/ϼ
;��^?4<��C�;�7o�+Kq=XF�<��o��.ٻ%=[[�<ť=�n=�
=@�<���yk<_ �<ޙ=r�U�W�4=�6��祺���������A��=eB=�9ۼI�μ4��<P�.�A7"=4�D=�x=����<(>P�y�"<�s-�)�켸�3=,;��*��4��f�r� <�!y<��:A�=l���Ǜ�Ge=��=`V<;������,��<֫���=��;��(<D�;ɾ!�w&J��e5����<��#^<f֥<�˾��f�<����ڜu;@O7<w<	�:=W(k=��N��x.��B�×m�k�$�<�d��=�>�2:�<��<��p%=g��<Ij?�re>�Q�<�ZƼa�$=�_q<8�B<�M���E=�l=�S���Շ��`ι��0����<We{�D�l=p&��&�<�2��k�<�ұ<�C$A���M�br]�tdC��|2<g.�,G)=���<Ǘ����F�s%����<��I=� ��IR=ɮ=�<%=K�^=�a�<��o=�r�<��8���=f�#�0����� F:��"�,{R��$��G�G=��b<�Oy� �	;��)=��#���~�G��;�F�������=���8��n�F��M��~<�G=�U=����=D�=���;F��Y;="QF�g�5��J^��=E��<R7�<]�;=$�9���,;�. ��l.=c��;%&-��R���C=���qV3�EO=rj��b��F=S�<�e=� K<xJ!���<��#���[<�k\=l��<����d�1P�<��<d_=��F<:+U��M�g�V�ιg����X���-�<�j���<�AC�w%��@� �#=bz�U�Q���<9m���<,�p=�����&��3�=��x���<&\.=��/�r}a=��2=�ڡ���ՠJ�����S��R����j�l���<)�V�qw=N0�8�5�O_=�=��v��!0�jO�<t�Y<D�A�DJ��}k<�ԙ�7?<��Ҽ��]=J�<{���g:��?����#=q�Y�6�f�-=P�!<�І;׸/��		=�6:";�:��/<q��C����/`߼p<�fӼ$�Ӽ�_�=�+��QW<�=뼚r�<C��e2"<��9=�E��O��YO�<i4�<^Y=���wb�<���<�_4=[��?,;�mN���$=�/�< ���D�߼ܓ1<�I����!��D<����V�}=>�ݼ����,D�r��0�A<z�n=<�f��A(�GT�^�U=��0��R�<O�~=�1�(5=�s�<]���:�y:V��̼+#���=��+�g���:��X<C��=ӼP64������`���De�H�L�<)�x����ﾼMf<!��:��<�L��N=n�<�%=BNʼ���<|�@<	«��3��Ä</Wu=�[n�.6Z<�Z�;�a;�N9�x�g�\�=�2=�!��t��=���qm=�q;�+Y=����u��<�I��J8�8�~ռB= =Qx�=���<K0G�i�I�ߊo����;�c7�:�.=�<�ռ���wF\=� �u[��l�<���\@�����'v=�c?=�5�FFX=��8�n)s=oY=!M0�)~.=TTK��F8< @ػ��3�~3���=���֩<�����<�%=xiC=�x~;�<Ԕr�n����P����b�	�`�I�C<G<�����q<e���I����;�:3��/=�J==�θ��W���m���S�m�<%d�<|7h;�<=��"��>�=��4=��źm��/�����r<�Ϛ�.����>�Gn��΄����j�����ӻ0d����^���ּ�mW=�s���<�����s<h1�<�?̼)S��q�g�]@,=a/�<��3=:P��"=ZM;TYG�7�M<E*�<��<P�ļTs�<^�.�.x����<�c�<��e=z�t=kr�c#�`Vy��G�<���2d=�$����5l(<O$�@������[ּ<�4�o<ύV��y�< Z�<�b!��-Z�Hi=;2�<��<�z���uo�Q�h��9�<��W=c��PB7�>�<�O��Wݿ<�>6��	�<�~ڼ&����"=�[7�U�=Eu�x��;|)�<��Ӽ���<�d�5Q��`��l=[�=�7<����
{>�n�>=о��L�O˼b:E=�;ȒX;J[m��c`���<��u=Cc�<�Ǟ�K��<y�!�Fۀ�櫺<���;���x�
=�y9:��4=�$��l�ȩ=\'����]���=l��<��1��1��7�2���b=*?�=�5�?Y�<w�o��z޼�����:E�Y�KJ=�F����5���aۼ�=/��<��=�{�����!a��mh=PQ	;SZ����u�[�F;��=U==�0=A���%s������y=�7���<����6U=HV�$��;��==a�M<��=$c��==XU�<�l�<�g��S�=��;���<�_u=y���|=�ō<�PC=�@=�p��"p�7�<���=`=7<�ܩ<�A�A�=᪋������<��ɼA|�<'�l���=��<���<�-	=�P�u� =a��<3�N���k��㸺q���s8w<ļX�Ԍ�<;��<��������;��;"Lh<�8�<��� ׼]��<;갻��/=D��<��<����*=��a=b�V�T6=�P =��4<�ᇼ̖=�����̊� ]⺒-=]��;A�k��<��.=�a =������/���4=��=��9�� =�`��=�kc=S��<��<O�5;3F\��_�< l�Y�X���!=<@��_=?�<|m=��<�q���6<�k�]ﰼVv=B��;����O=��<19<��o=h��<{�k;-�P=o�[��+���	<�&�<d��r)�<�� =��;����<|�b=���<c>/��@g<���;+ZG=R+=@'�<��<����<�ύ�:��<fF�<�˺D$�<��<�h�g�i��m�<n��<2��<�߉�2��<\^2=-=�=� ϼN!��ih<(�!s���f���Z=y���f<9	��B>=��	<�X������l <�Yh=�"��+
���ފ<:�<����L��ɼ�	��9��]}<GO_���==�Y�����<W8�:s�W��=8�<4�OyI=�ټ &=%	=AH��	 �=3�<<c�����m���c�����<��0�F�e���!=j��<�#%=4�;$��=���<IY=+��<C����=�YT�n��<À��@��\��ʊ=[���PL���H=K=�=�1����󤊼��=�V����<�^=8<$T��?�<՟��������H=AV�;���<܆9��=��<�9=��=<�7R<���<��u���_9R�B=��⼷5x=ۿ�92�<Wz;愨�J΍����<ݵV=!�T��7*=uI=k�b=l�O2=�^3���-���h���X=��<.�p���Ѽ�
D�kY���S���9��]=�=p�2'�<���6�X=~c�<v�.;�μU�=r/�;��~=�ᄼ�Ɏ<r�=�;=�dN�E�_�r�?�亮<��2�-�/=�6=�v%=g�߼^#�:�G�[G<�e<m*�b��ɦ�D�<�T =h(��D��S<T��(S�вp=��</6.=�����:n�5�ͼ$=�`D=�żԶ�<�N�*=-!a=�$==,k��* �<>�	=�.�-�6<��k��Rq��O�<��d��;�������d��X�7�;���<�D������1=�em<��w=��ȼ�<U��<�ꅼ� �=�ܻnL4�Ht<�#<��=~g:(��<>�W�M�y;�D�6�����;u��H��v� ���.p=�=�V�<�<ޒ�K%��#@��Iq`=auW�{�R<�����I���@=(��*9�<e�@���^=����;��Z�ٷNp���;q�$�W���������CЧ9���;�&A=Œ[=nU�G4=����.=��<�U7�MiS��6�&d�ԩ�;��8�x�T��w����T��{2��~*��Y`<o��<67 =��b���k<�я���1�g�<A�p�[�B�n�u��8O���5eI<�A =*�;{�e�:�V={w0=-�j��|#=�9�<��H=��=�\�<Y��<ܸ<&�=��fQ�<x�^�������<��I��!K�8�}=d�,=J=
������G=$?5�v <��<Ə���{���G��HA=�3=�D��uV=ޙn=4�:(]<	�I=L�*<��$=)�:�{��2���=�6P{<�kO����:�X(=)Z��n
�H�<O�<�X8�26C=�ur�,Ў<�;��=��*=�lv���S=�*=�g��
M=׈�9J�A�c׼�<<>��;��B���+<C�<���<�2'�B�<�l<;�<5�T��q� �	;��S=�`=�/=k�E<�ٕ=�j�=0?4��b�������8=rJ8<�<�? <��L��k=lt��N��w��<��r��%��J�],5���s��g�k���=L!��E�<��o=0¼��>�x/X={��<g�-��v�����<
-=�z=d@�&�w<�	Լ��O=QtM���{�>�5<���<ҟg<���<��(�K�0=��<? ;���La=��.�7��1��f��7=����=�����;�B=	��:��V=�GA=�� =��ļ������;0�r�̏G��|<Ɓk���=yvo�)��<�ߎ�wV��[3��n��t=���y��Gἶ��GȖ��fG��i=W솼	(M=-j,��2���=Ŵy=�����c<i��<��*= ��8ZM#=�m$��G8	���<��#x=o��ظ���b�<gh��9�<%;h<߉ԺK(�<�m/=�5��E�������Ȼ\[U=݆<V��<��B���r={�<�{<DN<=���<)n��1};�4� ��`+=�p=�y��f�V�?=˩8=d��<�^�����_L�<�W��&s)����<�T����24ؼg�F����<}�N=mw>�B�#��	l��v<MG�<�l�<W5��y.^��g�<���i�N=�<��8=&�ټ�Ԛ<F��<V�^=�a�˖D<:9�< �=�%>=�Ѐ�o�N�����|
�<�e =���=l�;­ۼ���A�<*�x�ۅ�<z,r;
g^�E�����<�3w=��T=�@���)=��)���4=6�N��ć<j\k��<�&�L���a=ѽ�r��x�<C�g��s2=��5<��R��Г�6��<]�i<Y�5��`=ط�<F�=tcl�[�r<���<p�����Mrb<�m�)�`�d��:x�3��e�=:���-��&6�œ��XWB�m���a=g��<k:5�݊��L�IT=]�1����<���A��<�n������(����	�Ux��(-=��N=(lƼi<�=�I���@;<`#�;�O�=�HB=V-=�����=(�$�	��N���S<$� ��#=
�v��<P���#���˻�ɻW�A=���A�<vH�<T��<�hO<�<��(=zl�uu�=��=��$�X�=�9�;�[$=�2<�*8=�7ڻA,�����<���<��*=��=�@�=�V�;��;#��<���u��<�}2��WM=�r=O�+�T
 �Y򼮤=��(�p;�N<�0N�7����_��(=��/�����
U����F<�?��린��s�z�=�x�< w޼"^��c0�<m�ڼ��<�n��Y=�i�<vD��c\$�������c<��~�&�t���<�8=Ԓ�<�!]=��ܼ C\��������$�Ҽ�O9=�<��<Y�n��R=ɋ�n�5��HV=��D@��g��j=wR�r �<�M�VI=�iO�$��<80߻	��=Ko2=C
�<��=�#{<�;Ѽj�_�1���6=�����G<�;vh=ip=˖N=ΒP;z��<�Á��=��hD\���<��=��;3I!���<?�����RAV��	���B��bT��C�v�"<~�ܺ�f<�U=�@������-=���<X��<�.=� 2�K{��zD�<�7=�os������<1��n�f������o=��]��W�ԩ�<ԑ��G�<����[�=e��M�<c�X�$�=��U=�[��i�<�7�<Ӧ8����<d�O���`��+��o���_��OW9�Z�Z=��H�`i6<Ԑ�<t�Q�l	��~َ<N�f9O=$J�<֖��#���%���˼���<?+=�NI�a�L<�s-��d*<�Rv��xg=��; �=}U9���&<$|���=�'w�e�=š!�p�Ż/=-��aQ=-��`l=��Q�+ɟ����5�'����<`�$=#`^���<p�<F'��=(�&�	M���W�eW�L?�;}�
=��<��<�����w��7����<*�_;�̏;�t�;F3���U=Tn==�+�}�=��d<	���Q(=PA���%��(P=�a<iY˼�!=���;��H;ď�;zB��-=by��ʪ�	��-��S��o"g������*=��V=�׻b��,d�=�CU<j��;��.�=���=�$\�Z�G=K4�,]=d�=��)=O��<t��<ll��6���<�<-��;_;2�z�&���<t�o=%=��������<��#��}s�b�3=�P=�4=_��� =�����5,��}>=�Ƽ�&�:1��v;�<���<�Ϙ<o3L�<����Q=q��&=��qc
��ۜ�X��<Z�h��^�<�'���	�ȼ{U�<��*阼��#�I��i���M�����B�1X���jϺ���<����*-�@{�<���t׻���<i�w�7��V���R==�K���<��D�Jښ��0¼/Z�<�	Ҽmo޼c���n���X�<�g4=uL�<^M�3�;���;u�4=�&:<�ρ�����aF==�NE������7=��	=m���f�=p���=_�U=��#��X=��;F�����:&�Wǹ�M˼�ټ�g=����q�Y�5�ID=4i<�^-=Q}��M�<^��g�<���:s"ͼ��<��<r�(=�@��_����<��y�Z =�s=tr&�Bٍ=R	�6'=�%H�<�xż&^��}��:���5=ݷ��V���S� �H��R�}O]=�@�;��l=��%�yU=��<��!<RU=6$��z/=�B=�0=�wG����U�9��Df<$M=N�˼�N���;[�M��Si�&�Y���></e�=�=��s�&�#=�i�;}sM=�e,���q���!����<�ۃ<�Q�B�j=��R=Pϼ���;2g��3�<�=z
���� =3�=[�*:=O6{�C�ݻX��;	#G=야��1 =}���D�m�ڙR=F��<���<O���R�P<�'�<�H��d, <�7X��t�<�9!�̪ż��<��!=ro=$ɼ��-=�q;����=1�<�^���9=�ħ9��?��!.��H=6f|=�&ȼ,l1�ub�;����}<b�L��}ü6�(��ź�%=�*��d���"T�;�!�<�B<�"ڼfY=/f��h�:��<�g;A2�<���?=o��;\�2=5&J=��;��R��j��-�O�)m�Xݼ<���;�<Tv%��^��P=�~f��%t�*����յ� p=q�<�6N= y���1<�,�i�<���<$����?7=���<���<\R=ϊ:=Uށ����AZ=O4���3M=�Dڼ{�P�L�Ӽ�ݼ���<���9aI�F5$��z���;��;�����<��r<�<a<f���Vk�<d��m7���2�����8�=�	=k��	�����;$�<�̼�3<��=-�'<�g����<]�=����
C�Z�}��n =.��0��i�=�y=А�9��=�K���<F�R���f=H�0=}��<Hm�<h��'�D����S�(&�;U�<3Q<E���3z�;��O< ��<�T=�3�m��5=� ���:�>}a�x2���F=N3)=��A=���;�A�}T=�	4=�$���.=�+j<�F4<�:=�rQ�!�=���)�o�>���b��<��B=yv���?�d�9�ln�q�}�7����<VzQ=ܵ<`h=�HX���&=��7]t=N9��V�<��<:{R�<̙,�Ù��u	�ѕ]=A��������l�;ׇ �/��<S|=٘=C��(9=n�����<Gȹ�&c��ua=��|<�32=g6��A��<�٤����<r7=?|���6�L��χs��{Ҽ�45��}ür�U�Z�>�@�9=2-@=I�{<&"[<HL=<��<����^�M<y��<��;q��<_a��%$��=�<��[=�U[�T���5����D=}��~=�=-6=:l�;̛�;qR�<h=c�\�8�K=�
=nc��m�;���;!tͼU�����Z;=j��v�y='W=Y��i�*�wp"�[�!<�i}=�T�<��O�Ȓ�����Q�W=q��ӵ#=��6=~�8;�z�;T�A<	;��EPf�E�D=`#1��G-;3�f��N�;1uk=��v�/^��Ē<�Z@�2��V>�s��<��Y�o1�<3d<�G�����8���7<R
=�Po=��<��ϼ�Zļ&�*=z�b�γ<�=}��<��D<��=J�Ȉ=��|=uwV��y�M�Kd�<H=J������^<k<�
�b�r錼�!�K���AQ=R\�Q�Qe=� ��m�����ռ���uǼ��N<�� ��6=�M����w#< �H=���e-=�rD=�N�������@=���J>�q��%h�v͚;��^�Õ����_<\�4���$=���n��<��"=���%7=��p=<����<��(���I�11�������ڼ��?�����9%=np/=��0=���&}4<HT�<��S�#=��/�~�<g7��{��D�8C�<��b���u��~D������\�<|^��VZ=�pb�3�<�3=,��/��;e!<�Sb=�r<��O��R���j=��=jO�=6O=A�໺-+=ZhH<���RO�[܏;��;�t�３zZ=��<�wV=E�{����<��2�kR<=74�+�M=}Ũ���<F�e���q=U[=���<��;�9e��9=&c'=�塼b���PO<�^n�Р�;�=��UT=Z����ә�-�U=�\�<�\S�5�=���;���j���kX�$:u<�M��q����s��8��2	S�ӌ"��LG=��<q���!=N|=?�=��=(?6��=4����pT�7F���=N��<
�Լ[j���lP;H���1;�yT=�
=Q����K:;V�h=M�5�q:��@==��<�#�<-D���Vu<\�d=,d<�����R=k;��$�<w��<��,=n`S=�6=w�e<���g޼ZD���%�˯ѼK�D�0^n�Ԏ��e���I��S�=Z�TCw�g�l�+��ł�6�<�<Ӂ�=ҫ3���<�b�����o�Ⱥg��N_h=��<d�l=�P_���+���/��«<��;<�%��q��ad<�"a=��O��?S=c\l;�)��0t���Ѽ=v=/�Z�xi����<g>]=��<!�����ѩ���2���]���{P<�7�;93�:I�N����<��ɺy�Q=�iT�� <9G�g�e�� -���E=!�a�b�H;�-�&;Y�<ź1=>��������;d<�<=8�<�Ѓ<��Z�!m�<�y<=8=��߻e7_�X�.=y=����*�<��>=|h=* =*�����r���e;�F<e���2�<0}G�h�=)�9=㘫�m�"<$�k=a�;��g]=����=����}��ݜ}�
G����l�~���<��L����c-O=)����o�I\�	I[�lob���<���,�F=}^;O<��A�y���ֆu���?�4!_�Q=F솼`��'F��u<���R��;�=��@=M�[��6�/��a�$���ӧ�<�=T`�<�H�<R�"<��W=�����ӯ<�1u=�]=�/�d�w=Ę1=W)Q�Ȧû��"=�\����;�[޺_�q=[a�Z�:[+&���N���K������Vݒ<�3_�-�"="�H=�Y;R��<0�=�5��7���Y�D�Y>�<'v�<b����gɼ��<=�<��;<'z;P�=!&�<� m=���<s��x\�<r���v˞<5�U�$�<�b�<_����]=─���&;�W=P&=[-"=�k�<`75=��żQ|T���)=���0A���<��<ґ<O�=�s��Zq����Ƽ{H<0ڀ�/�¼���4�X=V�4��CM=��;j`�<���H�?=>&G=��;�J4=�6<�j�=�Ci�5< ��<�<V��ʝX=N���f�+����4�$ǥ��?Ӽ�Y�^��<�Z,�Ƞ+��q���=&�4�� ��/ļ@�4悽���Du2�nz=jj@=�;�<�K���:�o�:Ū<�*v<%"�<�T��h�=��5�u@��v�=�&:��$�'$*=��G=ߟc<�q�<'�=�F�<X==���ք<��|�����&�<9h;O�W�9�o��IN=��V=k���[��QL�;��;N�=¢c<S��<�?�<�I�<�8��i6�t2�;i�<��<��<�3=�6˼D:�;��R���O=���:�{'=xW��`Ἅ�6=P\����dy�<�1m�W'�,�������H4�<	��"���p_���;6ü�g�={��<�`�;�C��j�+�P�O<�5+����S�<�`ϺӃ=̙���|�<��O���_=���/=��<B�=]܂�3��;p�{=
����c��~<=.p���B�˾�<ih=�a2��23��K=:�d�\�����-ޑ<4�ռe>�I��_�?��_��p�<�Г<M-=U�<�|0= �=�T�<<�T�����g��������OԲ��ռ�e;��N�����<�}��t<�)�<�0�<XA�<�Og=EG=2RO=�5�Ln�߭�G=Sl*�#���>=��[<;��<\� ��l��˺���;����ջ�L=�u�<R�����9R�鼿Q��<8��B�����6��=�G��A������Ğ=_��<���kH6=a�x����(��<2��<x�����I<��3=�+�<9I*=�~�JAp</�����Q�@��AW=�V�:��}�.8�:�=~���/�F<��V���<ݻn�=@��;����s)=�!=W+#<�P=N���b��WS=M%�VW:=殌��x =?D=�c����=�#9=zzB=���9y�<�m=��n<N�;B[���;u��)���߼�XB�3V��Z�L�C�
�iv����+=�A����d� G^�yI����"=���<��=#]X=\��<ST@���W�i�=��7=�&��L=
�w�f�B�����BwU=�+��(k;�C*���=ŵ"���C��:�<��=���o<�;\=�B[�د<���< �=;�R<�O=	�<��¼���<@l=���F����L��z��ڋ�<�0R��0�<߫�s�	����<�rV:I�'=8�=��<�=���oY:p�����G.7=-��:�<'9�(�=B���N=��=�?=�t[˼��;=6Y�<)u1������2<�	<2黱jO��e=�ݼ��
�5�< �����<R�s�'Dǻ.�	���=Lr�+�<�`)�s�<npE��(;Fg=c@a�[��� ���g=	ə<x0ۼc��#�W=��<���;���`3�cR�<}��<��<��s�
����<�p?<�h��盻g|�<<�eX�|1|�-D^=�IH=��F=�3\=��^����;+���Ƃ�=��>=����r�˻}�=X,�< ��hĬ�y�=9�q���F=�'�۾T<���҂�`̯����<�kۻ��
=W�6=�84�h=�b0=�1���܂<���3,��d�<Ő�<"��<MS��*3 �W�j=�9��]0=�<f�7N7=��q�.�<`���VF��J�h����A����fc������$�=�E�e<��-=���.$��t$�hi��.8�#�����r��=u�9=�W�<�;�<ؽ�$K=�Iغ���<H�>=M4(<Z[�;Ju�j�3�KV�cv�n=�<�s�7�;p���� һn&��, �h$�</-p=��=�&Q�X1x<��<
�=`U,�Ү��:f<��M���h;��<��h�L���=Am =���� ��X�<���;3�N=�S'��Ʉ;W�W<O��<�1�<:E�<P��=���M�x���t�;%Q;m�<���<��m��Q
��jK�a�l�sV=OB��Y=kO��Uvc����jh�_|\=��\�u�n��_�����<nL=�3H=Ќ��q��{�;�i�=N>j<+��<c�D�A&#���<�p�	��<-�D;[0=�1� 
��;X=�=��f�~Xa�����ռE1�����/����<��!=&g��]�<��<��]��� ��=g�a��3%�.BF;�3����=�b���`�$\(��T�:��^=��?<�����	�r��w:b=�9�;Q�ɥC=l��J��<�~��i==8o=��� <!�r<���<�G0=�#�����+�<_ʼL'S;�m��:���0�Խ=��B����H�@=gN��=���<�
#<&��<��\�����H;dXͼW�<]�p)�;4в��==A�ݻʻ�#���%���C=5s<	��:��ӌ3���A�G������<m�-���(��D�:��=�l`��w.=�#��Q`=�A���<>.���)�<����1=<S=�c=��S=#�p<�_ =f~��S�D�/ ���UC=�h�\;H=��x�=�ͼ�1<?�<�Z ���
�*���4�3�5=�7g<:5ּ'����0����<ߠh�~���h)G�y�<� �
yּ[)=��;ƅ���i;;/����j=��j<�{/=��a=,v=r�<���=C�9��?��\��]]=�dH�բ<aW=��Z<��`<.��^k�<$�<���<��<��H;=�0�"w|<���a6=gT�<�R=�x�����<��p< �;k=�<#�û�23��n�"�=�mF�q�F�$�A������) �[�;�<���<�/1=uXH=<�*���<`��=��:����=�6�<�`5=4֬<0�;�-��;c�#��{���<�o/���&=J�ۼYc^=ֽ�<�!�<U�9��p�;=������ż��漻c��@O�ق<%�=d�%��S<����x�`��4����'9=���j��5�<�����=1<�Z�<ж<Y�^;pt��ӿm=�U�:�)y������{ż��<H*��!�<��j<.��Ҥ<��������=��e=Vq�<�k=}>B�p�4��v��#:s��_]��}=a�!=��|c�<8�d����;��T��哼ް�< I�������Y=���=�M<�4L=֏��-k¼=X�;�)h��%r<.%h��Xf<�]� ���6���,,=z�	�'�~Ѕ��@�q*�<�z*=�-�у�<z��<f�߼�5�b���\=
���QQ��']=�<�^Z�;�� uV<��E�</R���n=w;����<#��<���<1�'��u=Fߞ<G��<��Լhm���,�<2��eW���D�ʼ�����hu���B=f��4ͬ�F�.�$/ʼ�87<Jh�<��k���Q��,=O]*��2~������=�6��߼z�;=�WR<��c��n����;zs=��ּ��u�5k���#�<í�EFn��렼��Tn�<Z���-��Y=4�����6=��4�W|<Y����� *[=Xʃ��g=Kc����7=5����==0���L=��<q��<�Lȼ�`@='*=�g�<��=�R'� "=�Q�œ<�<�m=�Ǳ��Ж;M�*=f�@=`"�5��Q� ��ɣ<?1=�燿�P�<��+��Y�+�'=,�<v������P���ؼ-=f��<(2��\1=Bv=*��;�H����C=��==��<�s�<m�AѼ�=i���"=g�(�m��<h��C���b���<M�<�Y�$w;�b��e�/����/�I=S�	����<?ږ��l� ����q�U�<`✼P�B=X���(#=|�»c��<^3$�PA���q0���<��X�ی�<�K�<�)4<�+o�'��<l9һ��f�IB�C/z=��=%�6=6�;�ׄ���
AJ=0?�<�<�<��A;Ͻj=�+'�'�o=d��s5=\��<�̔��3j��H=3I@<[L��<�v=�@�BN�<��#=�N'�����+=
����L�:L�Z�������R�GB��떼�'8��Br=��M<��-=��&=m���ˤ�<�׋<�8z:��X;.W��m�<o�����,n�����H��{0�<F=2�pP=�T��h�<6��;!<N|M���'��y9
/���.�<� ��=5X�<�@�<� �[����f�a�5=��<w�:=$�ʼ��g��ؼt���d���=|�,��>=�?+=.�<gg
=!�:��=(�ԼX%��A=��&�wؚ:.T�;�� 	����ۻ�N|=4b<�����s<��0=b�<�2=�a������d��E+�a�%�o%=Lr�)*2����<W;ʼx�K��ܒ�=�}=I$<b����%�����ְ�;$ø<�.�<v=j�9�)�Ǽ�>=��#=W������<C}p<K�r=�7+������u=�.��J��<\|-=��=�y�;�����]<��)��C����;!=�k�K��<�As�0w��mC<e=9������[=��!��k =a�=o�.<��H=��S<₱��Kw��za:�n���������:9I=r��<z+��z:�~ ;�AQ=s��=E+�����<�l�<��ĎK�"u.���9R�wEp�B�YIM��z��g=!3=��6�{=�U��0�<�C�<5�Ἃ����Kټ��z=ک=R�8��� �����=�_�<v�����V�+=Q"�O��<�ω<�e'=�
�<ӣ<4���0x�����d=��+j<$̼+��M=J�<%Br�!CR���W�&n��FGX��3<Ts8�M/=�o�������Y%��C�:%_=�q<�<#���<ί8��A����k�Qj)���:�"&=-|��X������.=%�K=���f5Q=�"���B�1=��=��4�AA��
~=䗵;��/��'�c:=�%ټy s<�V<*$�r�����<$4�k�_���ϼȆZ=�?��mڱ<��i=��o��-:=O�=��D�`ŕ��=lk]<����R��.��p��*1<7�����=�u=vX��މ=<0�<�ʆ����<#e=� =�B�b�"�b� �G���q�U�N�E����!�=�8��s���"�4��:�;ܣ�<z�|�4��HB=�����<;�2=(AH="��;�׮�!�h<�$2��R���=Tt�$J��$W=ɇ=�g���j(�; t��q��r9�<�	�<�X���US�ZH�<k�'=�[=�0���$ɼ��=��k=O�=B�����̼�J(<�t@�a㼩�>�*~0;0&���n=pD<�KR=+�e�����Hg�/��<�'��<$���ɩ=� <=�N< ��0=۬4=�Ap;���<�P=�]���Y<���<�4<W9=Ε[=2����e<0缚�R<��C�S
��^sL=�ݢ<!�]<����\����;9���G�-��N<�λ}�X�7=@`��<;�f�{�ֈ��̉B��F���,='�J���<D��M�F=���@�i����<�/켠���R<�_Q=���<��I=�Z���3=xB�~~���z�<�E	=V@N=«�;�&4=6�[<��޼���;~�*��q<l�3�����v/��g���=�p=CB�:Q�L�n�;�=�����*D��ˁ<C�X=_.|<걺~=(.I��ѩ<���,3i�-���nM��������;7-�J����-�D�w��J�;y}^=wH�<�]<n �a���3<����=_:t�-�<�'Y;}��|3<y4:Be0��X��~�6��BѼ�	M=�b`;]�8=��:�<a�&�B�S&O��?��wJ�<�b��pa#<�s�<	�=ÚD=�����*=;�4��=��l�=g�e=��d=OO/=���<��<� [=�y��V<��Q<w��<TO%=���=>��2=bw�6��<qd�<��:<T����<1��;!��A $��GD��=wx�<��:=�`H��m==|�<�۶< o�g���݋#=�F�<�ݾ��z��U��G�����<��;�0U=��<��1M�<`z�<9o���J=�&�ލ���z�q8q��׬��k�
-O=�2><Op�������<��� K��~޼<$�ǼÄ��E�b�m���A3=�7̼d1=��=<\}b�U-=�)���dx=a��<�uM<-�;8��&�<�)=��ּrs������i=x�<�&)=z!�y�~��Y�<4l�<b��T�=<���1�¼bD�W��KE.<�@>=K�|����\F��=uE��3=P4V����<�=]&<����������-��	y���<��"=(��������\=v�?<)��<��<��<n�1;�^{<�]̼2g��z�6���=�j�<�c2;̌Y<x�<���iW��d:=~�;�*,��3=�a=��+�u�"=������<���<5Rp=�NP;i��<_۫�[���=���<,S�S=�}�hs�;F�����<q��I�p;(�<��伎�����<H�3�2=�7��/�?:�<�D?�C�?�u�)=�'ܼ6�M=C=���t��<c��]v=9?׻�W��iU=��Y� ֞;�<Z��;RU����p�_�����=$x�;3��<VT�<��Q=d��"��<��0��;��=�����<����|�4=5�<M�h=ZT�<z�6<ʷd��&=<I	^�wtb������(<�o!<���;�r���L�悛���]���������\7=šF:��<v�a��@���IC��!�;��:=��=_�����%= �;����^=�&<e&L=WyP=����hT�M8]��AZ���t;�B���˼�87�����<P��7�U=3�;hcV:5��:�6���=�_μ"="=�A�2��Ƽ�Yq�e��P{-�Yn%=�"�:[u�=�ڜ<�;[�;�@���\=x�F6�=�=e�'��:=�?"=�)�����
"�;?;=�r���M���<S�U=Z�<�@=�J��ma��\=`��=��=y��<��N�Z�-=��B�Z����Y��r:��.(=��U<_ �H�1��/��yPa�y�F�d</Zz�k��<8'�<�IQ<>ļ�^;<�ϰ��ݍ��Z=�+��;fY��=�~8=�>=�l����:�O�Ƽ�����w���<,��`�=oc�">��8=�ci��/�;�T_�qBB<�!<�U�f��<��"�;=QgP��b���	f����y����6<^�H;�6܀�����͞���=w�"=�~�;�Z� ��;M�	����r�� =����<�f�� 2=��?�^?�<��-��Iv��0v<4�=R�弘�����;5�7�*m(=��m�}X�<d�<�7=<����j<�a��[<=�AR�p2=TP�P�#=KN��_ <dK�펀=q=���=��I������Y�<���<�;�Z�Ǽ�=����:��=��=�)�<�[�<�>=۽���`F<��@<�Ȼ��e���x<�2V=4���%)=aPͼG�_=��+�Ye�Zͩ<'��:�0#<M��<�߼:�����<��*=��Z��L���=��=w�����60=��@ =�U�<�<u=�st<���<�b�<}X�<~�P���}T=)7��
I=��<�~�1�<���<���<���<����o�:���<T��<��;���<R�<��@�󯷼'[��.<�x;=<%�;4zW�HG ��2�",=��N�|�/�Nz�<L%�;��*=��\�j��<���+{=�LX=��<`��<�+�==	�"�W�Y�����.���@��wX<Vt�<@<��ﳂ=v[���)	�?%2<��s������O��E>+���=�9�z0���(=���:�E*=^=� =GSd=�+4�mK�<������<<(=������G�P�$�z;�ϼF�S�4�A=y��/T}��mz��X��p =��Y�/=�.�<�e@=~�:;��`�l=A�D=і=��UļE	�;ei�<�=^����Y�<��7=JǼpp=���_=�<�N�o�����	;Xu��u'��e<�MR�c5=�ҙ<ķJ����H�.��K:���������F���O����D��9�r�t����J5���=L��<�x�=U���q6�W~;�ܼ�� ;���nO����4����<k("<K�= %^=�V��-=�M��*��<5q��Kk�$�!_I�t�<�+j=�F�<�E���-=u;�7�׼�s;7�� v]�Z #��A�/x�=6�-�k�%��Q�;���<8y�<���<�,<���;`f�mĹ<ϋ!=2]U��<��&�?b=�F
�����r2:%���k���H�<p�g���-�L/
�Ւ�:�>g<*X�;/�Ҽ���8<R=�B==�<�d=�)�;n��'	��;��<!=��%�]��뙼��'==t=eQ"=#�x=�:i=4�O=���� 	�C�ɺ��	<up�<���<uջ�U|=�v��ˌ�R!̼x���5�<X�!�+��<g=Δ@���\�)���9�<z�F=��U<3�)�����<oݨ<UI�<��2�$�/=
8��Ĵ�L+Z;*��<��<��6��L�'l7�i搼���<�D+=�J��UE<�@����wϼX���cV=Uol=�)�<�e��GIR=��eI���,��'��<Yzv��9F��񹻂0-�m9=7_��uX<S�=�5ϻ�&�<��?��@l=��R��X4=�p�<�86���<-˿��a"=j�U���>��Vp�6��D��<� <6.=)�&8;����M�p<��-�'[1�=�c��䄘<m�B�����
;=��:�}J�K���;B�<�mr=�4R=]�}���Q=h3<���<Gp;<�Zj<��8��%�<�#��v<��;�'<g�<f�|�m��<��8��V�������Sm��[<���<��7�&���9��o�;-�|�ZѤ���^=Mr^�L���N��?n)��/�<�H=��*��3�	m;h�8^��2�=��M�;=Z�E=c�<�bw���v��� �);0�=8=��#���]=�=����5Z'=x�<Z31=�
==4
<k�f�q���{��rK<�\�</���E�u<�I=�j�<���<R��=lD���D=Vi�����<z�ݼ5�"���B3�̃�<���;��ػ��7�wW�<�f����.�� N=��=mF=�k�<�]A�O_���
�H\%=d�P=[���Ϫ�<B_�����pT�������:��Y<�r�<�0�<e� �9̼f�;sd"�����x�<�&'��缰��<4^��M0�~�R�H?M�8�`:,�L=M��D��2����= ��<$���"<Ny�w0�������<kM=n)��l�;��¼ �b�����K=qL%= �E<�J=fS��sG������2�{0����̼��F�ٞB���E��0���(=������<�5��{wP=���<�5+�a@8��ì���0=d��<�9h=�rH=��7�����o�<��<'3���-=�5�;�������qL=��]<��=�b.�tΙ��3�4����`�z��<ݹz���^�AԼ��ѻ���=����1��Q�q/�U1=+-<xn�y��;:�d�L<J�<��91A<�yƼu�9.�� �<V=�<�$��ݗ�kO.=6q?=��%< �;= '(=)�=�z�<n5��]<���t�<a!��*p���?P�D��<D���3�=�mL=�+3=r[=��<Q1�<�.��܁�B*��ZR<��V�I��������DJ��(���a=Z�:w���d7�<�C��K��&Z=�s?;���>�Ќ��O+�4C����9^8>=�b�M��;���T��)�#�8�2ϝ<a�=�e�;#��<ά�<_$ֻ��[�d�<��L��<f�<*�<�O���F<��=��)=I�A���X=��!=&��l���32���b=.��<�z�<3��<��l<	�^��7`��Խ<_��;�w�sT;=�9����7͓:�T<����<�u���R=��;o�=��<�	�Y�=�UF=ؾ��0x!=�8������<ږB<�v뼇_� �d�j�p<���R����#[=��.<�#=���<ӗ<��D=i�u<�Q�p>4<�T�;��&=�h�<�c���>@���9e,�0.;��j���)/�ztؼA�f=8#�</:�?�5�D=��=$��$�x=��R�Ne���S=|Rw��ۼHA9=�U"�^��<��<���<P�=f3g�M*(��K��!��<��Z�i��;]�<��;r�F�����$=�S{<��e��zM���(=I+=e2�<#A=�˻�jL=���<tD��N)=���M�<�7@��-i=kI]=B=;�/B;�!��ۧ�<��;-R��s�}�b��WR�`�;=<e=��h;�����8��=�<aSü.u�<2= ��;3߮;n�w;�[�<rUt=�<�<�[]�SGW=�����#<i��<�v=]\��O�<�v�<_v�;�D����Q�=�<	��x�={N¼-N��E1=��x=��ü+t���F�mˉ<��p=��ߖk=A�=�M���=M�x<��;��6}�Y�6��a��"=��=&K=�̖����<�?�$) =;1�&��<�%<5qb���a<x3����$��;��=�I�<.+=�Ƽ�r���u4�%M�<�\��(Tb<�8�Q�9=�#�<Dx"=�x<����kG����9G�M=��A�8u[=�Ź<��=�^�<&�= B=� ���=j@=�3/=������}3=��<9��w<�< ��<��<��==��R=o��^O��<$��Za��!�<E�к3���FE=����DMd=&^�<-$=W�`<���<.R�9�����C�&.f��_�im4=��<��N<��<��<m+�<���< ��<~��"�r<mVf<k�뼬��<�[���=��Ǽ�5��l?=�g;���<(��z�&=�GӼ�%?�Z���?/��2�  E���N=��a�v�G���<)�	=�5��es=�jy<��<���<R�=0�C�'�Z=e����f��{�<6�Ѻ�K"=g#O���2O==��я��w#=j���T��f��<�k����}!I=c>�z�p=a=g����tz=�V�;�S=,œ<��";��_�}������>v=A��ɺA]�<^N	=!W�|A�;_Ý��!r���)<&)�<ز=�$��+�����R�E=����4<�F�?= *���G�;��B=��6=G���#�=G/<3=��p�Iu5�ܶ�<Lyc=�i����֭�<7�T=$6y;(�<N�L����)Qr����<	4ҹ��,7m�v����;�/�=I=��.�Tм=L�Y�@=	=�;��7��=�S�<��C��s3���Ẉi�<��&;�7���^=1�ڹ>ܣ�����j�r�M���F=S�:�)����5ȕ�S�M=�=�>�<�CK�]�;X��<J�d�J<�[+���<b����;t1=c	=3�p=���)f=�f�<F&~�n�F��X�-��<(�.=�����=E�=�=/���&�ʊż���;��<8BK=9ܼ��M=��<Ճ<�M���S�D�@�CW�i�t<%�<hx�mW=�'�= ��M��7a��^=��C=�!^��$o<z <;�Yˎ���7��1μ(�X��O�<�R=��3=��i���F=��<@�5���;��3�L%�d�3=I�����<��S:/0=G27�����z2�@�;��<�v`��;=�z��`�=�����M3�G3r�\h�����-\:������=��=��<�d=!Ad=����&�R�e<� 	=���;i�7���f<V�����O?=eB=Hx4<��4�����}	��B=1[�<]��<�����V;�c"=��O;X.�<��� a<Ǩ���:��Cש<�`���l��]�)=��F<m��<7��=z�;׃0��-'<��K=�=>3j<�9	�I�(�;V9>=J=��<8�U=a:F��,J��m<���S�ּ�|�����7�����<��#���j�7��<-�����<O����楼#�,�������g�<в��c���R�<����3�;])E=�O�b��<��=�}t���;L=q^;�`;��ϻ-ٷ�
+��M�<��Y;��y<Q���e��<�ռ=�/�^/�b�<P���4=��$���F�9x�<�b߼8�<7<�*$=g�!�Z=� ���,��Z�C4<D�=GY=ק&=�=�ɻG�=:�<H �;"�5�vVR�|Z�<5S�<z��<~b�Yo �9��X�ͼ�%M���X�ػ���<�ܽ;��m< ��<;��={�<L�==�jY=�E���7=O�X=�S=���<����1=�P�<t�-��1��$^=~�.�4���*��t��t伩�l�j�A�� ^�2n�<92t�/Z=�L�m�V�L;�E��<@�l�H��<��A����<��<���LU=<����A�4���$�
h�<`w~�({f�S��!�;�Z�;��;�W���uQ���<��D=�p�;	���F@�<�&�<A[=q�!�a�z=��D=-k=֑=�w\��J=־-���.��<+�����;#:�ѥ(=u2)�̎��e�D;�(O<���m��XfT�#���I<���}*�<YP��+�f�~�� =r<�6���P��e� �ö��������;�j�<�Ju;L�@�cb����D=)��<*����#=6gZ=� ݼ�,=oa=��<��i_�O�ۼ˺9�����˼��N�E|�<r�=��C=Q�Ə&= #�<�Y=�˼�h=k�g<Չ=;T=��@=���2a�y��<L]���0�I��E�K��<8
�<�=�aM=~T�%V�<s\-�>�<=���<%8=��B=иռ}٢�5�M<cVT<��=G�<� ����z=:;�[	�(�=;I�<�ľ��Oջw��<}�̼�Aa<��	���w��<z���~��=`]=x�=�o����<|���˂� �N<��G=�1�� <�w� 	k=��<�2̼����x��ԝ�<��;
��;��H�r�-<��<}1F=�̘��M=����?=�ؼ��<�� =�5=	i��2�߼�jk�-��<!(8��L������tA�/��=a�!�U.Q=x��A�:��t�$"f��s���ü @F����=�+���<@�<�rK;��I���<E�=�(=�;�tw=��=`E`=]��=Ԋu�l��;#ׇ<�D'==�>;I�=�.2=�~��h�������8��'2=�`4=�$=�:)= C(=#͆;���<`B*=UY=XE=���<��*=뻞<(2�Oe9��< ��x�<}�s=ɾ�<��S=�W��w��<�q޻����u<+��:B�{��G<���<��i�9����C<�=�C`=�W�ь����I=rշ<���<N��<��*�;l��<�3�7+���{�s]h�%v��ME��}����J�X���5�=F�C�o��<|��ީ;���<0�<�=��I��<l��kl���6��@<,H;]G�4[��5�;���<Ά�;a@7�D���?��l;y�B�'�#����<�V�<.�B<<��<d��CCm=�֓������ܼ�G��{<%$�<���ƒ=�����@b��0�� 0����<*=�<� �d�(��i= ���=���f%=�>���=Q�/�_��=�������e=AG��3���<ܼ�?��7��ɗ�;����픻A.e�ij�;4���4G��2�Ɇc<JhH=cH�:�= �=��L<L@=Do������c�9��<��]��"=!sڼ�M@=�J=��#�1�ݼl����=�=F�=�=�<�!)��O�<��	=~�߻�5={���s��R=�J�<X=��.�go޻�_��{,�xc��f�;n�&��k=1�=�R��r=&�W�M�C=O+6��?�V�+=bs�<���<�{=�lH�F�<�{����<�)c���<�A�<f�K<\��l�`=�!�;1�2�Z�<�E�<A��<�S=� ��L�NL=*�"=&J�>^o���Ƽ)Eü%<f;�a���<�W���G==;H=�JD�,^g������%���+��3�=",��M`[<��9=3a��0���r��q��<K�<Ht�<|�_=��U<i3=��;s�O=߸Z�@	%<'���TE�<G�=����	9���&�<�]��_�z���V=�:����oڛ�m��<��<:�Y�8� =��o�i�x���c�b�<�l�:z%����Z��8+&�l"<OG�-����i�G�[<7�<��q��&������+��m��;�A ��?���u<�����,�a�<�zм2�ؼ ő=ۼ�<e1<Q��;�L":w1�l���;�<��<$0P=�`��*�E�U��B��!4=c�@=BF�<�"=�NQ=��U���Y= ,6<Ns �Y?=��\<]ڼ�=�$���n�<�rg�}]�Ձ�<eِ�J3=��b��� <�^=ZS�<ղ�:f�<'FM<�c'�;^=��7=�a=ls����<�6=�IA���]�ļ�h<��8���J�j�@�mM	�z=��
=<�=�22=q���S�-�8���K��;�"�<� =W2=ǖL�}J6<�f#<)��Y��a��<���<¸R��*e���&;~�C=�.�<0�7=�(�O߼</^�_ϓ��苺��T�u���k=8�;G2T=�K	�ň�����K�gX����<k	2�A?����'��[=���;
d�<~Sm�K��;�0�<ٷM=��4=)�5�;Iqk=�=�	M=3�<[﫼��>��q<�Iu<\ؓ<�G=G�;D1��} V��ID=�h����=J�Y��0M��遽=o�;��d=�s�:6]e�C�L��=�<R��[�<��=�rn=#a=y7��F)<W�=-^�<�=���1@����м��H=��i��U>��t=v�%=#�vMh=Z�?�}��ַi=�J�����<��Y�Qq�������[��=�dؼ~0="���T<IƁ=�ZW<d��<<�~<��9<��g<�<R(<��q;
�*�=�*
=�ד��L<�2�<�x=��:��L<�zx=����0=�yF���s�<�	�J�B�Z��<.�*=�=i.��������� �W�[���=wZ<�@�:�b���ȼ����j���2��.���v3�T��4(�<�u�<��'�ܫ����<;��<ԇ�<��I�yKѺ���6R��'��M=�`Y��E���u7���N���>=K�d=R7<K�(=W��<H���)O=<y���==o�<�.x���=�h{��G=,������9���<��J=Lr\�$�$�¿�<ʱ�=C�@��¼'�V=N�<A����b�=yw�W�=�-8����<�~��t���-������K�#�m�l�H����=t����<^�<g�o�l&v<u��t=����ٓ�=7Y��Si�t���H<��E���4�f`���@:RQ�'sX�+�l=��g��?�/'��P�(�3=-�ɼ ��<t.�<�<í=L(=,���n=L�	=�=�uH����<)D��W=�������<��A����$r<���f;��~I��P=�߫; v�s��<Èn;��C=��Ǽ82޻��<,�<��4�,����$;�)�I��q���컫���{�;�} =�~�<�\��ש:�w<!�<og����=ܧQ=oo꼷A<��8<��`=5Ǝ��mj��Af�nO
�C����X���O������"��7�js��I��Ł&=��v���=�y1���c�.D~=7��<9~;={vϼ�E4�{�=�
�;��0�q�Ѽ���<����e�<��y�s��=N�T�|IC=N�M��)���aļ��	�#�R��G��7���}��U��O=gAk�!H=���k���%=�S]<�����<D=�$�<`�)��;����B�R��$�<*���ָN��-?�<�k��D�=�#�h�n=��V=��N=a�<�犼g��<'�+=��}=�x�;�u�;��W���<�R���m��΂�ס<^��<�l=�)�;fN�<q�<�{�>�7�-%B�t I=;_�}�k<�BH�_C�p�+=�E=�	+=�p	=�.7= 4/<�"��,�<䳰<.�	���<�9ۼ2d��#P� ='��<�a_��[�<�VC9G��;)<n<��
=[=e�.=�-<?f�]��^J�6-�hP�<5��<�B/�����K��	�f��g�<H�T�V�s`=�?����%�K�h=7���҈<�����p�����[������L=�O�<c�=�F���{�E�;�_X=oa�:�r��N_'=�.廏�򻝉^<��N;�>��'=�WG=O?�\�/����<�w̼�9=�ë��9,����0,=ep�<��;ߕU=���;��o=�冻��P�٠N=S�E=�6����v҂<���Y~j<�.s<�6ͺ9�"�:�=HPżF=������<�$߻;��<��K�
y=�>��K��'�	�_�=3Z���<?&�2��<f�;�䬼��.��V����<xbh��ii=�G��n;����v��yQ=��%<��;m(���P<�`�<��V��<�W:���c������=�3=���:C="��D���.=��$<k�=�zHe=w�_�׼@H<o[��w=x��<�J6�����<����1s3����<gv�=V����O=��&=�z���ļ��=�Y���L;�=����='��;v��:��\��Lf=��<��r=1쎽4�F=�!�<�*Y<�	�=�hT=����n�3�&��<O:��^��(r�:�ng�i�4���<�=��}��h�!��<\lʹ��7=5��:;=��*=��K=���<�YP=ؘ�<��j<���)N��*/�쏤<��QB<T�?õ<�����=
B���ӆ<L�̼�����MD=M��<�#6�cΡ��~(��)�[J[=���;�9W�"�@��S����;.?�;�C㻀�o<0��	`N=��W���=U9�<V+���=H��<X[��o�H<m�N=^�Z�<i(=�d�<�H�0MO�$Κ�C��<NՋ���=��޼c�=����M='��<:���1��f^!=�'l���w<�_+�z���y�����)����q;�Ƽ1�a�x�<��������y<��<G��<�0X�������o;�G�;��;X<�<RR=�X:��SI��+�;�����j�>Z�;y�O=v(�<�&�<�A:/�=�>5�C�'����57h�a�h,=a0=��7=�I'<��K�/h�c=Z!��[9���t=-��<�o<��4� W�<͙��=��:��!��&=s?����<�1\=ma =
cI=(��؀*=he<�਼B?=I�q;ɭ�<���YR;�����t=�N�]�<��b�e/;=AD�<�	"=Er��ia�I�.=��ϼ��<������<��=��q)=�� � �N=���<:�L=���<8��;�$F=�U�*� =�̙<Q�r=7c�<R�<S"=q�.=�|=���<��_�P�N�<=�����9<�2�<7\9��Z�<L#'=��a=R� �1�;wꦼ�����B=�!<:��7�:n=��<4�5=i+�<"\=�v�<��1=�Pf������N�_蒽�G��7b =�g#�h�=�+��m���?�^�:����?=�`���]<�Ф<��
�1sڼ��f=�j��vW<� �=�v�<\�=��м"�޼v����s���=3q�<Yh��r��<��=���;f���.o=����_�R���=���<t��V�j;v�K=����t|Q=wmR�ֹ8�{��;��)=�\o�%�<m��<���<�����q�n�<�0ϼ ~����r�g���T9�5�"��-�<V������-0�Z���k���ǼEE�<u�J#�C�=��?��4ʺ��y=-�Ƽ]�����8�-�H=j=*rK=��"=�q;I�d�# ���%=���<����U�<�=�=0=��h�?�<��<��7<kU�*p�<<=,�q<�����m&;��^=A.=&���M���<;NB<�p=�*3�
Z=vC�;�A��Ng=Z,w;S�%<�_�4=�4���@�\��}��Pr_���E<�c=2�<�JK<�<@�ςK�:�:Ǒ	<��=�O3�<�l/=c�:��޼
���_�ܜ-�X�_�����<ѵt=sB8=�5<���;�ֈ<.Ѽq{��$�<��
������q=�o<�o��=��=��Xy=�X=�}=�{I�b�=��=�X���+=����p~�w��;\TG<�B��G��+�9eV��}r�&�<�B�<"��<}C=�m�<�^^=2/=����<h`�U�=�ʌ�1�=��Q=��#=Y'�<���\�=�::��6<�;���m=e���,=?�#�GY0�CB;�aR��8f���¸W�<�B;�i�=B���<ϼs�P=��=.�f<l�7=�4<Sv���ƃ�ݰ:���<u�C=��<P���{�; �ݫH��t��W��a|	�:^��ʯ<Ƞ˼(�4�������'�$=e�<>"�PP��+Ѽ/VK<�qS��BW�$�R=}>�<IT�v��;���<��=��c� *O=��G��/ <�?q�G\3��|C�)C��[��ė =�O<3��:*�o=��y<u��dB���/�,�Q�k��Aݼ�렻���բB=H��ߪX=w	����M��<<�X=�¼�oI=L��<#�-=A %�#e=i(;G8=�i4�Kz7�s�;�yQ�� F=Yn�Sg�;wut;�L���ջ#a<	k5����;RY\=W}<�p�n�/:X=�8��1��G1<���<����>=�3޼z5.=O�<�%p���E<��A<�`�S}���4=���;��T�m�#��<�<XK=9�����T5&��=A:ݼΏg�?�<�UQ9
�8=b�Ѻ�%=.?5<O���&�����<�����=�;��5�c;*i�:����2�D����ͼ,ڪ<?H��{��]���R�mn3=.��<��4=8:�:�`W<�[W���ڼ��̻�u�<v�����g<j
�nG�|T��,_;�m���"��$p�~K5�����t'�$!�;���;V���!�����$�<d4��1���<�_�ъ=ev�<^������	q0�3�<��!=�*R=9B<��7;��T��<��<����Nj�<l*������m����b=��e���<?0=�u�����zS�<�!S=��U����B����_<ݔ�F��<SH�;+;�% *�͠I���n��aһ5伳��t���Y=��s���<A�f;I�+����=wv=g3�d�}=t��<��=�n{<����+F���u��K��"'�����h�<�S=_+f=`Y+=��2�t��dI�,��TC=��M�u��g�U;x�9=��<��:<�z�<Ӽ=��)��=���<EV=��=��<�>A=A���^�<���F�Ƽ�f�dU7�N�@=9�
=�<��<[�U<�-Y�Ĺ\����Ȧ����<�-��Z(�f{�<�}-=h��i���)�;�5 ���@=2��N������S�O1����<t� ��]=�D=1��<�
�; `�p�<E��<�_^��x�<NF<]��c�V=o3<��&=�C��Fi�/�2 Z=�H�;�YS=<�(��h�<,��b���O���d�B��<��0��/�<6�^=��'=�2=��k<���;��t���L=U�<|~Ӽd��j����CXF�~��;��<�&\=$�=q�-=evԻ:6�<�����'6<�=
�&=��H��z�<���m9;�f(�_��wV=�c8�յ`<�{�;ZO=t�C���;����+=n#=�F���<��H<��<���=��<[a=z��<6��������D=�GQ=��<��%�cG=�>����;\��-=�$G<bF���a4=�}F=;�ܼە��1���һq�'<�S<�:1=W+�=��$=�hR:�)6����ɍ"=h����3�H�?�D<-$���{<�O�Tx�<��h��+=��%=��<�W<l�%�TJ׼�<���c<�Z=�B�<��F=��=2|<=|:�<�?���� �>ԉ<����P��<>��������v<+��bh��L2���=��;�0�<k��<�8�<�24�K�)<�����G:=L5)=��g��-=��#��Ņ<2�<��A#�zT=M�=��0��e�:���=L�J=S+�<;V������]�@��el�n�0���D )�.%��Zk=�;�Q=��g=ݟ0<�<��^=��T�gk�f�T<Gaq=L�<�8�<��V��*���e��=,6<���:i�#=t_��[悼 ��<.�,�c;��Y=z��q��;_O���ը<Ğ{<j0%��.�[d�tX�<�銼�ڮ���E=t�;?��<+g��b���V�)=�"��#'T=�Yr���=��";v���ˁ7=�^�;8�<�߶<�ԉ�:�<���|���;�R�� �����<ӵ�<
�r�_��;��<N�><u%�	5�5�{=�n^=��=n��<}�:��ۼ�4=�&�Wy<h0������O�D�BH˼��[���@�:���"R?��4i�������:��c���<^M =�+G�D�l=S(�W�5�7��<L�U=�z<�M4;�>�R�=��=�E��ܳ;',)=8N*=��O=�dͻ.L#�J��߼}����.<5vH=��=2_p=��<#��U�2��Q=�>�<N�g;^u=*;��4}��5��z�;�;2V��z<=:��A0=
�=���=�n7;'f:�`�A=X8�<��<�7+��=�Lo=�?�<����l=�@�<��Ў=ݞ�<��8=��6�hh=�cJ�;�=o�ɻ�}&=��B=�X:=/�,�:]�<��,=�==�O=� �=�G=��=�p��na<e �<B��Y?�:��M�0Ƽۻ6=�2��z̺�t���D4�ꅂ��*����м�NY<}6:_���e�i�k���I�W����{��),�<�F��,��k$<�"=���:��c;�ϼ!%=�n��K(<�߻���t=)����Z2=�rM��d�t�6=m�v���t=��i=��3�L=�=輶i�<�b ��ʼڎz�,��<7`Y=׀B�S�<,8%��l@=��@��5v�5��@�X�0=FyJ���Ƽy��G��;k,��&=��i��2�?�}<�<�;�<��=�f��2�0�2`<�{��׼U�.=�=zzc��hh���лԚ��'�]�-�?<�������<}�$=���<�J�<y=0=z4*=,�<��@�/]!��#w=I!���VU=73=�N;��=�H+�F�,=��<5eb�1/<��K<$q�<ٰ*=X�o���#��C=ߎ4�h�e�~��<�l7=d���T汻�Z�<�#���*�-Ů�[��<���< KȻ��<%D�$��;2w�Վ=��'�UT�"v����=�?%=+�3=��=XL=��=��[=n<,@<rv�
I=��;E=��4=l,B=s(
<}Y���L;=�P�<�,��B�;�F1��&=��a�`c�;b�W�.�==�h�<+&4���P=g&�O�=?�+�@=O�ټ�m�<�Jw�dQ���<�vZ=f=��@<�9;<~L�< ���a���a=��$�Hۆ����K�q=�����7껎�O�4�ݼz�żTV׼�k�8�Q=м��Z�o;޼shg������0�]=B�$�+�o<ƃ;�8;��N���8=x�=XG`=�<��=̹�:�t����/?^<Emʼ2�,����<aa�;^�;d5<��x�S��< F�)o"<��a��=Q`�<F��	�;V�$d1=�1={F���ʼ0����6(��_%=#=fb2����ZG<>e�\��N�<�Gq;��.<��L�Oq=Ԏm=��bd��k���1�%K�< �H=cz�;y[��D��<y2����;�>=SA�<�!����<�G<�;=5&H=��Q!f�u˃;�~z=�N�*�O=���<O�;����S&�ĸb��K��#�=V�j=��w���ּ�.�u�G��]5;Z�<�5<�޼�}�^S���<�͗�?��}j*=�iH��T�<�*=�n+=I��8��;�s����c<���<r��r9m��d�=��I=���Uqo=]J=8�<�f=�����*]=�F�� <�{׹f�9���5�ۼ0.R='p=t�=� �<QCz;��=��:�Jټx�<v�^=݆���%G�Tݻ��?=R�޼�E="��t;<SS6�
�@<��:�װ���=�1+�[��va��^��:rT=��5����< ��<�\v=ʩ�=i��O�M���5=bn�X��<T�&=c��A#u=��!=P���%C= ��*h<��X<qe-�4E�<�ī��T��͓�}.$<^�;���<;�>:��j���b=.g�:��;���<q��;��d�e��f�R=�`p��^G��bA�
H><A�M=?ذ;���<�2������<�/�<�T����<���-3��+�C��<Zؼ˻�;rO���)=�rj���m��GO=J�+��#<�E�ܰV��Og=D*=��<=����'�;�	=�@=��a=���<0�����0ph� ��</	�%P���<=�4�<��4T�J<v#=�q^�<$=�#w= ����L���+=W�f�nѾ�^\
����<��������=`N�v��<�Qv��-�;��U�iچ=�e=�mҼZp�Vǃ�q3X��]�;[a<��&�X��<��&=�Ym=<x<-Ҽ^��<Jؼ��9�>�����%ջ�2����<�t~=�4�|� =OSs=3W���K���<sC=J^�<�S�II=�90=�X=D�2�#�=��<�l�������(+�9�˺#pw�9Z���5=��/��MD�[Om=eJ5;r#R=�Mż�$(��0�Aͼt�2=a�=@]�<w"���V�;�Q7= W����+N=̼x�;x�;�##;R�<s�R=q���s��<9��
yڼP[9��H2���!���=��
=����3��]=��]=�4�<성�"z1�S�q����;TZ��Y4��L����=��=*��p� �q�=X�(�K�Z=�м5�<Sf׻�.r<y3Y8���@�� ����寮�� =^�=XJ�<`z�<�J:�p�<waؼa�A�@ �<��΂=�ʼ������==�NU=��=,ޛ�1�6;'=~�=Ռ<�<�����6=bX_��pļ���;��|;zk�]W=!L2���M=��<r���d=S�G�#�G�%�ݼ��|���6���<<�!=���y���[U(����C=�<*��/]�����<i�*=-�0�[�@�M=L?=㚮�/.=$�>����<��A==.ƻ/�ѻ��=�!=?�.=�@�<U���*��<gx8��_<�El��sV=���-l6=L� =��=�;[<[=��A�U��mW<BO��r�b
]=��#=�п<��<ʨ<Tډ���O=>�Ҽ��J�q�=�e�<|�Z����0���!7=�=0�=�h=RJ;���1�@�f=�}=�
������<P�B=6���Ȅ�\v�d�<v�S<>_E=��r=��6=ќ�<? �¤=%(�� )�<s="N���<��<��?=~��<DK=���<�>/�m0��*=g�#=��-=Ȫ��_�B� ڔ;k���D�!=Ć �7�R=u�<n��;X���א�����&�X���d��\=��F=7��g�u=�;l��N��\yC=����p��̗:��z��5�<�W1���C=��;e�=�qn�����\������X������粉<J���[2���j�!��:��<��<� r<8Ď<�sh=�5��:�S=o�F����տp=��ڼz��x�<5Y�;䨜<�/X���<������[��<�&��K�����̫9��;��Qe�"�=�!�Y�G���=��=����)���
��B��")�~��;^�H=�C <z��<I
��=��q��ݼ��m��bۺb!����<��Z=΀<,���mg�|ʏ����<_����8��G>����:�=<غ�Љ<�y!=��;ԇW=�5��i�<�������s��9��=�E�����;��^=e�<�-޼���r�s;��<k=8nR����<��\=���;��;�5�T�����^5=�?=�����{<u��<�.���D��,�˼��"<I�T��]�.�p<��`�h�ͼ�==�<��S���Ѽ�����L�{�<9�_����;���<�S�H.�]U<��<��X8S撻e�0���:\�H;���<ԛ��-=+-���ߐ�m|�@)d=(@=sv��Qe=Tzݼ�ą�5�=Z�ټ~$<���h<��?�<-R�<71F=��8�%0<o�ü��0=�沼m'=$`ռ��!��j���`H��Y�����U�ΩA=6W�q�Ԗ=�Fмr�B:l��<T6�;ݺ�� �׼@.P=h!�<O�L=�(I���I=(m����*=�r	=��	=妙=��;
��<�@o�Z�4;ǲ�<����<�⼐������< ��:�9���Y<Ux��0�{Wd<���<m =ӇY=�1�����:�������7��-t<��
�g�A=q0���p]���X=/o�����VN%=6,]=?�x<#N�����<t\˼��<Ι=A�;�0�<N��<:�T<�6��T�ϼ!<M�I=��D<�eC=pd�<�mw��$=^��<1;R�^�m6U=V�=�tY�F޼~���3�<��;�G�]&<me5=_��;��=��	��\�5F�;3"����h":p=ע��=-+9=/�N��y��	����<�j=��,=�={���}d�<|�C<|1f<�=ʵ~;`��2 ��/=d�<���;a�;�+��ѼsQ%��B=0�;t|��ݷ�u0���1պ�ᏽ� ּ��C=����$AW�4�Ժ�0;�{ܼ�<l-��	��>�:ȅ =�4�M��8{{;2=����<4p=��>�*�<�^�<�?=<�7�{W<�S=�K��,|�X"���f<��U=wV=#�'�e�f�=h_�<i{��p�<�:A=k��m��osI��[=u�D<���@�<0bL=Q�*���ؼ�x��H���AI�y� =�`=mdc��E��P0�8�����<f�!=��L<ՙ�`�A=t��EG= }󻠁@=�k=�3��6�<�;�I��<�%=���=�4�����&�<��5�5u��z��<ǌ�:�v<US��
S����5��|�'��8����;�=��p�j��_,=	L�N̼�Z˼�[��t&�=?K=�k>=�I��]<�W=J�L;[��=ّg�ۉ_<�c�X�=�|�%)�<��o<z�$� �?=�)ʺy�e=,���l�]o��NR�"�n���~<�G��|�&/=�j=�k���R��|�<V�Z<q�`��{�<�Z����,���q�<�9z�7����9�L�<t�<>��<\��=�<�+y�S��f�%��_(=r�#=�U���a�;*��z��,|I���_�;�<C��<�#����*���*:�H<i���<\���3�V=��<~d]<��ʻ�$/�3dļPN�;��=�ͼp�K��ﭻ\y�<� $=��Y��r�; `/�r��<}=9��=495���<d#�;�}��6�t#�XQ��-b�<N��<x��;�m��P9����=�"W=���fl+�ç�<*�<���;cÏ�� ������-;��<G4��x~f<=��a7��!�<ǧ�:�^�,�ֻ8�</)���@�*R�/�p�<�»M'T=��+=�Mt=�>���/=|b�<�4<��ܼ��;KHN�����<;7༈-�<$�	=T�:=n=�<��o�=/�<����K���9>��A)/=��'=/,A��S-=��":�Q���/A=N�Z��߾<�
<h�L��}=^ u=;M9���<N�p<��	=�8�^V�<}������e��u꡼xJ*�n{	��=��̼���BF���<�S�?;<}[3=�}�;w*=9�:�&��G���xB����ꀀ<:go<��<K�!=���<�=��G=�P���_C=�e����<��=��U=C5ܼ#��>F=e�'��o"�c��;=H���t�mϚ<��<n�޸��q��J�����b��t�¼ց�<V�p�FT較V3��V�8\y�/��hM=é��h�ؠ�<D�<*��<�ւ==k ���ŀ�9�;���dF��7=�=�I7���=_
��}�<�+�;$=\� <~�L�|����?=�ݭ<j"�*�<��м�@;���;��l<�i�j�	�oɜ��o�<o�-��_��cC���4=3���RY=xJ�ջ�dB<<�eٻ�/;�A=�.x=�'8=��[��K���cN<Gs�<�ҹ�>(=��Lp�<����&b����p��6<�=]Av;���<~t=T�;0=_2Ả-�=� �V�|�b��<4�8=�'�<�%=q��;��(G޼]� =���k�=��<��&=�����<�����Oc=u�=�=IGs; �-<lk�<�K�<;<W�g�<��<1�G=�m��6��K"=�$E=�z��3VQ<���i�Ƽ��=���a�<N=�_=\m?���"�<�=%��ye=����ˍ?<m���Cv<��d=㼸;D_�<����p�<��n�<c�ռ	�c=��r��G= �<``2���F=�������l]j=l�<&X��<Q= ��<a��<jx��㷶�oJ¼���*��"C�<���o@Ӻ���<��N���>=�:=��<�&=�~��E;=C�����8�#b;ro=9b5��*7�`�=�᷼��r;�üՂ8��(T=���<[�< ��T�<�a�dw4=��	�μ5�����|��<Y�)���%=E()���<:ؑ<YX��;�Wj��L��7�_'ּ��;=o)(=n�:=��8=Jߴ<�ۼa#<!�ۼo�\=�/"<��=hN�:x�=ӵD=�iӺ~�:~�;�r�=��<�
$=�)�<��R=y��g��<�	�At�<�HZ��h�;~�<��+�}�%=�@`<=2�;��O=��<�Z������R�P�[�(Bw=�B�%�;�A��	I�Q��<ĭ\=M�$�<�����yN={�ؼ�ũ<`>���/�<j����d<�L�˥�\#=�~%=��S=IR�� PŻ�t���
��)�*<�N���;�G=�O�<�L=�}M��!�|��=�@`�斣��R|<xЈ�K�a�3�?=��;:��-���=�n��Ya�Mw�X,̼E	1��=,n=xt=0�����Z��N?=��< �n=$ă��hͼ) �<������F9�����=*&��RJ=<{��(-=@=@�Y;х&=WS=�\6��� =�^y=�tt=ל�<�m-=�c�<6�o�`�<�@������*l��r��:F.��K=t����<�PB���(=��:�\/<�U��n���>m��3u=0���O�Jr���1;�9oB=(<)�����]���!=B_���P����<3���,=�Ѽs�`�8f��r�7�����L��������X=�Q=���U#�<��;Ն���
==R��ȻLv=����=�h=��W=5)V�0x�����%�g�.�*�ϼ_=��<;����T���%�#�=����V�6���d+���E=�!ɼ�껰��< iļi=�;F=��޼�;�OO<E5���=�yl��P��F�>=>/,<���YJ�<[O^<�cb�;4����>��:Ǽ�bq<�E�<�dּ�R���3�<�j�/�Q;�"=��Ѽ������?��=9x<2����1=�*U����<0R���Sq�f��������^=�Kj<#��<�����8��-�k�;�%�X6=��K�B�8<DXḐ�ɻt�\�\P<,59=��X��Pt=��<�L<'���f=j�;����a�M;�&���<<��b�q��<Ub���,=jjm=jY= =�;�&=��m=�6��$(= ��v� =��.�Ѵ�;&�����<^�?�s���|� GA;���UT�D��a�;��;-������<Ѽ]�T�nd�;_�X([=O�<�_��~��Ǽ�&c=SD�;
K�B����� �һ���/�	�};���-�����<'�;�}��<��E�>��<4y3����WT����J<?��<��
�V��/��p ռw9N=�P���J��?<�'�;9#�:�-�{"Ǽ1i�ÛQ��fB=[/r<)�,���
=ȕ6�qQ��Ƚ��,����:Q������<]N�Qc�<#�(���G<��=����݃;����}B��i��	=^6�\�5��*v�\���*�w�)k��g<��E�O��<��_�Uk[<�
1=3m%���%�[l=�,K���-9څ;�y�?�<4w�;(�Q����9ݬ�`�O����<Hu�<��S��M�<,=v%u=3b=b&�;O��W}5��9f�u��:~�ʻJ�= T�<��F=��F�Y�<T�e=�J<��N����;��4�����F�:�/����;+p=�.�<ʚ߼�4=�����h�3<�9��ռ"�7��<b�:�� ^��Z�=p	�!�� ���<8�@��k�
�R�OZ8=�@1�$�=�V<��%�'$���u<�%���
��=�ms� =���<��>=��F<��C����@��k�:G^�<�߂<�Ɍ<8t��.b;��:=�r �v��<�����<1�L��{=zK6=\��U��<���?�T�"�5�eܼ��/=;���p������<��;��X<��D�+=���&=u�c�Oժ<��,�r >�Y*R���<PE�q��<��-=4\;��=%��5��sX�<@�:,���4��a �b��;/���E�<�Zh�lT�5-]<ͻ�<4��}XG��?���,=�<#��<��)=m���r�<�/D���H=T=�p�<�	.<�Zm=W�D=�sp�$
�=)�b=��5��( ������;�==j�v<ˎ�>=�ϼ����ϼs
=���<J/�D�[=\ ���F��O<��Z={�<'��;pJ�^�L=�����7�<��/;�3�<����T�<YZ�Nn˼��=�$���n�<��:3.1;�o����<�쐻�'��ﴼu�9�V�5<`qV�]�<d�=4��QE=��<�7�/�^9��ļXHD=��<@ 	�{��<���<7	=L����B=���Gv2;l/{�^�����q�=�!N���;G)�<u=�<?�d�cWT��]��r��E���K�<}d?��%Z����.=����@�PP$=�CP;�(z��Å<��T=����t�f�-���2�-R=QO+�����^E=��0�{R=�n�<�[N<{����o#=���<ͧɼ��'�Y��<�X����`=�us=��E����$�:F�%e��'b��+�0=q�<�V}=#�<�P�;�L�e�<u����?<�����%߼���<mn=����b�<Ae�;1��<��C�/�
���;�G=,��<����Լ�@I<Gr�2	L��w=��d=`���=�3�Y���jn���e=B�<WG�<��4=g�-�~zH=����n����.�g��<�4�;��O^p�[LM=��b��P�<"/�;)F�3�:� �<�FϼN��<
!@<����<���:�L�E�V�%�<:�[�)�Ļ-D@���O�c�=89= o�=A*r�2q�������=�
|��s=�ƥ��� =A�O��Ĵ<�2u;�XR<h�_�ex=��/{=!�<<�¼&�����:����G:�<��<D��6%��d�3�^\u=�����X�T�\�AB<'�b=2`:=�lf�f:����V2b��H=2:f=����\=Sl�����9<U�$=�_)<�L���9=W��JS�����<��X�&t=�tؼ\�Ｃ�}=�=�����2N�y�[��Z=rWQ=���<�=v҆��7�<!�����;��=Ɣ=�`;r�P�C݅<��ƻ?dC:>z�;9$�C�<���=���<˙�<6�<�m<��¼�T�<��������K�<�"V�X?6����<{����ʼ:ȊU=��]@�_�!<-8%=�$�eT����t!7=���<		�;}�\��}m=��l��;�G=b�+=��m�*�<X�ͻ8)n<ͺN;�KA=g�{;�Yʻ5��9lW�<�����{�x�<=<�	��	?<{5Ҽ�y�<�;�<r�H=}K�8;#���K<̲�;��;��I�h�c��fw=�$=�W:�F&<�=���P�=�nI=B:��K�����Yr==�(,��fH<�X=�Ȭ�2�B<�F
��@0=��`:U�r������[ =�JV=����=�S��ư<a�:"aw<�?��Gݿ<�z���ӼV8���q�:�O=+�j=�f��Ա�]o=���9�`�+�J<�м��;d�$���*<�zL=�&U<F+-=<"�L�+=�_���z�2G����w=���<>(�4�5=i�H�I�}�(?=�3t;oN4<�H=��-���;ח8=�IT=(�<�p!�q�:w.�<���������;�?x=}���N�;nv���nm�6���7\�ί�<�O��=�C�<�R�;�!���+�{=�W��tt��~<m����;)�=w�,��M����yX�;��-=ۨ8<zw6��x�=�@= -=ܠ ��5S;t����<ݟ߻��+�"�d=,�(�y�S=X��^�;��>�����ǽ<B���|���E'�
5��c��==�9=��=W4U�+�=&�<�����o =,�,�r�&���@�@�?�(�	�w����f=�D?<��<-&P�a�$H��]gB<�T�mS��7�=�w-��&=�cT���<�=.�[�`fv����<�������J���r����;p��?�?�M��<s6;~�5�+�C�͞�����R0^=U=��<��<�D�<�>�<���=|��Y�1<<�W�~��q�<�\=ؔ�<D\=̃.��B-�~�;=f�9;ڨԼ��<F�E=M$.��t<�����=|��r.���	�'�˼ݪ�;�0�<Ru*<kP�;g�i�!�>��<:�j��<o'@���>�3=U�茻߄���-=�;<x4<v'�;�&=��e=Ӗ�k�2�����"=�/f=J	*�4��<�H��G=�R<����L��v�;�+!��gI=���<$����<l=!�$=9����� <��;`k=�f7��=�ռ�s��h@�?f������_����1��uC=�\�<H�<��V��(�<(���<l�K�Fs��V9Ǽn$=~SS=��ݼ]��� <Lo;����T�*=�%�3»��i���=?3�<IW;ǂn��T�<���<�g9=ڹn:j�Y�]���?;�!=�r"<:�<F'��pݻ�u;���<���<{��<P&5��qp�[�<�x�M�]�$��a:�ܠ�B�:=����/��W$���垻}f���C<���x����<�W<�ٽ;lk�D�l����<�?�<�>u�A�<N><�~O���<�W��y�uK'�<8 �$�'ZC��(x<z���IL=ǦR��	�89��rB=#I"��}��a�<�j�<�r=�4$=�p,=lz8���]=B�+��Q���;�O���:� 	��W3���=F�����:>N<�����5=�f>�1A
=��<;�<�<I�5=��<��%=�s�;�,�۽�<��!=�L���6�����cJ�aٖ=F��<z��W�V=�n=0KS���:=jXe=Q�u���9���ڼs��:����#ѻi<2�n�t=p^p=��=�= �������v��;��w�b!�ve/��c;ܗM=$F <��<b[=�(�H��������uS�<�S=��+=K+�����E�s�=�f���ܼ8ﻕv��`5=�$�<��7=��<�g��z��~��eQ"=X<{ӱ�.
=�G=�C�;�=�OV�i�4=GC�<n�3=��Ҽ�pG��#�gI=���)i��M/�牛�n�-�!�ۺ����;�I%A�9<�l<s�<�\g��~�z�<bn:��=�����k�V#C=B�H��Q�X?伮b�=f[�;I���د�<�#j��w=�[�U�軚0=3.�<��=\t:=Ir:�.��)�0=��<�t^����z�a�b�G<ؑr=����($:�G����<h7�<kp*=�6�]oV=g���{^x<<��:�"c<S�m����<�ُ��v׼��<~d���\=�2�<�,�;A"I=��O�s=k�<�t�;�� ����<O~���C�������a��<;�o�<e͉�**����<ж�<�-=�:=^�0���|=$�/��3=w�8��eP��94��Qu=FM�<2L=�~�<4�v<,n¼C3f=�&.=�� ���=MA=�O=�	�������<h�;�3(�Bc=�β�H�d�`�_���H?��*�$�м�H=}��;ۓA<E餼L=7�E4��?�=QQ�<�jD� 	�<��	={�]���;��Y�=w���Z;���T�+�ļ���;0�C=Z<����(к����<�U=��(��"=�C2=�F*=뿼㜛<Z_`<�j��gC<Koͼ�U���<�(U=��м���<a�>=V���b�I=-X�<��`����%o<��Ӽ�"=��ʼ���<Jt�����"$�3ޟ:C���jY��a��{'<'�<��/�S��v�V�/�5<����P�<r��=��g=�����(�<|i2��ke�������<�oм��*=&�=87��;�� �0>?��J=��"<՞d<6���N=+5�;Dhl==%za=)���ns��P=�P���H�:_=�e=n�<�(��<a���\X� 7<J��<�,	=��{'�<��L<�k�ላ<�L�r�e=��C�i �<Y�Y��5�z]=�!=�h2��s��=)�ƚ3=�Ex�������(=�u�<j`�6X�8B�;���<KU�+��FI=r'=w9���v<�=��`=��t=8N��=(�;_?i<$�<�<}�
=/ꚼas�����+=��G
��*��|54=��D=X�d����;�#=i��eF���8=�=9�5/ =���<�O���j�<P9�;�{�<��N��wO=m���x&=*����'�<3�7��k�<���~���5��<�>�;���X8�[kP�G2�ON=��^<~/O�����ԝ<Y�=�"N=���A��<G�P=.�S=�=0��d�<��Y�LU��f+��G�<���:�E�=y#���{���¼<+�|�s�=c�C�A=�����<<���!�<��8�^;��M=��{=�Vg��\#��a&�:~߼+���Fx�]$��dT����?xP<ѭ4������>������=]����<a���y�;<�V=�P{=7>�<������<�xg=J6�<Ķ������%=Mn'���j�6�=~�+��t��r��Uq�<��<�:�%=Z�.�G{�<d,$=d<=�'�;MC����T��f�r�C=R�m6=�i=�����Rʀ<Jv%�+�;E�<�N=4�o�S�Լ�a�<A��<�7��6V=wq���s��>�kY�����<����b!�<G �<���ӛ� ��<��m'T������dX=�9�;x�<���:�\=,.V<��L=�����T�߀A=����I�5;����H$<xU���k(��=.;T����}	��Wa<�Yd;V\�<7t�<
�z=NP�<�T <��</��=�W�r�(��<��G��)<��X=z�S=f�)9������8<Z�C=�伱����Ϳ<v�_=f�c=�:.=Xخ��Y<ǝ=��R�e�o<��=,Ǽ)=l=mD�*�;X�q���]=�9��V=P�@=W�ּ��C=��,����:r�ɓ\���=��B=�򰼱�=~�x=y��5zz�.���u��;�r����xe*�'��I݈<Үv<�$����W�<��զ��6=�iU��|���"=�q�:�2=u��<)��߳;[��"\��u=�=�-=d�<�&=��;ǲ��`���h�o���[XL<��?=�n#�a^��� =�cy��$p<�>��D��xV=�_%=�J� ��;��N=B�<Gv=��<�LH=Ɋ=;?��ּ6�>=�=8m꼓�<�����~x<�4Һ�绥А<I+��٨<=�{�<j;�=�>����<�\9={Gӻ%�<:N�<��W=�A�<�ʼϾ�(�f����::�=�Ƞ<�}=B�<�9��X����=,�ټ���<>�<h�Һ��=4& =�5���2E���T��M=�g�@'��?�;���<_�=��>=7ِ<OZ�<Sd�g�n<��7��\���xu�!���D�:��?&%�	3h=�f4=��@=�������<t{;�,?=	m$����<&ǀ:b�����<�"=��[�`�߼���<�Z�<ol<S@'<Ƚ�<]�-�[q4�5y��}.�<IoH=EQ弑/�;~!���#�j��2�<Y�}�=q�o������;;�(�&���x��A]7��������������ր�DOܺ�n;>��<��j-�<7���F�/<��R�<15<>�<+F��e"��Si���<���<ę���a��CF��}?=�H1���=w�M=i4=�!l���z��;C�=o����l�/������89<c=� ,=�A)�IM<h�]=�~��x�<�7�=���=��h<�R<��=�T�9���;Mռ"�k<kTI<i.3;e�<�q�<�Y�TO���V���μ,$Q�Q�=Xm9=� ���ڊ�R�c���<� <�~=^q=�O=�%���<<�~���=plG=�<4=a��;�� ���`<֪¼6��;�xE:�mG�s�=_�u��:;]�=�-ü����-#=���<bߛ;5�i=\����i��|�����;��P�a�(�k�X=w�=�`o�8Ϡ<Sf�<��=ª�<��<�/<�<˟.=f+F�e�)��%�ł\�t}=rղ<ƛ�V�S=��<�ǻ'm=� =5E���=$u,=L����p�(��[����¼a0���=%� =ɓR�
�y��f=���;����<w�<��ĽO=��O<��=�����ü��6=��0=��3��7�w��<��5%���l<n�0=��<(��<�_�m�8<'�F=K��dC�~�ż��!=��O&=F>G=�N�<
�=��<YU���<�5;����I&=[��������%�A߻������m�!�h�mk=3ei�~.m�y1q<�����<��\<V�T�Ĭ�s�B����J�P���H�����e=J�B��Ig�f��<��e<�D��CD=+N<��;��0�W*
�u=+���>=]��<�=�(!=�lE��'#;z{=���� b�EGn=�=�;mIj<�J��,��
��<</�<���<`
<���<3�S�ԉ���/p=����2_��\�i�q��<:4�q�<�F�wC�eO�����<���;X�=�D_=�+<�e0=t�=�Os=�f���޼��<=/�;�6�;���<xy<���9�߼�λ�?��b�ও����<=U��&S:=�1�e�N���
=��=Jtq=W�G=7�;`��D�W=����f=uM�;*��� 1� =/g�;�a�<K�^���?=��ռ�!��#���y7=� �'�w�I��3�����A��<HD}<��k���Լ�|:���=��<^��<�0E��&޻�+�;��W�}:T��<�ػ,��<"͙��rN=��`=3I=d�p= u�����'O��Oۼ�ܞ<��E=���<Dq<l�=�Q=��<��=+=��O�=?���b=)t�<A��<`἟;I�����!H;ȥ��~��<�ἉG���i�0�%�b�m=�����Y:<����ﱼs�y<�𔼎	;�8"��=��<�����ž<�������5*</�T��Sf�q:z=�� �����I*��R<�_�)"�=8H����c<n�?W	��&i=�Q�;��(dE�xb׼�q]<����枼+����<琢<�=�=�<e���<q2=�#=YB7�y喽�	�}v'��1V<I&t<��<C�-��̻�2W��c�<_.=ܺ��N1μ��b;C.μz���-ZA<-� ���P=â1=9�a����;�K�#=4�*��<�C	=n�/<@�<Q�[�+~�<hՠ��l,=,U;��C=��L=G�����n=�? =5Ma��X��ּ~�<��E=��<G5��kb��R��@�#=ʈc=.�m��һ�=�}=��ǵ�V�3�AG �K��'�2=cSX=/-� =g<�T=x	~� �"�!1�<L_d���k=�Of=�ʼ�24=|�Լ��=������<���<����j�<��0�)Z;�ĵ����Q<zT�<K�=�2=pӴ<|��9E�;�<=(7�VO��ѣ��ߦ��ML�oI6�JH(=k
=���%H<�"B�MC�����p�;*�D=!��,oB��b����=x�h=U�=ƻL[<�1:<����X=໪��~B=��
:o�<�"&90=k�%;籹W�}��
�JO=g�>=��6=T���=�<
�k<��>�Z���I��>="@=���<d�m=�J'<v�K=�J�E'��B���<��,]���g���㼭��u��<pK[=�ǵ�Kf��6⊼���;��!���,�{N�@� ����;�9�(�=���<��q�̌�<F%>��<�\�*�b}s;'�
=�pY��E�<���/W`=���<�B���vI=�~#=ɕ��q���'�	=,�&5�O��<�3��q=��Q=?u=���<>S�&�<|�&=�}�<V��<���<}T=��D=�o����<��,<b�m��b���.���x��%7��QO=�z��G=K�<�%'=��.��kﺾ���ֻqZ=�� =)><仵;b"�g�;� =��}�9쉼��%=m��;ռs���λ/5<=�8�::~%=6;=<aM�G�f=#��8�Ƣ��.�pʋ��f�;�,G���0v,�B �{ԝ���c�-�=�f=�f��ּ2Q�<n�<���<�<d=v���0;�� L=lG�<W��<?�=/��A=y@=�K=%0=��<K2�m =<�>���=|�f=*r��5"�=��^���m=ś׼�no=OcӼ���.�;���vK=,��<RtؼG�=�����<(����<\_λD	e��� {�<��=�������=���<�<@iU�f��<����m�gYS=��N�bqT;f�;K�
�WN<�Y�<���ۯ<��>=ŀ��C{�����^{�=�ͻ�:#=������	�4�C�#���W=��dU=���:�i�<� �<��<{��o����<����:���3=��ϼ�r�<]���l*E=��y�J8�n
=̧w=U��=+|V�����.��<�Hm���<ɇ�;�?_��#��R��J�<�3]=��;�q=�-�<��輜��<4XG<6���0_=[����<���UJZ=-��;E�==7�B;k�<ba=�]�zr�;d�<���<����ܻXպ�C-��<��$�4=:1���D<�]0=;�=dQ�<d�'��G5=��<�y��<��6�	a"�p�=v���=� �[�弾BA��X�<��=4-1=i�^<��� ���g��^HS<l"=�t�<��TK��E4˻5�d�m�q��7��:t;�M�&B/=�;ۗ<F�@<Pj�<ԣ�<$F���m=URȼu�μ�<{��Ai=�O�{���<�"C=���<���?���@�<=��A��'�<cX=<e<��<�<>�	*`=�}@=���d==��̻�+�<b�q=����փ)�9E=Vm,� �A�9cƼ�x=� 	<ᾘ;�yl�b6=�����:���	���*�<Bc9=e��Hü�L<P� =TQT=�t�q�<��<���n��&�<:0=�P�!��퍻��P=}v=*~�<B=�W���8vi�;�4=��)�z�=��=�����a�����/jJ=� ��g�y�<i�|�k�J=�3�<�����+\=y߼�S<[�cB�`�켖@o<|0�<5�;�5���n;�w�<�91�J�<�"@��B=2�м��$=�x.=�S����x���4=�U�<��=��a��2P=g��<ҡb=ag�����C�;�ۜ���<2$=�`�<��ƻI;u���x<2p=�zi�Ӏ�<2���L5;�O�<�i�]��=Z��9����:��u�<������L=��L=���<kgD;��̼TE�K.�:&9�s�3�V=j���P=��-�C�H�Z<�˵�0}<{=�ͽ;>��o���ɻ��$���]=d-A=7�]��$=?�û5����N0=�ޣ��z<�Y+=9�>�E*�<{r=��$=�?h�0��?�;9��<�㼭�~�\࠼Uy��*�=��A�TQĻ�=�	�=Nw'�����!=���<M����:���=��;&��n�$�&�@=�e*��}��o�xO�j�Fq+��r �H=~�<&Oh:���<�f^;˚�<�&1<��s��VƼME=��]�E�(=f��<j�<6
�KS���{<$a
<V5:3��<��ɼ�;��*=��F�f�3=��<F[=�`=��<d�<4�;��r������f����Sͼ�I��y�$=�=q�;=���@=H=�Ȃ<��w���˼���<�9���p�<Sb�ʶ=�<O/F�m��;jq�<Kn����ͼ��<=`M���N�:=��2����@1=`�B=�S���X�<jI<�q=7uѼ��\<b�<}��<�JT��Ռ���&=K�D��09;u�=F�<y��V��=.=ˋ=+=<Ew=T�|K<��v=�s�<t��F�G�����ZAu<e�o�>%��缑<���'�?�N=H��:�w<$���~X=�w��A����<��<��[=��`[b=���<���<���<�+��s��;g�<���<2��=�� ;�E����<�n3�T���k=ɪ	��/=���;徏<�*�<��=�9�<�P��f]r=��$;�9��'=�<����LR�� 1�5S<��xrQ��J�B�>;0Hi=wlz<U~���]@����<d���jȳ;��=��+<\F=߲�:�ӻ /S��f`=%�/��{0�(�;�N�y�,�>�V=��I��/`�`H�<R;�=���<��=��	=�PU�.��;�-<�=.�S�m	��9�ôS�6�z���d\=(�<;��<E�2<��<��f�m�<�U��;z��
"=��=�p������=c�MK=v���]�;��<�Lĺ�./���8�<=9�:)?�����<��<0�ʼ�p�����X��~��\׼;;�u�F���7aw����=��pn¼��=��<tN�<���<Td^���u�Թ�;A�,���$��|+=RI)��Wj��݆<.װ�U���/=��ڼ�kH�/I@�21=~�������䆼<�=��<��＋��<�L=2���Z��\�����R���L���\=Քl:�\�;lt�0��<�b<rY\<q8k<��H�\V�<!��i���ے���3�R�J�t�S��
=�v�<'�=�L�ǥ=�T7���<tLj�V�*�f�'<d�R�t��cO�;��.=i;=*���铼e�;�ל�U=��{<k9k=,Q���N =��<��Q�t)z����<98�<�+>=�c�<cB��_�a�����<�4/=q+g=U��< ��<żȰ�����#�V<��==�J=�����ȼ1=�<,��<j��+ݻkYu���8=�^�v�<:pļ��ݼkն<�9��,=�0 �s�\= �3=�Q�<q�b��߰<G���5�������;��<K皼
�;��<5Wg=���Ű9=m�z�/�1��<+�����<N��;�0���]=�)=�\=+#�x��?>�Aw�ڇ=Vf:F*��pd����6=x�:��+=��\<�켨���E~=ʔ�<,���(�<>�<���<�����9=ے=v�<���׼��=R�(;�C=\�B=;.=�I����,�J=�[X�<w�Y=Bl8�� �<�A���B=��tfʼp�E=��_=ͩ<Y)/�-�=ׯ�<��W��������#��K���=��}=Ny7=��:�˼�et;���ʈ=on(����;7�D�ws=�����=<�����x���<�ty=��̼4ỗ�G=��O�� ��X�i��x=0+����.��1ǼK>�ϵ"=�s������t(��G[�J�K��Gм_�w;�Y=C'޼��3;Чa��	����������2/=� =�Z̼*l?=f8z=z��Z��E��<I�D�J�	��{�;����;J�ik�<��L���<q�5��"��V=0C���V=�`=���;��<�[<Vo<�m�:s{���λF�U��o<7�����;K����L���lk��k���΋<�ƀ�^-%��x�<FY����\=�蘹ck%<�]����^�o�K��Q��(�==��o=9�A�D�;=q�6��K=�~4=;!ؼ�Nv;��=�X�,�<��c���=�U��"$E�@J=E���UP
�kS̼-QK�!ܼBS�<��L�.����c��R˼��D��˼�v�<�����Q�n�h<��A�$M��Χ=�Z �Q��<��)8=]>O=KB�<�%=�`������i=M<]�3���=	�4���g��\�R��>T=~-<��#μ�5=g&Q�W�/=ťr���=7$;<�Z�9ғ<6G��7�=������z8�<JK9��м�G�ӂ4�+
���4;��u�)X�<@��<܆�g��<X4ٻ�#=ޞ
�\K=ӯ�<�Kc��=�P�~=O�#�f�<��� �d�)AH<_S2<��=����==�=������꼎�=���g=�=�%��j_5�W����%�<%����Ժ1<<�j��1�c>=B=�"<)�;$�ϼ��޼ON�;����s%=V=�ӻ���<߾��3?=˟�L8=�h��?�<D�!�r�;��=1��F~0���M��Lܼ�G�\U=��%<�_=O�s��7�j 2=���;#�ɼ�8y;��8=���:_嗢"�0�=�b=��q��#��
,�l�����;T�z<ז�<!9$�)߭:D`��$Ƽ���<������;1;�|K��a!�`܇:T�=��e<�b�<�h=4,*=��81)�f
ۻ���\�=_4�<0�B=��s=<���2=D:E��Q;0]S�|���Z�w�����=�;��#=zw=�G=qP=����i=��(�g�q=l��C!��G&c='�
:�F��I=�H=d=*�U<hl3=��b��6����=��=q]�;Q�F=p�ͪH=�K���K�����鬂=0�<�R��dW��߷��	'��R�<9�V�#�M���ݼ8U�<]lüĲ>�I��<q)�;�H;�Y$��k�$�=ôM��K�<���KW�1[��@���ӭS��tb=�D�<
<�=̼�=�PK�˾��,�=��;R-�<�#V��V8<Yg=a�?=NV���J�g��;,;��G=�4�<�h�<� h=s�E�\��<W5&=b�s<��R���N���hD�<̐�=4��":�~H���n<�b2
=��ٻU�=w�,�r�3=}Ǘ<��#�4v�<'��<��M<����7��;/}�<;�`1A�i�h=Z꼊㿻�N�<xd=VW =��-�<�X���N��x�<z�!���F�J�a=���A�0���.�Xc�<s�<jB�<���gi��:P��ZC�#�>zh=�0=}G��?X=�n��U� ���P:���ʼ#C=�*%� A׻�)�<
W=�^i<�"o=�8�;��?<��c=6y?<��z=��*����w�~=��<=�gy:#���Ƙ;��^=�Q�<�>=�f=}�º�S�;�=ʼ_�^1~��*�����9�\<�p<o�<X�Ѽh�==�ͼ�e����_= �f�$V�(���=��<�;�b=Q;<��׻|A��׀��N�u/��C�Ҽn�=�t.=O�0,>=j�2=�%}<a�&�Uk�n"�i��r"S=H����1<ID9�w2�<��g;ͯ�Z�9=�饼�ռ�T�<�K6���K=��^=�n��
<$=W=�fE�^�T��S}<B��f�S�a�8���|ӼAPK=��C<}�*=vXE<�c�����\�����w�=�첼$��<w�i��/I��|����<"$���̼�����4<�}���
��u'=��S��?=�KT�w�<�(=���&��}�<���<Ghz��Q�<��<��Y�U��:�^w=)U.=^Ӽ(A���P>��Qi<�t��wf\=l�.=�vQ��1�M�J�݌�<�ʻ@;j0�;�]�5a���$�<��=|�;m�O��w#=�)=�B�<�]��:m�H�S=�t=:�;0.c�+b<'�]�s�J=��!=��6�芩<�Z\=�s�<R�ޔ==c��<`=�5�q�;>�<�m���<����6ּ�*�<��>���'=��X��9�;���o�; H,=�5h�M�G�ThA����<B��<Y$=��۹�!��_��;O�����;
<`=A*=��	�4�5W��J��p�<�`�LN1=7Gi�I޼æ��R�4�m=��c������Z�<z�j=H����<;�@=�Z�<?�G��ܼ�Ŗ<h=�����w=~)L=��L�dS�<pK2=�͑<552�v�;�9
=�H�<�7=��(���U=_l���<@�Z=#�Q<�ۏ�}�F�/�.�2��<h�=ހܼ�c�u{c�-��C=��=� �j�W�g����=q(+=}GV=�U�V�tc�<p[�;U6=J�<����J���� ~�u���M0�!4=�$4=�a=S*= ����I���<��,�z{=vмw��<i>X�A%��t3<Z�<:~�<,-��t<�7G;��D;]��Gb[�|H;�+=\]��5�5M��5����8��
F��<��<?�V���/�E��� ��<�����Eع�K=���<��='a�!/���)���}=��A=}�b��<;�\W���,��H�K��]�#��ʼx8��K�GKd�8^��p =�ٜ;;0�d��4�2���I=��%����f)�%��<�
�<"Լ9s[��ۍ���-<4��<��/=��0���L=u�<}�T=�4�<i���e�s��}��L�<J��7�ݼ�=�:>�>=}1�<�Z�nҼ{����2=��<?=.@�*2���<���
���
<�='=�]��1��<�5=p �;up=� �=������%;�0:�ݏ<�6�A=�2O=g�)�bżkL���<]t�:�,.=We��L!�Fl+=�μ!� �n`⼟�a�{=�E ���<�a���_a<�I;ӭ<�(�_�Z=�&�e4]=7=F��<�E����~���x=�Q=^h�$��ͷ3�~K@���x<zܹ��G="�<��h=�<����
�<�H���#$�2|Y=��j=$����
=ˇ<μb��9=�(;;Wb;��<R- =ʎ#����X�v���+�k�9�ʞ�aF�O9�DT�Q1?��|�<�$�<�z=��<�z6:�{��H4=�5e�[���r-�>ϼ�=�=�ʹ���֓�9?�V:����<:S<}}k=�=�G]����<ƛ��GO��=�MK�2�;=j'��ve���<�&<hP=�հ�oC=�<��|�<�E$��Ls�;�n=u�=w�<'6�t���r�	=9"<<����;�f�&���9<�N��CtE=��Q<�Ɠ<�=_�<�o����<���<q�w<*9=��@��I< b=���<�����F��4-R=�_F<(��<�z�J醼tU#��m=��\��Y5���-�:0�=�
=Qi%�ڝ�<�O�t��<2z.<���;�C<���=�-==Uxl=��@��=�}p���;L5g=�O���=0=rҼ���<��ü��߼��>�$5���=���<� =я>=�O������B�<~S�mKf=��V<����^
j��3�<�z����<��<̞�;#�<c܋��"�7�ϻ	l���=;��:���<sv �1�P�C�M�9=��
�^.`=��E=^����<�~^=��=�k�;�[�<l�����<�
�<j������<��ڎ&;��Ҽ{�_;�za=<�Z==[��^�����;���<a�꼙E�<�{�<�/=r�H�ʼp�=�x��m��~$�;�r��;��AP%����=��.�����sO=��8��A���:=��ּ% =⊄=$\�<ПT��P�<�#;�c�	=	�,�։��V'�6��0�T��z���}=��<�q=i��Q/��!��]�<�܅���m<�KO��A[=);=��X<O?=$�,<�*�I�m�$�'=�͍;��+=��z=�|!;�帼�P<Q��;o��<�K��V=���9�(9=(��<�Ђ=��c=3s��*��Ki<�5����XxĻz���g��H��n}~��Q��%0/��5c���t��D���������� �<_�<b�ƼB�J��������\�<rB)��J`<z/N=�����<����G�V�<�V��۔=O\=J�<�̈́��Ǽ�
�<O[n<l���|$=V��<�/=��@�:�K���#=ߠ=�5=C<u_r=ٞ�<;{*� ��W��< 0�=a�;�O���m���~={�����b�=��:������֔<�~=�=�A�FN=�1�<`��J�нN=Y�=��Y<����(��US=�90=�]���?U=#3;<ڈ=�=�<�p=�V;1j�<�m0=p�����<��K<t{�����<��<H
H;;��<W�(�3YS����!��<�<�;ߺ-��[��,e5�|\�<<�C<8f�<��=p	��W�$�*=l�Ǽ�A���<w���l%�c=�3�۹W<}D�t�`<; �`Ф�5j��"m<������<Ԛ��U��1���t\;c�;�Լ�E��-�<V�Z<IQ�;��C=�r=Y�U<4M=��޼9��<fqA<��2=I[_=�>=�o3���O�s1��FC�-YJ=!=ڼ��%��TC=�O���SW;�=��H=)�<��"<Rd��a���T<qoټXY<�s=�q8=g^��o�A��+�<�*�<1h4;�Ȓ���9�KX=�2�Ճ�<�j���@�IYT��f>�	�-<�xV=79x<�����<i�<�9����3=&�'�|<٨P�Y�
ּ��<�D5����<�=Րἴ�n<�f��l�=�F������}�Z�y=��C���4=
������<��s=��?=F�<8+H=�i=��*=�
"<2�<��v=���<8��;�����o����ah8�u���2��<�\Z�qN��"I�|�=���=Ol<�S=���<�^ĻW9�;S�ц���+�/AE���x�<�M��
=13<KP=�L���*:��<�`
=���<��<Ibt<��.=�/=�!���L��R<��S%�.�ɼ}l� ����,�<�<�S<Bf)����C=��E���=K0������`�N����#=I����<����0��=4QU=�]����<��d��5�<jpS<�]����s�=���'�;y����j�=�K�;�t�w��<���$�W=�U���3=ޫ"=�0�G���M�(=��W=|ºu�켊�����$�\��S`:�-�Hax=x� =FlA�j+G��7�W�,�35y��v;��2�'�[=��<��-={�<��Z��H=s�c��7��R=�x=A�1�aO�9��:��<0�<?Լ#�<��K���S����:��޼����SSz�Qk�ĄӼ�@=�oм��������<
�k�D�X=0�X)��g�;t��<C���1�y���y�N<f�䬻$���U��<uq=��r<�{<���<.� =\�l=�s,�H��<TE�j��]-x<fL��tCW�2�=��=��=�I�#:\=Tjf=�H���<�������AC<	�<�5�<���<���f1��4S��&t�~���^M<�g=��_<gx�;y� =9�ܻ|E������k<�/N=�Oμ��<=B�;�U;P(����Y���9��^J=X�@<���yoK=~�;�;=TG�<��F=[=����>=�s=�"a����<U\=��z�z����F���a��ɬl��XT���0<vM4=��'�1��<�m���z<!;I=g�=t�<��D��[C��������<��<�����<8���G?�v=���<R�=(�=d��C��<F6l��'=��=mf]���J=l<�%<�Tռx�м���-�$=[)e=q��<>�,	���&<I�P<�ti=�� ��@=C��<��$��==���<�H���3��E���;�h��c�!=�|N�b�Ѽ��K<[=�1�:�ɼ�*�j�J����<Ǻ�<6���ܼW�ܽ?��o]9y�;�ې�wK�<ҩмɷ=8J=y0.=~��<���<W\��c�l�h��<������������;��>����<uN�Ck�oͻ�=
=���<�Y,�==�4���K=c-�<��*��WT=p6G�1k��RO=L[Q=I _=_�N�-�>=8޼�hY���Y��co=�8��kh�A<�,߼�)�!�Q���q������p=D!���{:?cʼ%	�<���<���=��<��<�R�<���:wC��R���*�������/��<:g=�w_�����.u�<X�Ef�M(�<�
ۻ��@=���<�N�F5G�m]��#=
�ȼa��z�6=�"��:O��� =`h=��O��y����u� ������s߻�f��_=ַI�(�b�i!����;��z����.=�6��H�<%��< ��^/�ߒ�;��=�����ż3B=�.��]�	���O�i��<�Ƃ=T�C=��<k��>x=�k�<.�z=h���=5<p�O<��}=�J<6,0<op���`j=Հ�3����:�.��<s��+�=��<�. �d���
���.��z��y{6=r�+������x=�Љ�VM�=r^=e=�䋼g�f=pi�<������,��@:���;�ü~�=�C`<���;+��:�$�(0=��꼌���+�l�pz<�0�S:���sN<� ̼	ƶ� 
x=;M&==F�{�m��%�=��?=U:K=G�<�!�"w�����֐�� =N'�捼����C�����ġ;��M�~�~�A~q�#�&�O�24>;?, =P=8�L=SW��b���q��-@��d��G�^�5��ղ;)��l���9F�.�M/E�*�<j���L=Ȋ<�
���Np=X����x�yǎ<7�˼eɉ��?Y=$�e�B�ceԼ�}{�p=הM;�*���<Yٚ�Ca=�
��i<��<��-�U�&=_鑼Q7I�%�=u]R�S�;k@ ��Z�<4	==�9Ĥ�5K2�ܒ�G`�;~�g=�Lx;@C�<��4��JF=Y���<�䥼� ��}޼
@���	=�m��Q�7��}�98���G=�����:=�	=��~<�-=1�i���;Җ������n��5N<��Q�����ʼ��;�
���缼	@=�w<�ϼ5/]����<(HU�)}�<�"��RZ�<�9I���Q���]�M:
GH9���5�L����.x	�o=%Ȉ<��=L-o=_�U=*�r�k�<�I��a6��F"�V����8��˩�6���E.;!;Y�I1<�l�;�.��@�%��`��R=�M(=�o�:���<��?=E_�;���<;{�<`[(=U�0�.�ռ_H�aХ<h�<��
<\�o�4�-#;_�#��_K=�$���f=��6�D�9x���=�3���G=�̛��%5���<�=�f9���'�������<t�ɼ��<�{{;�ߟ<�@�<f�K�[A�;5)�;	�<3�a�v��i�<����X;�7m�>q!��^���z��<�e�;ꧻ<2%)��~�2�$�6"� C;��m=ǝ<�1=v`t�(�1����;�Q��>�^����4���>�پ�<�rl;T6J<��=�s�;��[�����O.�q;j��b��	�<�"y�d��w���/J���H<�K=�%=\��<�ZA���$9�`=:@b��kH�D�>=�f�5�\;X ]��g^=]N�<�p��Zb�%4��K����]����;8����Ҽn���#�>�OR5��=�k(=q�D=� e�����s3<D@=+/���x��Q�<\��#nj=�����;-��7���&��:C��TB��e(���'��g�<���<�y����+H�<U��;�����R�<�)��$=i#=q�<ǉ<���<�4V��K,���H�� =�����i\����;@�ּ���;�ֳ9�<)=���<�:Ѽ�B<��4=�v�<,��:��n�_���)D="�q��qV���=�˰� �)=cm�D�˼�;=�����}N=�f@�y=�<�B	�T��bH=����O=�5P=��LI\��H4=�:=�K\�2�V�@���(��6���*=�#)�����MYM��==.Yz�W	�<�q����t��p�<�=��e�x�=	��޺�!�Q=��V�4���I =!�>]:���=�<���<��O��`9=5��;�8/�f��<��;��<@�<���<Ԅ=��C=��� [���M�y�g����<��=��ü�C���a}=G0V=8;V�5㼦'ټ<�λ�C��=�Ƽ ��~�c<�=�mǼC�ȼ��B�0=1^�����m�P�D��==��L�|̎<��P=3r���-��i'=lh���9��1�<��%=Z+��w$��5���Y�b�R=��<vhO��q�n`�<m:�����F=��!=)�����IGX��Vݺ��������.!�E[�<U3�ɨx<$A=�(R�_=��aY=�q�<�h|�k	N=\�V�%伜�%�I8�<��=v�E�--�@<���D6=��=E�D���W��s޻Ɉ�<0�<�:ƀ<�I����"��dh=x��<%�Y�ڍ���H��?���I=��/=p�<=�4l�
.��X{����L�5�J��ơQ<?��3+���m�=��<ؐ=��3=0Lg=pA��=367��6/=
wJ=�L/<l����<~v<�%�<
P��8e7�y�<��=N���4���ʽ������,��ZԼ=�"�j��Q�����]�K�ڼ!<=�q��ZM����
=K=	��<ރ�<6~_<�d��v��<��L�ѭ����8��=��;���8x�<�):��g"�����Iga;�gj�{B<��%�JD�G�
���_��=�22=��7=�V�|�[�B�D�=�^�0�=�$�;�Ҽlr]<d�;����F=�S�,B.��VQ=�n� ��<�
F</�u�$()<p����B=�q=��2�C�/=3��<6��n�8:JF�F*��V��u��<N=�*=]�y�Y��<�g'��m �y��;d�<�<
�9r�<�n�<(�<�#�͐S;�M�;�h������6���8@����<�L<��"=��~�[pG�=2�<
�����;+�=�4=���<)yb;W�W=�,��f�=�|���!<�fh=q�j=a�q=��� Fϼ����<�8�9�=Z�[;��h=��˹���<��7=~1=�0<t�g�f���-(=p�P=Y0�n�`�	*q==G=A��;��Q<�J=��(�/-���	=S�6�h��8_=��=$��M=��Ǽ��<V�\�'_Q=�Ż;���؄<֯��Ҡ���9�T?$=��T���;�,P����<]�F�z6���V�<�Dz=�=?��<��<�I	��\�]�j�ƻ�-�<���<�����K=؁z=6F��q.V��V��?�;�5����=�o=�^��Ө�������
�z�8���P=�%��R��<���K���y�<Gf
������`\=e#=M��<�=��<)0˺�N���$=,��<0L�XI
=ۭ�<� ��h�=%�T�Q"�<ӫ����@y<8��<ˈJ=��<�=�����
�B=�:���¹�m=��<+=Gļ�N9����;_b"=�k}����E�T<��]�=|Y
<r��;B=��=�:��d��d~�;��<�e�;��<DUF�Ƞ+:�H��6g�~��;�`<J�̼�&���G�K'��})�s�<%DS��f�г��r<'ې;ծ��Z���X[=C�"=
��v꛻_���,�B�='Yּ.=2�X��4=�D�w=�)��+e����f2�<zn<��m��@=M���������<-�2<�d�\(=��v<_һh�.=u�č<�VM=۷�<-�.;��a�C=/��<���;�X��A_N�M� �Л�<d&/=��	�A����=�<<�}{=�s�����<�w�����3�C��^w�=�<=��Z=��w=0?T�ln!�`0��]_�6!=5�<?�����;Ͼ��!=��;=_dļ�u�<�Fb=�(b��5�<���;�*ʼ&���jr�<y(�<�WF���=r��<�	����L��+=�
�<Nȼ��<����U�=sZ9:@�A=�k#�U}�;�l�o�i<���d� ��-W�=�f��c�����^=L��<8==��2=��%=x끼H�ļ���<��g=��r��Z<2�@��k(<$x׼ ���X*<ˉ_����>v?=C�<�=L�%�ռ�-�!i?��=�<��<����<�i�a@%�`
�<�C����~�<�;;�Z�<�N^P��F��Q���&p��򮼾��5qm��^;��<�f�=� ��C"=�~&�v`5<n]��s��q�:0T����9�:Ԟ=���<{�}=�3S�G��<\��<��<�dͼ3�_���	��/��D=.%���BP�%JI<�T��<��S_��l=����P������K�91n =���~��k���i��g�<�[X=��<х���h��Ԋ<>=�l�m=����
=¸.��^z������<��Z=1zK=Qz���L����y=�MW=�.=H�<e�*��I�R�F<�R%<�P�<��軿:K=�?���`Y��c={�0=	�|<���<�><��=��<?ٺ��8=�n=3��a#�4��<�ƽ<y�[���q���Һ���H��5�<O6��~l�-�D�'�]=F�$����;��<��=��0=B��aW;�@�.2(���,��b=B7=�w�7=�[n�� J=?ü��B<��=E�=@w�;�/���^�<$W*�$z�����5=1���R�V��<�2�<f�|<F�B��t��>�*>���~S�2t�;ɡ�<��=4v7��y#��Y<��ۼ�j%���&;��:<&�O�p�5�%@�����}�W=(� ��@<�\�
��ó)��CR=��/<���<���;��<��+=U�=��<�j�9p$=ך�9,;���k=��*='?������x,�2�<�%`�k��< �!��i-=z1��^����҉/����<�<=x��?�<F2��*�X��gO󼫉H=f:�# L��=��P=<	�<*�)=`�=�=W�G���Ӽ-�<�gD=�g="��<�co<jc⼬�=`֚���l�����9��<�珼��@��W0��"b<��=�,a=!=�Qb�E�Q=��,=�`�Mռ�Kb���|=���$Y����*��&:B���=�:�6i�<i=� �黥?��Q�2�w>=V�9��<���ZR]�vg%=	ܟ;�%�-��>=5$�����2��=i|�<�	E��~<Ou[���l��D��w=*�<�)��,�Y�<al���(�"�B�ܩ�/�<�v7=!Z=�~��D`-��T���3���'=o�:=Ԡ���ZA<�{�<H����ļj�����R��:,�G��=�?;=i�=2���^���#����<��}��Ϡ���v<I�޼/�<l�=~<^�|�^�dX-�O�M��g��^�;� h���i=-6=+�G=�_����<���9P�	u�<Zw�<�'<K*&�{1a�UIZ�i:r��U_���8<�o��V8�:���G�s��9��w"�<%r=�>�<��=r��\�e�<lQ�?qn��5��6�<)�=J=�-��:�U=t��w�i�a �;�z����!�c]�<\�5�<Z��w=t�B����ǧ=��2�sF-�^ԼM�h=�0��8��c�6�1��=��#=��ۼ�lR:�h,�����k�<|s1�H�����(=��O=��J���8=�=��<����似|�1�� I���?��A��Dx<=�<2J���N!�mļ�{9��䐼Br���j:`�J=o����<�V.�g��<-�Y��Pl=K5<�6Q�h�U= @=J�W��匼��v���z=)�<�t=�.�<��@;K��`'=F-a=�)s<����Y�=��<�|ټiڈ��7��A�"�.=�d=|��<��Q;7	���T�ܼ@2��e�<���i]=�=���`��=�H�<E$<Sm&=�(!=^�=P:����k�%����<̓;�HQ;,�C=Kln�y2�}�e�K�L=�s�<�j�5���>=��<W�@�י<�:��d��y!��w�+=[��<p�`=�$<g<��X=.K������N�Q�<8�=O�=��b��e=KBL��xQ���h�;K�<��b;�a�t��/U=:��<v�b��$�t�<��W=v��B�w=��V<��'�zJ<�D3�'p�}7�Kм��o(�:�O%=E�)=�?9= >U=@=��p=MKj=1�K=ۦ���MR�L^F�]��<d�d��;l^�:.�=J4�\�z7pN��ժ7=5��!S��=8={?'=9��< �m��D=X�L�G�����[&�$�^����<�R�<�-��)*�z<��<�O���ѻ�'���
$�}����;�'�<s�:'���C�<�q�Z):=�0�5�N�*��E�;�=���V@(�L��<cB=���<g�<iw��O���D�RgK������o=ON�<�2�qّ<_?�<��.=3	ռ�/>�����	�8= �=�!�<���e��p�!t��"���*=��>�M��X�ڼ�6U=7��<C�z=}�/=ҽ�<L}Y<���=L����������<����TԼ�޼��a�یq�G��<�,=H=P�f��@�(x<웾<�Ǽ��u=U��U��}�M=�Y<�;:=��>=L;�����}_=
�=��;����kt<.1.�<��;�*���*�<t�<X��q+=��J��c�����������&�����`���|=�V�=i���<~�t=�K]�k�=�>$�,Ҁ�C�U=���u�7��.�N�P=��e=��<�t����N�u=�ͼ�Ez=�x*��1�<�����<�k켇@���7�Ea?;�+1��H��؃<[-������7=o%ܼ4�.���8���<K?����<����=�n	<�N+�Y�=�:�[x�<����=�c�<κ;d��;k�n=ZT�<�V�<�	'<�f ��L�<�t=1N=x�̼7��h�;-Bk�"g���"�����>������<�8&<���8�<�b�T�G=���<l����;�k̻��;.�R�3}J�=�T�;a�=~�=�<ѭ&=ֈ;��<�H&�����J��w�<��i�sPu<�#='��	������m�����<J]%����(<mC><=^Q�<�%<�9ؼC �6�<��!�\1D=�n=,�b�<gc�V�;؟Q=f���A1);$��k���#�7�ԼpI��70�h>u=yR|<�";=.׮���V�T�	�=G=���������a��<-^�����H@=�t�Qm��4p8<$񤼄�7�m\O=��<La6�����r<p`��A��<���߯=���e��z+=�@����;VO=	=���SVj��x=+�;�Z �<�0�<&�<�)�<��8��g���r�P	:���A���;�1==���؈ϼ8^"��ռ�ͤ�?��<�P�4P=�	<u=k�!=��[�~/�:�|�<���<��=J�>�=';� �k�G=/X<>��=m��<�{�<x59<�;k4�=�A���żz��:�T=7�A�*��<̮�<;�k<�1�;�r�<�='@"��y	�Qk=2?����Z���뼎����żY����JL��= =A��V�=�.��8�<�=��I;�;��<�z;w>��A��W6��8=�u��#�S<�Y=�Fz;b@����<g/�<�d���
=>lL��^m<M�==�r=�U�U圼X��=�� �wh�O�<s = Sd<]�G=
��<~ڋ<��<���<E|�<LU$�:0=�������g�8<gp�<�B<ay�S�a=����^�	=�{
<K[=.�뼾o��u��:K�=�I=)�/����;]�L=��޼
�ں-�E=�i:�������G�Ӽɟ4=��<��Y=a�P��2= �W�T=���b���VF���Y��W�淋<�4̻-ͻ�ԛ���B�k��7�<���L��<����Kw;=5[���<N=��<2#=��(=<B=��<=�q���=*8�<��:U	кR;=��<4S�<�T����8��6=Аm��=��e�[�	�o��[C�|�p�5!N=��<�� ���f�Ͻ�)��;��5<>�S��4W�ƔJ��~���/�<�pQ�D:���Z�=�,j;������d�q��<#��<�a<=[����F��'[�d'5=%]��j�=1~<�ב<�޼�嗢������<�6U���`=T=_�@�D���4��>Q㻢�W�k��<N=H���<��N;�
�����A�<�_<�d	=���;`4=x��<?��I�0��vA��L<�?��5y=���<�=�Ȕ��F�<M�������J<��A�:�v����������T=cE�P�g<�6���X=�j�s�<Qg�F�����/���
��J�<���g���#=y&=��<P1�<|I-=0�ۼ7�;e+�6/a���}�U�.=< *=k��IpP�S\!���Z��pa�u\�+�ټ��=lnS����<'p<��+�����+G�<3>���7<ʼH�;��_=��*��{x�;⊼|ߞ��Yw=�/�;X�<�;ϼt�=a�<g=)=[�����<s�������-�;&=�5=:��Z+8����;�=�@G=_ =O'��3�{}4�"�=�W=~�%<����b��U-6=HC<�"��I_��$=s=�<�z<̖<H ��:=�ez�<rއ���h�(b�<��1��%���󆼏#d���k=��<�GF=�({;��=i��;��X=mK������R=�e=:~�%ȼ�//��V����8; �=��=>���|���+.J=���<����,�<�<<]q������p}=��;����<E��<��=z�7��bY���v��E=c����A����q!<9�E��L�#�z�z�|�gO��K��y����=�/(=F�л�l�<wܱ�'_��"==1��� ��	�K���W6<	.=J�9��W�<=�zF=�L&<��M���O�M��<�@O=�=y�˼��4=��=�Ȓ�u�-�́��,��[�Y��Q���G=)�]<��;�yY=�h�<��ɼx�:=2a�<u�<ݦ���%�<薐�aPP=�?c<�z=��]��T=�G=�����l=�E�<Y9�cJ�<��)<Qa	��_�;ٯ�<��}�{<F+ �rC�Լ�7�:2x#=����
=�M�����<����\F�~LA�/k�����ã�<[�,�p��:\�S<���;]=��<�%�;�-=]G/<��=V�=$�/�%�<��:�k=�ۼ����4t��� ��L¼��;���<�R=G���D=��Ǽ&�g	S�s{C=�:���˻�[��RM=K�'�V=����[���#=���<��=�@g���;T3��0P�u7�W�E��V�?i=�H�x�<B(�<��<�҆:����xH=R��<�w��\-^��a9(�g��.��	�U=���<<��;l����^�)�"@�<�9=x��=ִc=��<(W=j�:�P�g�<�=��P=�*�<��a������N�b������<��:���<ca=(+=F � \9=z�Q��u��=��^;��'�))=pL�X�3��LN=�~@��Y5=�<�R�<ݰ=
��� 1<~]o=`�=�p��@%�<N�=1�Y��`<H�<�T��x�;���<f 0=���<j��<kl:<B1�<?�����T.��a�=�V<s�X=J��+@A=�d=9.i��Ǽ������;[=��<�|ļ�	�<�4��3H�j"�g�<���<���\*�O�:<q@�<��<(ݼY�N=��3�7���Ǽ�'=�/�<��-+=C��7@��K��<{�̼u�<I0+��`<�f=oZ��c�<�G*=��S�f��<�e�j���N�<O!U=��a���J��*���/)�)�f�̎�8͞;u�<4Ȱ�����Gy<`t ��U���1x<R���DS��e�;�i�}�=t?�r`ܻS��*(c�ż�y�"�ȼ���75C=�0n=p+����ۼ":��M=� ���|I<������Y���=ZN���2�+�k=#t�@]�<H =a��m
�)���y߼()x�2�4���|9`�t������y;�I<�4\���Ǽ� H��?6�^Hw:<8=��1�+cd��Ț����┻�@�<���<!�G�C�O'+<�	�<��&�*�����<�h����`=ՙ]�q�=z�:��}<GN=�0'=�^U�ۯ�)y=�-�; 	�<�[b=�$��8�<�p<�<��f��I���Xt���S�G�0<TH���<`�r=��Y=3�K�=ڮ<�dZ=�S�e���=��B�;M97=��:S~=��=1��t����=���7(�׹����؍<#����Y1=W'��jn�<�� ;븰<��=P�<=��<�vn�7�<Y�<� �<(�u=O�A=A�H��==L����<�$
=T!=�UV��h<z�Kd=w2��ܻ�:<Jg�����<��>���<��9;{ş�>�i=�}�4�1;4�o=�1��q;�o��ƻ@�� <��i�;Tj;�&=9�	=X.�rHͼ;^a=t��<��;)8��+�;e�<)�7�ڗ�;��1=��=c�H=�_�<5�<1T-=�d<i�ݼ�)B�Xs<���:��;�V=�og<5����2���X/D�ݡ =b�i�$N^=rO����{=![{���l=s<���="����7=�S=)����:��=�
P=���<]�z�IS��IV����=s���^�<~KM=�����`t=�g��9=�3̻����wI=M�,=�0}=M =�d�;�$����=Y;�<G���<|м<����vi�O���M=�n��g9,��qH�+ �Y�R�� W<�����PQ�C47�51�HL=-�.=��0=�A=�E �;�K��=���C=��><����G�|<3`o�|;��+�0A(;ǚ[�o�d<}�����X��<�g<=�E��,<�(
���=O�>�g��<"x7=oÈ=G5ż���<�:<u���d=;��<�\�mb3=b�O<
x�<y�\�Ev���$���?=�v3��aH<<��<I�=�G1=�5=�:#��e|���;=�j���<�.!:N�ͻ��=�YѼ@0o�n@=��z<�_�9��m<�<=$�[����;�V(�������K�yRY<��B=2����\=���6�<	�G���<���w\�te<L8��YG=���=n�<�Q=[8=�B;=R��Wu���B�<6�/=^�J�z�W�-�M<(=1��ؠ�<��)�{��<"�=���<Wy���`[�<犽Q�'�u�`<�ϕ<�.�=��=���<<X���2�����<�z=t�6������&�5ݎ�%s�;{�n=�yS�mx
�mU<(Q�<�O��\�<2��<�����A�<���<�)��?�j�R=�P(��}t<�j�:9����O;��E<=׷�;��ؼ�g =�4�<�U�*�=�`?�Z�2<��\=��F���<��I�/`���-5��z�;�B=6D�ZL=�� �kT�z��;;ya����<�\ �[A�.��������X�Hq����)���=}&��TZ�<;�;|M=m��<�}�;Ҋ<B���,�E�����Zȼ`�K��#d�^?���/м��;By�Z(�/�Z�Y��<�R{�>ٜ���b=���<�ޱ���G=��B���<�4�<(D=�m=Oa��=T��<��G;2n��+�n��'߻�N0�HA�p��<#h���g=`.��h<�L=A�Z� W��k<=TǼ���;�G��>�;a*�<�(W=Z;��I�C��=��=�V:���!�ռ �G� �H��|�<��@���<3���TX�=�ݼ3�=�q�rS�<M:���S="J=;�O�	&I=����=�W�<D�¼��u��=  �:O=~�ἢ󪼱��=��t���<���<& �����=T�'�@ʡ;е�;�P{�rl6���"���弸�ɼ,S�;�	'=f�i=�<�W��;�D�h0ǻ�QN=�s���[�@��B�����F�'�ᮀ��bU=Z*3��]�<z�c<z����<��̼2�<��>�xѸ<��<�0��1��<V��w�������<�r=��<��"=�w��h+��eZ=�-i<zʝ�l:�<��^�/z?�Q�<��E=�'==P7+=,	S�ƚ�"0]�e�<��!=B"=s;��#���E�<�p:�ck��n����C<)��<�Hh������[�K��jwټ�R=�hF�Y5H�2�=ܮ3=�:=ӥ<�<���������R@�_�e<F�&���=�-�?�{��<�c��>��<�no<��=��:��:��H=G��<  5���������<8��<�M���s��q9<]:=-�ܼ��ɼ;��Q����Y=!���ϓ�� ;=��
<�r��a�c��{<,�=~���k�t����=��	=R(;��;=�=�<޽�<m�W<��=��G=�8S�5�<#�h;
�q�H���j-_��IO�n����<o��Bĕ<��=z�:�s��\��|��9�9�օ���~=d��;�w=��<?!�:˗�:�EѼ��<"���0%���P�lH���/��R=��t���<Ӗ���鍼�z}=n����j����k�л��<���:�<�N=���� <4�;�\c�<���.r=���<Ic��M���q���T�
� =2e�<�o��8��zJ�<�|<�iH��1�/�"=�/��Ղ=�˻`=��=��4�~�R=�s=U
���ZL=�$=ʑ=)=m=&E=z���a����f�=�=��:;�I"=�܅<��X��&ż|<~=eu��-=�m�;I1=���=G#�ڭ�<$<����,�R�v=�a=�3��g@=�L�7����4(=����=C��*=А�<*��;4�F�����6��A�S���<��O�R�<�
(=V�<P�r��XѼ0B=�a��r���=�<j�6=c�ڼ�1�<l?�=��:�=)=�\�;�rS=Co<�=�+�ф��R��x9���ļs!Q�9�B��/�<�=E��=�
��\��ܰ!��d���8�<�+^���]����<[=��AD���<g�ܼ�5<�C��m�N����༙-�H ��H� =�R=�5<��<,�ۼ��%=y�=�n���������DM������{2�%/��0=�弱[X��FQ=�u+=E�*��j�Xg?=y�J������S=#�	4��J&=�y�<N���vR<h�<�[�<����W=�6W==Q�<���<����G�ш�R�=k�o�u�*��/;����a�DU�;� ;�O_��s=$K&<�&�;�W ��p=��<?�L���<4��<H�`�~��;�R<�J��u=�v�;��o��E9��=��0�pJ�<1��<���=ܰ<�%�<�E=x���'m�%�h=��-<N�!=��H<PD�<^hv�b��k/s<R����;�"$���A=Lx�8�
��R�<3B�QF��J�=��T����<Db���"�#���1� m(<� '���P<�v�<+qn�r�0=��!=BL]��p�=
ㆺ�4I����<��^�W=��=�ӄ�Τ�;��C�F �%K�<�z"=n"K=�aC<g	޼1��<�6�<�%�t=,=Z�;�f�<�*G�D_Y=����G�q�<�*�;̉��X��v	�vA=���:�)P��y%=��1���d��<��u=�i�����;��:=�����:=1��<Ķ4���<�]�T`=�ot�eʛ<�4���=E��<�$=y������g�Ni���'L=~4׻y�J�=��;]�=�󼻺�|��W��f ����<��[=C�W=�
=d=�W�<�LB=L(�<׹<=��<�o3;'3�<] /��Ƽ�i=����λ�τ������po��N�=4Ff����<�¼򁽣�!;&b^<��s�)�:=�^B=a&�<	J=$M]=�!��`�T�뼫����9�[�d�=V�9=L���u����r�伄׺<�=Q�h=d�;��_��U=װ|=V�=Y�̻��|�����wp�p=�m��s귉�J=ټP�s�x<g�;l�=֭r�V�<�N��A�#ud<��<��<>U�������a<��N<�V9�1ɞ���;odY���<���<��t=Р#�ru�<	�=�g�|�����g�;��O�s���<.�%���=uq�<5I��0 8�Td6=�7^��P=(�����ʪ�3ռ/��<:���G'=��g=p��DѼ%�z=�����L�U ���^;]>�<+�"=�<�.,�u&(=rYU<;=!�B��Lh��1Ӽ�cS<����I>=zN�<DY�<M���7Y���1c� 8t��"N=,�����<���<��=���=Y:i=��/��:g=���;�2@�6�=�J�<߄[;��8=�h�<ۜ����<����	�=��X��<��=�9)�ot��q=+���*�<@`���=�)<J<��g��ӼeؼU��<4{(=ٻK<�8��H���X�A�-���;=�I{��$�.΁<2�����;�E<tK���#d<�h=S�U=zv>��d�=��L��;CN$�N{1��v{��4�����<~�)=����X)=��=�t><��`�Om#<�[=%*]����<[3<�!����<�����+��~�===��<CGp=�,�<��<o��<�)��H1Z����l<��<Y�e=E��<��Ƽ6Y��*���;v�<�J��aꃼ��ڼ%��; `B�w���!��<"yp�5���߻`�e������#=|�7<������W�c��hd=�z����W=��j={4�;�|�Vg�c��b�:�4%�ʙ5<'A}�͋;)�L=B�����U��2�����ּ֮����<����6��X|G=`���]d��Sv]=\*�7�=(�z����Ƽc�ؼf�]�`��[�<����M����+=T~!:{�N=ΰ��+���e;�`!�9u=�����ڊ:6| =5�;=�8��&<ڪ\<gxT=�q.=��9�b<�Ƽ9\B� �=�{���p�<���Q=_���u`=M�������}=R���$3��a�}�<=�"���V�<X-�<�c%�/<ߗT=�������s��Q&��b�<���<�U=k��98=m�B<p�Z��T�<vճ<?�U=e��<������ni=��d��nT<�5���y=�D;��û{�����0<�N���;�w��'�;}�P���m�L��<j���A�"	�<�&��&�Ji!�7y��?�,�����V�<
�bp��-<���34c�h�?=M�=Q���=J�?=�-�'��<~�Q=((�;{��0_u��)=v�	�5�<1֥�T�=�#���e����9���<�o{=���<	i@��w7����U��:Ƀ�h� =�Є<bpc<|�~�SQ=i�<��<2�=��	��q�ڼCB��eL�B:2�d߯;7rE�bR���=jp=�f<�u�<�S�<�"μ�I?=��'��f*=Jr�=~<Vo�<AO=�@�=y�=���<zd=S=�����ʂ<Y��<[��|�X=�=^\;��\=�u��e��b��� =��;���i=�̓=��
��a;<7+���W�T������Dc�:�,N�2��^b�<�.�<�s�<�#=-5�<����l�=��W=3�}=�E��rw�W��;&�=�V4���s���<D&=���0�>��� ;�|Ԝ<)�&�[(m��\�-�<���<�U󼇊��.�;R~R=����g���2\S��g���p��AI)=͋b�zd�j�3���t�`(<u\企�=`S =4�&='�E���F�/�.5=~H9=�>=��<n��<�au�B{3���=�$���$%��7�ʾ�Ч�K��<8!�\�G=à@=�4=^�%=G��=L=�D��J�< H <n��;�F��N= i<�zm���;��<=�{3<r��@�����ab`�P�<�;��Q��<�RI�]d_��~�<-��O�~�Nc_�C�<=ǜ�������;�u�F�?=x@ļAm"=�<{�ļ�9��i=���r+<�2@<c�g=����0=B�6�ת�;K(V�C�c="jV=�R��K$�������<�,�����o|Ѽ��R��d"<v\����<�z<�k4��UM=��?��=c4!=b�<���u1��XT��;�`��+H=J�N�a{6=�D�֊B�6�=B�ɼ
Ҽ�h<2��<r�=��y��8���������H��c=�-ټ*�=n�	��!��3E��~-=9A�;wO�<��8=�4=9:�;u|��߻��<e��Wf=#%Q=���<__�<�9�YA���<���O�v����l<|==n��ɜ%�$�p<ss��x���H�<���G=J��<b{.=2g��Z�����<�k<��<���b�<��t<�)=��<�!��_/=<���BA<�]<) �<`<��E=o�e=��g=|�<��<���:��s=��&=�wg<�U�"�=�d������"M=�K�<;:�:�?�8�,�V�U]U����:�=�vE=ʴ:�Ll;J7e=�I�;~�?�U|��T$�!ɼc�G��G�;�j=db=���@:p<T^�?V/��>��i�=���;�?�9ˆy��F=��|���V=zە�j�m�Z=�ٺ<�o&��j����z��q_<J�=0�2�ɾ==OLN=��X�:�����V��d(���F�00�;x@�<��<h#�����<3�(��+��@��b4��=v1�<�l��z�:=N��- �<b{=�<���&�畄<K`<<d����	={�:���(��Y+=I1=P��0�=Wqջ1�Y���@��<*����*?=�S=�d�<�������H��>L�<��5<~�R���=��B���������/����<��<��f��Zr�L!<�{"=�������=j�a�n��;@��Ŷ=;�5	=mzB�>�N?��<�ûg�d<�9n;�v�S���q�U2��jʻ��������!C�<Tȯ�upK<��Y�@I>�"~q�*<]3���;��B�Vz�<v#=��L���>=S�#���<,�*�g�c<�=:%k�<��»N�����:="�^��I���<?��;�e=_��6.=g%�;�o�/�?�3�2=��g���u���<�T�<׎�<�W=�.�M� �����;�"=d����	��z\=8�
=ɜ�:ă�<w�r��ۄ=����̈́��9�����8���
��d�׼ԝ(�puּ}�9ՍD=K=�q6��D/<�7;&0��G@��4�<)*&=��=�h)�ݜ��<�$�)��~T������<��6��=N�L�3�=����8M�sTT�Gpf={]F��N=��U�8�;�A�k�7�$�<k��;�౼���K�8=��#���;]�ɺ`��i=:�};���;e���y���g�üco�<E/��R����9�A�=�"ݼ�5�� �,�ɼ@��Vv)<t��A��4x&< bl=wA;�Ӭv�T��;��8=Z����y\�<!�Y�
�[<j��<C�=Rfe;�3\=����܁�)g�9��$<� =`y��>q�秼�=4(��2=�3@�eO;�����}Ѽ��%=4;Y=6��ؤ�<��=�~==x::�I�ʼHf�<�z�\�<��r�&�<�}q;=�v<ѿQ=o/=i3=�"8<��V;`���J9�=�#�.�E��dT�� <K��I���2�<�2=~��
�r<���;RcN�J1�<��::X7t� ����ͼ9x�s���ޱ<��$���=���y�\=�ݻC$e=wu�<�5�]R�����<��"=oJS��EK=~�޼N��<���}e=�L=���z�/��K�;���Oz�����k�Z=t�$��X�<Ps<�0���?����;�#��<\i�q|�$?<��:U;�<P�.:�0P�<�<�>=���$�Լ��;o�(=X�n=\%e=�l�����_�a���n���n=�R=g��A�1=!К<���Z=�ك��w�<����W=3�==�*5�6I=o|ܻzi�<�A=R��<f�h=�?��[o��u�&���э�<��S<o@'����;��<�:��{RA=��<�)�<�N\<�B;vM=x��<,�� �m=y���#�= +�9;��Q�n<s��;s�<G��< �I�ͪ�<М����O�+a�<��*=�I=������{����<�V�<�ا<I1=�!=��<g�享���J����=���<���B1=�K�� �E0׼1G=�j�/�c=�ӥ�L�T=��Լ˝ϼ.�:��P����<��8����4;V1+;�:���[=��X=|��<Q:	�СI<��Ѽ0�u<u����V<զ��I'=���<,σ8UE6�x ��0�<ʋ�Q_缕�=���;Iq��/K�<ǳO�eI�;w����C�mI���=�,λT4.�SB�<.��<�U!���<�-���5=8<bj?=\��<#B#=����w���ق2�O9�O��s�<\��<Y��<.g9=�>U=;1�;7k��K��o=�x;��u�\�(�٨�<��T=��G��4<��l��(�N�&��������<���f_=�4���M�#�<PT	��]��I-��c=WF��N�U<]E���8A=��<�3K<,L=��5=J=�n.=EZ2��#�<b����t�<���;���c�9��o=�����o��R��.@�!Qټ�x=af��W��:�Ǽp�G={a�
[I�l
���=?�+=S!"=��P=�7<�G�<e����9R=�ؚ;�����Rk����*��
���8�;�E=�G=�0[=j�%�1��qHʼ�Mռ�Z;�W��<ط����U�e@=��<$��<y��[��;Ij�<�kn<q��<���;M�x<�ƛ<���<�'=�?=rL�]F� �t�ɬ�<��:���<���:�B=d�<�һ�DP��u)��Zm�2�=A�=tf=T/=����d���F=8�&==�;q7<=��%=�D=� M��J= ���Q7��V�<
M��4m�<R���s=m�b��6�9�{�<qI	=K�ӼS�
��=����<a��<YR��M\=�E�����<��S=��Ӽ4�l=V��<M�O=�(�	(������=p�<��=�uC��IE��*�r����ح�/�<G�b=QP��,�߶[��S�Gt�<��]�fU�<2���+@x<���$�zA=��y��=����;=t��<�#=9�5�����&!�;h�~<	~����G���M<}��c�D=�9��%��ϼ�L?;45�78��0<8�<\_H�	J�<��A��9���&�K%�<+�U��:3=&�h�v��#�]=C��<��?;�=`��;�m���)U<!�<��3=.K�;v츻:���Pr	;��ȼ��=R�m=��J�q9<�y ��`�<�朼JW7=H��󴘻]c=��2�}�伇="�w=�P����,�=���T�����;��0=,(�=6�����<ƄE=�`ĺ�L=u�=%�d=��<~�p;�/w���K<�d��ꦼ]���'�-�~=B��<b�4=ѪL=4CY�ϋ�\$�$57:��<o{��&;}z=<N�;;�U<O��.�=�-�<#k8=��;�#�;^a=jeI<��p=���<�DR�2�k=E��<"�.=y猼ⶼs�ֹ��-�O�]���C���<RM?��e�<�a=i2�;�⾼rQ�QZ=	����P%���|<6�;�H`�Π�<8W��!O����(=A_=�+H�4J�Z�=�Y<;8��<8�+�������%=A!;=�g�{`|=@g=ԗ�<Z����'={�N�y��7=�W<��:d�<_b���6=��v��=Y؆��0Ѽb�E�4�a�F��<���=��;�؏��L�і꼹[�<Uy�<vQ�����+\92�<,s��+ڻu&v��h���y�;;ޓ���;K3<�����<["��x�*<��b�M6���%
�1&==��j;��P���ּ�(:�]�7=��[=T�	������%=��ѻ�L�	s�<N�i�<��,=:�^�'�X=�c�<�K�ú��,�u�5l=�c��2������<g*������1$�+���@��:�=�<�[W<)�<�=�po=�<�߃<�n:���[��>�ļ��C�"Ue��;�����G8=9�����;��;�X=�9���r=YT�<��=�����p<������x��<��g��=�K��!T�<O�}��A=I<��,=��X<��y�2�P=J*<;�ڼ�sM=蕼��=��^�{��� r<�I��|�<�놺��q����<(t=���<[P��*���=����>�7=�=�53<���<B��<~T���q�0|S<pN#�=ï=���ZM=)=6�拣��X=^�g=�󼸴|�� ;�X$��C�<���o=r�����Uf4<q	ǻ��M=��=c,���;׉=���<ʻ�h�`=��8=���<�<9�q�9/{=�FԼ,���x�DBz<q��'ƻ��-��`�;�,̼w;I=��U='�����<$f��_i=h�t�	�K=wo���R��U���8�޶�;�5Ի�OJ=s�r=O�B;�޺<��5�à=z���qz<V9�=�^ �P�<�d�<a�޼G<=��ź�W��!���R�y�U�����<�Ż��9�.l6=�8[<�60=��O=}v+=8� �)-==\�����4����8=F=�?j�O����C_��J<�F�<��<=�#�<�<=�耽6bּ0�5=�ы�yB��
�<E|=_��<�f��0�7=��=�~����<?E�<�<��V=e�F�¼�)�L�G=�:?��@Y��Ef���Լ,���w�<��q<baU��B<�N�;j�=�:=����W�C��I9��:���B��Ł�L=�<��I< ����<��S=m��r��F�4�6F��NXl=�VG��Ƽ��F=�(�\�2�z\G��i=fR[�b�8=�n���F��mH=��J=��ͻ��<Yݻ-�C<.x��|Vk<�:W=b]=��w=�R��gH=�a�<���<��=��ܼ֟Լ�uA=��$���=�9��t/=b��X�\='��<�G1�������<�x_���=u��8��=K=�	O=*���,^�<f���_�z_��1C���	=��ݼ�=��n=�\=w���C=��=�l/=`�9���Z�<q�B:4��;�&=_a=�V(w��,���=�c�����P�J=b�.��J=���<�f�`<�mY���c���D=�M=��9=�}�<`#�dT�>,=��==W���<�h�i� ="A�<�猽G{^�-�D;&�<�M.=��0�� J=X���뼫;/�S����7�<�qX�*Ŋ�p�=@��<j�=�"4��u=G?��9�<)�<4C;��\=�>�;͗�<8o�<�M_=>�=��.=�{c�@�W=�߉;y]i����`�;I�(�R�]�K����I�	��;A*�ڇe�M��"��:�&=uX���}=��+�+_$=�L~;�<=��P,껖c=n��<0Q����=���=f�,=�[;=9";��(�q�~<�m=T���4�M=����W[8�j��� ���e=�D%=B~��F=�b���;����ƼMV=y�=�80���9=�*K=&���� =f��μ{?m�YG2�T�<e�)=���;s�<3ӕ<2�==�������N�&��:�r��� =�X=J���L�:�g8=��^ D����`q���ʼ���1=U�<�E=�]<w���N==^4��^�@=<@%���<V֓<V���\&=22�O�;=�;�9R�<>�]�݁���N=W*�<}X=���<$�<��?�gμx�/=V��h6;���<�IV=B62��1��:jӼoM<3$`;i�#=h��t�G=�c�<�L=��==���:�,�D=؎B��(q����;&��<��-<�G�<��=�.=��p�}��<W�<_)<�؏;�/�<�k���-=�E��l�;��<�nB��c�<#p�B��<8�8�4׺��,�,y��n��W=O�L��P=`��}�>=���<��1=gB�<���<�/1��������<g�l��HM=s��ԓ��~���\S=��=w�=r4���e;��<�r<{@=^';3�F=��E���D��'=5;ͼ���(m��]�<�7=�&=��9��49=}Fo=!P��g� ^<<oK��#7<���<�P�cj���e%�vv=9��<��s=E��<k�F<C6`=�?��Ž"<��T�4���-��u�p<��4������E�p���=��#�#c;���6��%���	i=��|��C<�=���<����+�<HC�[���V
�: ���?+U=���d�Q���f<
 d=	K)=Y��<����<�<=הF�m�ܼ�u';`�q���=��<����4'"=C�<ȝ���$�<k��;������y����:�r�w���*:V=��^�n�e����_v&=!hK�D%9<�<�<�o:;!$=�Ng=� ���������Z<a��y	='�G=��U���<z�$=�����<+З�<�=(*�;[��0P��1`=Ϳ�<�%������E�_��<F�<Z�=����ZzP=@ �����6�;<���<I��'Pk�k�.=S][�E�=i5=87���g�0��>�;ʁ= v��wt�g� =��P<&�:��6=��=䃖< �ܼS5���<�Գ;E<�:4�2�~T �Z�R<�P;��#�8i�;w6�;mJ��C=vi޺t8Y����;�ׇ<�y��X�������S�-��J�[7���=�=���V3Z=��X=�������or;�P�μYv3�yR)��;�<b�E=^X=tI�p�`=4y�<�GF<��=��Z;D�q�=nO�������<=<��ȣS=24���P;@�0<�+��CR=V8�]�a;Pm0�zr��	�,�I��:	��;==�?��WN�<��B�2_==��2;4�L�sc=�z=��0=M�<��K<�?<¾<�a=�4�<Q
}�k�&�~�:���Voּf� �Ǌd�N=*H�<)�	�S�5=���<�׉��;�C�a�`�է�	�<���<ˤ���:�$�=�M�<Ө�m�<�_;%gT���?==���0{=�ԗ<(�1=��<�B)=�`=0�c<��<U,��j� �=�s�1rY�Ȑ�;���<�н����?eA�V0}<�Ư<��<OA4=Td=/�,���i<��<դ���&�<�/�=E�D;I��M�=�'=�W�;��3���\�:���'��}�<��@���<m����x���=u��<6� =��¼N"=�%<�`�<4�V��d}��q�����x� ��(��p=�l��먼~�<#;�;��z�^q�<�J^��H=���]��"=�ǿ<5�=%s�:9b(���8��x�o|���-=�����q�<�P=��v���%=�"B=�@=j`=�F�������E�x�H=csS��+�<��B�����t=zs=f6o�c�+���B=�S���<(�f=8���!=�=�)=Y?��Q=aH<�����G����;�;��b=\f`�h�O=�<1�=\�<\�T=�B8�PƼT\=��?�2���kd�ˬX<�n����a��<!����O���Й����<�J��.R ���}��5=�W��9�/T=*��2��;4lN�~ԻP3��	3:H嵺.�`=���0�7=j�g=���;���;k�="HȺo�<�����?}<�E��[&�<DxU<4�< ]A=z�=A��_M(��Q=A����T�K�:���7��  ټ\L5=��4=��<�LO}�Bd��d��=^�2=0��r<8��\�����	�g=����>�<j:��<��=��:=�� ���<�F�<�-=(��;r²���<�,�g����:��R=#A=��=��<��[�L�Z=p
�<Y�<E����Gx��()�O]S�����<⚼� �<`NN=>�;MA$���Y���_��:'�<&��	�;��X�A��=�Q伱b=6ۻϕ=��^<�Z'=���<~�Y�,
Y=���n��<��:Y��<e�-�&�s����9�1E���n���8��=���<��e�n��;nx��֭Z�7;���:�<�;G"a;�j���(<� ��m)=s�E��>�<ѼA=䝢<�b�� �N={3�;�E�^�ռ��0�|rػ�lF<��=�켒�@=[��xma��$n�^�^;�RD=��=��<��;9r�<�3|=![�v�Y<3�#�y�����@=#�P=�3ļ��E=S��:2��<��U�$��
�;�G7<���<���<��l<���<��hF��b\���.�؜ֺ�yj=S#=~�$<����f&<������<[�:=�	<�Ħ�$o�;���<'[C=3ͼ|A ��_{=Z �;�����`5��H=�=�e��o<���<.45=�O��� ��R���=��N=�==]^"=dV=��.���@����<�Cd=��A=��#�@��;� ��b=z�\=KX�<	�k=��p;֠<��==8$b�%3<��*қ�����?]����'��K����;5Sż�J=�	��[L=F�ͼ�tR��n�;�;�;�Vw=�m��]�����;h8<��?�����3�e��',��;��3��u�;
+��ɰ;�����M��qɼl���s�|����jd=c�H=ej��_�c�3��<� n��h3|�di���V=(k<R�,<��=9=�3D<��<�~��,˼]-��g�/����<k7m���<*�g= � <��(=E�M�S���<������<n���z<�G��,@��B�;!L;���.=����̼�������:⌻팎�����#L������P����-<=�CI;��}���%=cD�<�7;F趼&���=_8����<��4=��.��z\=��<�m=�Xv<�!3����(=��:����.��F<�=�5��%8�<�=�<�m��3=���LO<̒�<�<{�<��==p����,=�MI�-V�A~%���M=�F=�o���[E=����J�b=��(�[����&��U;]U
�*̼m.��A#���Q;�-���!�_�<�����
��v�;����M>=r���o=%:=,pn=2j�<Y�>=Vl����/=�93=yB���1�"��<jz�<�H���A=�A��=da<��ü_%��q�<~2�E ��Fi<����+�� O��oU�]�麘�>��ڴ<��_=\���Hp� xP<+8'�Ba���O�<�9=="=μ�V<ZF�<�ͼ�v����9�x�<�q���]�X��<�Ң�ɤV=!�=�<��h<���`f=�k���"���9��X=�Y��<��<��:�W�<?� =�`z���"�C�;n�;�%����<�7��>m=Xv-�TX�=c�:=?�<F��<f3ļ�=�ϱ<=��Y=B"һ;�D��\=��~=�dU=�˼%�[����b�Y=�-<hD�I^�np�;p%�90�<!+ =u�j���<{�<�ȟ�B�*�i=�K���>��r�
2�<�����۴�:��7tS���;8�<,.�;�g���t������m���/���{�;�9<a��*�<�iy��+}N�Mzf����<%&��e�<�}8=IAͼc��<������-N�ı�<\�#�B<=�l;��
=W<N� 4=<?!�;�n�<���;�ǲ���j= LE���<��<cջ���<#�P=�o-=G�D<B�Z<u�<��r����<�}Z9ͣ�s[��S�)<�;�� =���;��
=���� ��G=)R^=��<6ol��\G�K��/QC�$L��_@4�6�2;�'� = S=,��<�!\��ن<�Y�e%<�2�� �<�?����gey<ۘ<��(��~ٯ;Ǵ;��H=v�%��_�=g�e���6=�Vi��k��B^�<0�4=��I��$���=�k���ػ�M��T�B=Z>=:;S�[��<���ll���dN<mN<x!=�6�<df=� �Tr�;i��<�-O=��W=�$$���\\;��ݻ=�d��<wă=�<������-q��;#=W_;kA�<��>��\ɼ[=̻��+=Q4=�ޅ�<�Q=�>�;�S�<XW��B�8��8=,<�᭼_��i�F�<9�E���3S�[$:�i�:�%O��Zv<U=�(����l=�O< r���<O�L�6��;h-{=��U=j�]���߻½�=z<�<6=]����r����x���.E=0���D�/���?=z6��.�S�<����T�X� �c0R��">�pD'<�g�\[X<�]�K�0=�Ja��kL�0�;$;�=<=̨��9��gK?=i��;�����<�=X<>��<��(=��<s�-=�*=��<�y�<�=8�<.��9������+<6�$��6H��0;�Z
�H9�<�F��C�<�=~=�@%��g�w�N=G*ͼ��e��?�
�I��k
<�=S�D=���6)����b;SS+���T=V��<ok�A�==14=�!C��N=�{�;�(�<�+�<ʄ1��`M�(�4���;{=��B��m�<�mM=��ͺ�f
=|K���r�?�=�j�<*�=���L=K��:�4	��F=c�?��
A�
q�<�T<�X�9��V�I���������;��5�I=�XKw<7��<#�Ǽ�=Kv=Nxټ�|.�?~�<#�������j�;��K��{/�b��:�q�/	<�E�&�T=;�=�Uy=�s��	E<1�=�U�����:��]=A���;��*=�;�<���|[�ڳ�<9FB<�X\=PaP���=,A;W#='�<#ԣ<��4=��<)M��ԼQDT=�Eu:aH =�扺p�0���¼?Iμ�=�Jzֹ!J�<?��/���^�C<�I=#�<��J<4M=V2���U=)�=R�=�o�;(�t<\		==�^�V�=U�=��N���ӟü�fC=�Z��`bl�ۥ�<p�=7e&��>�;R*��ϱ;�a==B><�\�t.i���;�=)#���?�8(*�$�����:���]��<���E�����y0<A���� ��+�3�K�9ʼgql<!fr<��w��3�3�Y����њ<ǵ��,=��� Z�<�Xn=@�==5�I��I,��=��Z��g=t��<��i�5F�< �"���<.��<����O <M&F92�=�9���E�<B_/��U��=�����<��I=Y?�;�<ȣ�<�N��!=�����D�<=S�+��<�<
�[�U�<�H�<�\<�Ñ=��=�s��L��B�a).��} =��<=Dk��#�:�ħ�;�6�<�`�<M��K�<���<��Z=�����$���M���t<B��/"�<��<�<]��F�<�z������H�2=l��+e=�1<�<(TF;�{˼�ޤ<*'=O&��c)=�;�<��<\	<��?=أ�-k
�Q�2���Z���<X�;��}�e=?��<5ۼ,B�;S<��u��,ͼ�5r�h�׼��>�RWf�ւe=�iͻ�{��?B�s���ZW��'-=�t�<�]�_MN�^������;@�7=�a��L�v`�|����/H= (=���qg���P<���<nK=�3�<-�>=s޼ ����<nU�����BY���?��=����;�=2=���<���N=��(�~ON;�q+<Ř.<=�漧���K��3�^*;ZDe<�?�>g�;V,=���*��=�=�[%�u��<�('��Xx=K�Q=���<���>��sn�������4$�,>M�+�Y��RҺ�����=Ƕ����<�v�<�kD=���I4�;yPu��=1=/80��ȸ<�(�;&#)��aC�TC���B=��u=��-�P�#=���<���<+�b=;0�+J=J�
���$=����~�;�bd�K�=�:�λq��;�N�%��t�9�2=���<�b<~=9=E=S�<�f�<ɼ����-���5	�<MD�<�32�{�;C<�k�<�nN�\�=u��<R+m=�<�"���V���t~����<mn�;r�/�wE�K"���;�;��N�<�C8�WVj�v3���C�^�1=�H�ϴ�<�d=���U�'=����Fd,����ۿ���A�'�����7��d.���~���|�4��<_4��=����<�W8�U�V=o�<�B��O���Ż�[�<�}#���,��1�<~�y�X��o8��Sz=a5ༀ�t���z��^9�!6X:d�`�Ӽ�;=4x��v�M=#�;Q~����&�#�=C�T=�$u<v�o=���<Z��<9����$7�[R���a ��B�F��<M��'Q�Z[=�Kػ���ĒI���=�="=�O�<y�:=�޼
=�������lz� �e=*yU=d�j�_���u�β�;q'!=9�D<'��<Iv=ku=D�Kf=��:��C��Y�K=v�$��81=�=]=�`/�ͭ�q�����)���Ļ�4���Z�O�<e�����weX=��u�=� �㱏90�=<W�@�Ѝ��=�ָ���<���<T��<'�]<�U��L)��<=��5:��<�	�=�ߎ�-�����<^{�n/I=���0^�d���<��[�Κ�<s��<����я�=��Y�.�J=
�V����<�lx�Ʈ�=}7�����
�X=f�ϼ��+=��S=%z=ůǼt<t��|�����S�9�]a���q;l�s=�~�<��H=���<�D��KS$�	��<�f�µf=�8��/R��Լ�ټ^���n�U���]�pu$��jȼ��Թ��[<�F��p�B���I�ʎ)=�*\��iA��˼�񡺨/<n޹��%	��'��:5�Ts�<5�`��'�IaF��bN=�Uh���#����<�"���<3�?�'�)<*Ψ�'DS��$=����Z� �CA�;I�O��b8����<s@n���J��u=�s��S��(��<��)��Ԥ��z=R��<R#��FQ=>a"==�Ǽ�N�<o�w=�RU�qU�s4��y�<�{	<̿�; ̼]ȝ;����_=�|u�����+\�'v��s?���QʼCz�s(��K=r%��3���P=��=F9=2�L�_g��2b�%A�=��8�m�!=ؾ߼��]��'<��r<����$�"���z=}*)��O����<�Cp�FY��ܛ���=���<�E=��i=�l���k��L';c�;�{=��U�o� �N=Wǳ�q��<O�R���B �:~�=�'X��U�<�ڥ���S��)�<4w<Y�1�<�ݼ'�=d/���R*�Ql=�[0��Uռ���<C[p=6������>�;n��y��=� ��D�<^px=�)<�*��/<����,I���<B��W����?�[<�%@�ؗp�u<==ܼB����1�<J'A��F@���T��Y�<���<5��<�rȼ��4=8z=���ޮ&=|E&<j��<EZO�O�j���Y���j=����/!=�IE=P��{@=e}�b��<���<����OC���<�=�D;&�\<:�=�5=��U=危���a=�a����պ�;�<�P�<ڳ�;�M=d�8=�U=��i=�N=�[;GT=����<�*=�5��e��Ub:trR=HR��y�]��ɐ<_7A=�m<��=V��<quF=қ�V&�m4��� =��<Qj��l���i2=.ff��9��~�<:�U�V�R�K=v�Z<�����3<������<pXX=Кa�.��;!NL�������Y�k��<�N���KY�L��<h��<6�����`������=x<��E=*���Nl?�e��<k�';���<���cE���=_S���ƻ���uw�<P�D=���<����D�o��<Z�;H:��s�T�Pڼ_6�<�v���Uh�JB6=������=II�5��<�n�</�0�-k��B{�"��}c=�#i�f�m�(��<��<y0غ��A<���<��;=ɹ�<��g=�$D��,N<b�B=P�t�^�3���<���eA:W;�kϼ8��j�X�(H�:�zn:ݢI��3��D�jK����T=�?m���t<3�2���%<]�Z��R�<~����"�\��.e�<���y�=�P"�H��{I߼�4м�Y=B�y�H=�u�Ԭ�<r�);ܱS��~F��+��<=�)�n�7;���Un;$�e� ;��J=�eR=�A��4�_d�;�"1�?�m;�=�=4����
�šμ�
���G=z�t<���Q6=��A�ᶌ�˽�<��$��P����ļBE=Uo;\e��[�ڼ5D�=�JK=��";��2<'J=wX��D=���<	؄<��=�-=����84=��[<�E���3:�WW��<;h��)��T,���F=*�N=��b<R���c�U<���;�#�cNO�*����v<$]$=�Ȧ<<�����]��<`Ǉ=�S�=f�s=Q^��Ǽ�.�a=Y�����;kVC;�ϼV����	=��C<
���DR�<�� �IƟ<�V���!=�^=JC]�t»�B����<�X�T���!A��j<1=h+T��򼇹�]����\����<�fY�6^Z=�" �kn�<Խ=���<�,��T|�(76�&�=b�]�4���<��[<`���	���)�t����<
�g<1Z;��;��L=�(Ӽ��Ƽvu�;�9�h���%��<��<��û6�2<Y���:W��W-�5�^�5h��m���ˊ���q�s�� s=���KgJ=ї����=�0����<l@D=^�0=�'=�ŉ�6xj=�.�7<"�:�W=�E���L��}�=��>�Y==���<�4<e�)�NS=�I=���<-<?�=�c�<��B= v<V��;u ;�{�Cn4<�([=�x��֑�T~�P��<Ij
= �l�E=�ha=[��<X�_���I���=���<ֈ<��������'��t]����T�[)�<���;'ε������x=�"��8�<u�t<�9g=��=�+�i_�<C���<(�;_�����=�$��,��;�X�����pNP=Qh���,='��;
�<����-g<����F�����C����)=aK�<���<\��1��:_��<e�9=�X<������;;�:<D�=a� ��hK�����V؃��g������Y��[�<O�w<\/q���c���7�r��vͼN��<a���.
�:��=����<ъ)=�>�:���<��=9s��G�P=��<���<��;1����D�����>���;؈<3����C=��<=�N�;�Le� �=]a{��0��}м�'�����u1��1Ȣ�O�M�u� <\�<�=�����W�p5�:0@�G��;#i,��W����¼��;[�1��?��A�<L9��#0=$=6�'q��>�� =t:��T�K���%<�-=(�"��b(�J�;��A��M�A�Z=����4��$ۼ��|�bZ�<�����sG�i,�ة�<����H�y��<%]�<�t���ǖ���= B0=n�#�9�&���<�'=�S��_Ӽ���9C��<�.=�>�w��<�5ռ��+��M�<#ɴ<np���[����+�*m��S������;'���[6� ��<�wK<�.=�ǘ�=�0p���&=�⃼�i<!�=X�+���,=��9}.��D<|��<E�#��[�7=�0]��	����&=���%m?��U<z��<�w�6�<�D|��*V=\��:"Ha��q#<�dʼ@q4<''��[ļ^mP=��C=�'O=+�V�L@2�'�#=h�(<٘}���7�!�=��/=L �<|���GS`��R����=͉� �:cBH=�y=�3-��X� �f<�t��Ez�<��	=�$�;5�;��=���8�A��N.:e�\�Y@���=�D���j=�G�\�j=>15����<Io꺡j�<���<��<K�=�v�<�u=G�<�P��ۃ�'��<�F׺tɁ=oR�WD�<���5�}�_�dZ��M�<���<�}m��S��+3�<���A"�GĎ=G=A��;�B�<�Ll���<���<G�<���@@R����<c=(�<4��==)�=�`=�;�
��M���c�<��	�޶���b=,�p<�x�]s�+2�h�=�)��i;�iW=]�$_��M޼��8�I
1�_�<	�L�2�-�!<U�*:��f<�3�<�|H�헸�'2Q�*༝q{<��<+�9��E����=�W�<�4=T�����:�~��S=��*=;�мKoi�vx�<^=���<�u�ƙ-�>�=Y�^G0=���;��(=�=�7<��T��M���.=�d(�4v�<�p���<&�f��4&��0�<��û��/��;n��<��r=KcƼ=?i��L*�<���<�2B���<tI='�_�v��'��d����������<�������<)˺<Hj�;���:a]��o[<z�=f��<:�d=QA><�)�<��<��=�s@=����<2�켘/����E@���=P�B=�<���<I )=}&��U��@r���<������<�ǻ޷�<�x���%�ː
��M^:.&P�p�<����=K�U=R�6�����7:,��=U���U�<i�<>r ��x`�T}�;����=��,�L��~&#=���(s(�ӈK=��¼|Yz=p� �����ؙ=�a��x���!����-[=u�A��ں&����b��k<s���ͼ�v;=p%����<g���X��l)ּǟ��B=�9��m�<5�L�-�޼�"�<rpl�����[`���M���x=ىV�-��234<Pe7�����5�=�u=���<���>B=�Z�<���/�<���<iM^�1ĥ��,d�uڹu{G�"�l���1k�<���'����,;i{�P�;�
w�?1�<�Z�<�
L�Vc7��4����O�nI=I�=㧅����<�XL�\,H<�<=-:G=��i;c,b�e�B=�3=7�#+�<I��:B9�������<��ϻȼ�s=�v�����U7<T�]=�bH�ȁ���G�^�Jo%<�Ԫ<��<Y�=�$���d=�z��'��:�;�8'=�?w	<�ͼo߻<�>(=�{i<S{1=*3�i��ۘK<O��=&��X�<��==�=�O~�܇<��3��HG��U=$���F�b���6a�ew�
�I<ʍǼ���;�D=j����J��b��z>���=Y5���M<�䐽��ȼSy���ͼ���=�!�::�f�<�.�(Q��mi;��.���ú�<�{|�j�n=�9=d���}:��A=�V.=�(R=} B=�KF=��/�Τ�r^=Ї�<��=��<��<.��<���<%5F��'�zf<��&==:�;N�漦l����<=��<6�[=�=��A����5j�E+w;W`=����D�<�<k��ő��lk�Ź8��"�� �3�ڄ�=hڼ��j�P|/���ż��=;?�Z<�g+�V�n==�S����=Tx<i���iL��N=�-B=��@=&�>���!��e�<C=\���D"=˒��LK�SXn<�;��4�Oj
��>6��k�;l�N�����*0�杚��#1=fu���u<�L=9fZ�v,�u�D��]*� rO<�f�<��?;5=~,����2�J1���J���a%����<g�@�u��Ѽe�z����;ہ��%�B�)G=�RA���=�2��'�i�k�J=���<$�s;&Z%<O��<R�t;�j�:P]K=g���vi��+^=�*�<��g;�>S=[/=����m�/=*�7=t� ���<���E�6=]�;ZX�;{�q=��-��z�M�<n�8=�"ʼ�oD�vA =^�=�q��%���j�<}]�����5<5�;��N=7�
m_;�><�զ���]=������ݻ��L�J9�<d���M���f=-��<#��=�|�<\����\P<��s=-'�<h��O�"�a-J=yH�<IA8=B$����m1*=8�u��U:;��=F�=3}J=/�=�������2��P<r��Yp�<k�x�MB=h=a�<���ckּ k[=��Ƽ|)s� �I��+=�s-�kQ��8�<V̨��X!=�<~������=h���X��a�<摞��o�;�>�<�ü���;4@<Z��p/�<f׼v�%=�ce���=a�����1��6��R���)=��8=�I�� ��;�X���G��tݼ_;&��aM=[{=Y��:b�#<�v���3��	!=�H����7��6<��D��1�+6=@gͼ��*=̆]=T8μ
n��bC��3}&=V��<�A=�R"=��4��쌼k2�<Vad=�y8=����l=%�^<MO<}[Z�`��o˳���<�9=���TB=�gu��Tʺ�R���f�<�-�=4�:=wT<:1���B9��K�<~w=��m�{ԩ;Sم<`믻�}=�'�<P�<�j<�=��\�p���#�<eռF���no��ἥhO=�ջ\���D	=�!X��E<�1��?��aJ���	�2��ռB�<�z~=nޯ���<�=H8U�{�!�������</����sq=J��<��R�K(��UO^�֫���Xq=.EL����<�<=���1���f�<��-;c�5�_�=�撼����Y�E���8ڼ�'@�9��&�̼���<��=�H����Լ�u�<��7;�X3��}��!��<:X�<���<V^ü�%=�}���޼?�"<֛�<�/ʼ6.:�� =����ۊ�q���Y�<�VT�<
��Tn���;����w�<�è<��*=��޼�!%�q��<���lv���<u:��W�<��)�vď���f��0=��j<or,=ͧb�`1�1cx=b�[=�Ȓ;5�T=�Cq��\�,�����Ƽë�9�л�fg�s�<��<�i�<��v:1`��-
�<)j%=$�|;=�:<h��%v�j�u����<��V�� I=UNR<�u��	�\�zJw��=�6N�d�K��t��'e=��c=�BϻE�-;��� Z@�|�?��GD=_�1��F;�)h=���`K�t�{<��I=ѐ=Ӓ�Ąϻ�x;���;���<Ҧt=�#<��,����46��'6=Tq�<���<lJw=�����[��K�;%�O��=��=	��<���e�w�8`¼��d���_i=H+W�E��gz�<����CH�*�m��F�<@���ڻf<����A�=�<��t���*<���y�5���<c�b=ꍽ�p&�/�!��9T=W%��!=�t;�!Y!��DP��tS���=�dp��Y]=ڷ3���T��H.=��߼%!�;��E=7%Ѽd�=���=�׼)�Fs=�z-��������<�`���J�=2==�4����q�G�7��t�<Ju�9Nr+<�����,4(����+��;ɠ:bX>�)�=_�ۼ���������<-��;�_=�L�=��< �/= ?=�a�<P���4���	�c���(<Ӳ�]e[=@.������!����<���Mw���0<�u���0=Sd��L�6��<�:$�C'��sU=��X:%�<�h���;%f���/=q��8|C��aR=��<�c~;�T�<<��C�u&1�/�� d�8ܩ��kQ=Q�̼�]����=JF�<�`�������;$���FL=���US����>�|�O�}� ��[;�)6�z�O=~��B=�6���� ���1����<S�P=�1p��\����ټC.)=��=��m�s�W�fW��ﱻ����<�ż��B=:���1�y���W=��6=��ϼ�x9����<��'=��^<P���¯�<C��<�]�<�ו�~ΰ<��5��'L��5�=�q=���<a�<@뻼 n\<���C\��f��vһӠf<g+=�Nj<�
=��	��RO=W㑼j����m�_�V=rw=8�����Dd=.�u����=b��<�4'=�֊;
����k:)��<��,=��g��d����<�(��'��4�=�go���L<�-�d����!�3Oļ��g=��V=1�~� ��;qa=�(�O�==���o��<��B=�|���=a�w=�!�<���y�6=�ߋ� ���Wi�5��<��=PjZ��,2��"=a����Y<�(��4�;��Ǽ*��0�6<d�=�QE��	�;��J�H]=pyx�f���M�< �R+�<B�o�@l�`�6=ފ��'��	�:�N}��W<(��z�g�ď�<�xx=v6������i�i�'����<�p ��^{�4��=�0���6=H,=�\"<#Zg���N��S�����Ș�<l~����<�%��xi��~(���f�Lм,=�\<�f���g=%��:�`�<�Y�*���|<��+=��p��ӹ�^�oܴ�G��A<�n�<UE�<g�&�y�<�F\=���=O�»Y��ߪ�	�¼�	=�_=|�;"��� ����:�s�ǻ"�����<R�:pT�;g�:/}3�9���E��;|�������V�P�<�!��=�Z[�=H����=�A�;� ����B=+����t�3S�wQ����u<��#=T5p�ހ�<����ۧ;�N�A������<����)=���<�QE=�e�!G�ХA<5�<ث!���<�w =�H%=!l�<�,<&3����=�2���<���W�.��-=��l�l���<M����;ŅP��]@�E\u�#z[��Q���4�<0|dz=Bh��<�b��tRC:�$=e��<�4<��{��P:�j���Y����У���c�,
=C�c���r<'E=\���A<�'�<�xe��`������iT���zD:�~=��'��t��jZ�#� =��W�.��"����*<2�;�C�%�=�8���t��=��\�ˀJ���D=����LY==rZ=��]��������w_=�^�"���<�-y�&�$��P<�r`;�d�<-,=��<<4����0��#��\�/;6�f=�82�E�;�DT�b<2:�UJN��3�^my�������<��1��ZN=���l)��@�<l]?=�'A=�A�{F�A�D2�<֞=�~���
=
�V<g���_�<$Q�<�F�<��߼���/���M�83��.o���|�����<*�;T�*����U]=\��s��<�B=�O�<��<=�=M�@�'=�0D���	=�c8�Cs��R?;u=�4f</[�_f�<���<|DX=�a�hų<{^�<9�\�QS=��/���z��ӟ���M=�0����a>G� .<�b'����<N��E�)��Y�<j�<V�=��ổ��<:�����jV��UV="d�����8�<��U=��;k�f�'�=:��{��<I���@j<��U��X�6b���ؼ��<��<Q���|<U":=)��<׵� [V�M�ʼ�2=�`��cx=c�4���+=E��=�+=������<'�i=l�<>BM����;C7=rJ��*����S<�rg7=�@|<�0=x� �ӲM=�`=n�<)�h���=���D9�<���ry�;�-=wF�7=Vȫ<8=�}Y=/=�7�<>�=��[�˽A=A� ��;<Ë�� �W?=XX=	�)=��?�n���6=�h���R�j��._w�{��<�9�1�����0�Ɇv=�<���\�.=❊�]db��z��p<��Iy�FpH==��c=`l��U��<�^M=� ��w���F�x�ټ~m=f<:=��;��K��;W=�P�p�=�/��pℽ���<��c;U���<��n="6�(=�[�<z�N�v+b�xԭ��c����<� �Ͱ�<�U����+N�?�8<�<�ʋ<A�[�<�	�W�7=kݸ<�D�<	t��X��� �<I�[�˄X=[8�<�^�<�6�<�O��T=\=�<�A�x	�W�>=�����l�g3<G"�;J�^��?�ei!<�$��:�H=���<\ռf�Y��:��v�O�;=u�_��zR���R<�({<��=˼��o=d�o�8<%=�Fo<{vV��c����=�t��#Z�;��E=��z���?�;M�<��=%����Y=y�t���X��{5��üKߣ�W�=��>��,���m�( �<]���>�����G<>=�a=�TM�s6���F;�+Y�r�=�('=$
j�df9=�޹$�<�F;����_���X�(�ܼ���=̟�2��� �<U�<l�F=Z�8<��ڼ˰�;���<�֪;)*=]nH=}y��<��=�5=dLl��Ƥ�@�����ۼ<�b��}��ld=�Mr<��=k�8����bk=�qc�6��D\=��=<�ȉ<��K��I�;���<ˋ�<�h=���;H�G=����.w������MF�`oW<�)���:I=���<2��:�bѻ$�U=��1����;���;7.�>E�����b�<�(7�Q�)���<I�A��=Xպ<z����:j=�F��5^���粻M�1���.���;v�;�x=�����ۼ�ƅ<�l�<��=��=��Y��{�<K�t��['=H)=&tK<:"�Qһ]�T�<�B:ᒚ�v�!�c9:���
=�v=��2�P���HK<�E<��%=��
=֙;t�;�Jjj��J�� �'�_=�|��o]�<�z<���
�>a,�D�=~H=*`a<�8�<��N=� �<h�*��=~ ���=g�$�?���H=@7<b�b<��<�!I�H�<�=�c��<έ	=�d����;���<��<=ӶT=(i=��<,�<��1�l�<�6�;��=�<ԸF=��|�hSP<<�<�-=��'�ǻ���I=/G�=���8x���'�9� =����:$=eY���0��gq=b=��@a</�=$�5<Q,��uQ�����O:=j曼l���<��H=n�9�c`<St��)��-��<(����H<�	#�io:��)�v�����N�<�h.=u=��q����ɽ.=�E
���ޘ1���;<=<Qռ[*T��i�<�c���#���L^=jJ��T�)<�C:=�_��Df�<����s�t=F;�;
;�����=.f������>=
�<z����a=��U=�
3=�YV<���<ϓ����J=x{}����<���<�9἗HE=l|Q��U��Ĥ��#h��2`��Ax����c�;��={�;��:�ݖ<b<��Q�=\S<����Y%��OD=�ߔ�߿u�	C=΁�9�={��4&���8=V]J� �`�;W������м�"=>�=k�Y=��<�N6<hH)�\�Yм��<��.�#U=�������T�?��ص<�Aݺ��<�(=�W;9����a<�[��\염��'��<��d��+���=WI�T��{��%�<*
B=P��;�pL=�\=/�x=ԑ���[��ߜ=�T�=�>��\+����"=�+F<�<B=p��;r�K=�ѳ<EV�﵂���&<0�<�\��iN(�h�:��#i5�6�y�L�B���悼,�຾���~�����_=�D �;}�<��񸜎9� =�$A��B=��[=�ޑ���A��@������_�<���<E"��yG��H�;1X�;����kW��� %=�]C��GZ=?=ؼ�z �܅< w#�Cƥ;{�ͼ���<l�ļ�[���N[<�[���	=�I=m8�;N0 ;�ws��-�u�M=J�U��@=��=n��<�.J=�^�;ᾥ��/=���;�<=������Ӽ��e=�u�;e{�1�&<�q�a�W����<
�;;Be=��D<�w;��S�h;���<�n=�ד<�P[<@�`�����]����<Ua���u��o<=VL.=��t=KN=J��<��]=uL�;��ܼ��b=2�_=ꐝ�.�=�U�|R�h���8C�̚	=�(�1���Z=P�M��{ =�p|�$�%��s*=��YW=�Տ;��Z�kJ=�_n� �<�������P=PO=�4�5�v�]=��Ia=)�_��O��-��]B�<	8�Y��<��=�N�<͌�ɖL=�_1���+�`m�[2=֙�±
<ls$���<Ι:�*$=��E<Xfj=�1߼0��<I<-���So];]�U=�c�����<9�=g�2=�}=�7�;;s8��<��<<7�����k8�ّ�<�!=�h�m{�����8�Q�M�K��s�;�\���)=�6<�w���<�?= �Լx�=�z�:��=n��:z��<D�<�ǡ���A=Q�'��\��Qcg�)sм�ɛ<d�=�	M=M��r�/=�fH��8��.T=���;�|09��)<ySy���<��<խ�3�s��ѼJ��<��<s��{��r�=�$2a�-� =ܼ�<xU��h���1=V|����<��l=N�Ƽ�'_��J�A�O��h������"=ߐ���T<���<u7r<>��k <�Ӑ<wA�q��<P�,=ڎ<�\=0m�Y�b=�F�<j����)���һ��(=�ǃ��p=��;��@=�[�P���b=ܰ=�AK���;�s=|�:��i=��R������;���<�7��C�\�W2)<�]�;�sf�:<=��=��:��=�a��&=!��=�7��ß��"�$�C<�a��C�"<M�<�=�\@����<���<�+=�F=�.1:j��<�O2�*�A�mi�0���E�5E#�q��-S�<h�$=�|2���¼��Yo�����<�R�<�A[���7=
�	��]=�<��<֦�ؑF=�ݓ<�{=k4=�߼<�����0(=joU�{��;�l��d=j��ט�;7�S�=�=�~��JD=�O�=�V���c=y9ʼ����I�==�e<{AW<ƮS=�R��k=�=�J=�')�<�	�R	��~[�<�0V�<�?T=cm�<���<#��;������	=���<K�6��`X�
��<��=3� =0#�,r)��/9Ax�;IRr���O���;�Xx=V�<H���?���<�\#=@_�=m��g�Ǽ���=a�+=��p=�@=�;Q�o0��<ot=H�=�p�<�}^�d�6=�ܻZ*!=R�<S4G=�qu��-����=�V�A�t�v�&=B�,�Q��5[��Z����j���(�<��L��e��h���;�j=��d��43�j�p<\�`�����0<Ȇ=����m�D=	�:�Rð<:�2=%�<W���R�f��0=~(a�an8�]m�<D$m;��s���<��޼�]*=�2����<�rc��=Ҽ�r4=��>���[���<�^A;.���p)i=S�4���G<��=�e��(���EB=�b=u�!=����<�[= ����hؼ�B;�Ҽ����G	=k�;�k=�<JX6��~�p_!��^��v=<�����*��f(=F�+<ȇ�;� ��͐��C�3
=���h���F��m==}�<�(
=������<�$n=��ؼG�R�t��<B�f�ޛ�<]�;s�G��;�j��<o�~<�V��i���	��r�;J����`=Ł�����`}���=�r��FL<��3=�sn���F=��)��2��dѭ<&1�<�+y����<p���w=ly�T�Z�"�<%�*�0#�}�J�����.;�v
���c=�@�k.��+M9��5��:V��7�=���k =~=��!�����(���=`��@;��f�<��|=�Z���<z�R��J-=Y��<�摼Dn;g)�ɼ�����z;_
<���Պ0=`�V��=�9{=1�;q�M���=�ܴ;��[�>���:���=� �<�6=�����R$�;$<-/�<��;� ���<�,�<u�<�<,���x��<�;�<��N=Q}F<uO<ݧ�;�
�:3��=��k�&�v�%1�����N�;@�;��ɼ�<�tX����<�Zj���OK�M�A;����B�;����k��.f/��[=�ó;T��<�K=�(*��X-=�X��+��K���z=#0u�p�)�����1�߼D�(�ü�lց����<�K���<+g�<?W�;e�����;<Oȼ)�<T�j��L�;�����Q�<�����[��a�v̹���;̰4=1.f=I���i�<��2=:}��d���U�<J��<3�x=s�<B���#�hO��*Z%=b�;��N�o�9=�<1�*=?���=b�����k��	����<�Z�C��<Ǜ�:?}��`����';�R!�%JF�C,f���&;A����h<"+b<�^E�i�4=��[=�p9��#S=�8;��+=vԋ�C�,T	=3��:��<f�Ż�9=�oS�!gE��/�<��Y=-Y����;���<t4=��Xy��G�<�K+�J"=Lo6��}1��O�=�r�;��=yH���T=�7_�|�);�����j&��l�<ȳټ�|5�p"�<=�L�6F���~8=��W����~$���<���<�Ƽ��<�<F=��һ�z���߼Ox�<��f;p��;�Bf<��<��p���<��~��T=^�<�=X�{=&ڼ��.<qS=�,�;�ԼUZt�쿼�s�\=<�=,�R��=:`Z=fQ⻳>=��E<�h=�bc=�hw�7:�;yJ0�懇<�1��8��<׮=t/^�*S=����T��t���T���)=3�<w���V�<�\�;G9R=�^����<#�O<\�<�3 ��f�<�%�Tu}�hUʻ���9�;�鼈1;�5-"�_��FJ%=���<��W����<쬻<$!n<���<��=&1�O�&<��J����;=�I���55=�[�<�J?=���;�<R�;�,Jl�)/(��X���]r=p�C�' ���!u�9=vF6�����޿��R�;�>[=/]ȼ,��������t���h=w���7ؼ��=_�$�"�(<2�g=03=�2&��l=r��u���W�;�aS<m�?��ȼ�r��i�=(���T��j=L�����A=I�h�%ɧ<��5��=[��zS=��ʼ�A���d<�D<(�=�d=�'2=��3�p��=Y�&=i����Mh���=J����^�Gr='�Z=�����D�铙=�=9E=6�.=s����ㇽ��c<�=�X��ż3���&�<mO#=$�0�GS�;[U=r�-��K��46��V�
�J�!=I3(����<Xղ<�m��	m��"9�J;�W=Qq���=��ؔM�3V�<�4K���.�
=q��<t�f<	z����&�۝��6�4�#=� �<g�ǼY�;L?��D{<�)M=�O�<��nV޼�!=�'D�nm��A�=�\�SBy�K+��d=߭�<M�=+<��ҿ�<��<U:2�	*Z����<��6���&=��=ƞ໧0�<+��<2��<�v#��6�U���#P=%����vݻ3�6=��<1=T� ;6���<�;1��j2��Kǻ6^?�wg�5��;sv<���:2�<�;�02;5�}�� �Nb:��C$��",=���X]==���<�J�<�����y=lme=҂�s=?���<=�g{=�:�}�<=�zT�+'�<p��<~�;�m3�<��-���!<p��<�y=�#G=���,*=�	P=ǨH���u=�
�?�<��J<K�K=ݜ=y@=7T��6�;�+p�	Rq=k�`�{/=�`�)�Y=�d=˫e��?S��'�<H�1��tc�[B;�C�<=P�<}��U�Z=���W?=��N�4yr��SM���C<6��<�A=�d�#�U=Y$�R<W���>:U��<�==ZN������c������U�ר<��<�S=�Ǟ���;���<�X=�(�r�+<o٫<� �;b�:=��^��ʼ�=n�S�&�^��9,�n��<�s���/N=l1 =�=�<	�$�^_;��kw��V��R==��&��C|�o¤<���;1��;O	m<i�)���;�F&��!��g7;���r��/�4m�<P��x�:��Kg:����D8���5=\_g<1i9=���Asw<f�f�U�Ƽ��c�S~���4���@|��;��<�D�<I����	���S='���d��K)=��f�	�;V�^��1==�����[�%�^=�z%=a���#�F=��A����$<s�a�A��e<��O�f2=���Ğ�<E=w� ����<˫H��Qs���=.����Z��Y �����<tpw�s�C�����4=�+#<~:=�<��e1=(�^�^!�;�\���+�����<"�"��|ԼUw	=�����<��dA<��I�~��;���9�P=.j¹�}G��Uy<���;�7=�R���v���S��GB<�ĳ�d]��!l=z��R(�<ׁ�<������&�8�PZ��xS=v׾����<��$=ʀ4=���<�?8��>=��<���<ǶZ�|)<�{���=1=k�+��"K��{*<u�k<��o=�'?�4==�a�<�ܾ<F=�j�<4<���%U=�O���<.1Q�֮����ۼ]x4��k�<�YH����+��<N:=,�$="%�<��=*�=ќ��F�=���<�/G=ZoZ�c�P����;��,��^
=�94��c=�?���=y��<�0=}mм/Vm9�+Q����<x��<L�<���"=z��<��</=@�=3�j<�?�<�kw=�Ɍ��L=��q���T=�6=����k<�Ph�<P_::v���P��A<ke�q�K�b�ѻK�0=)}P=�%=C.!=�2=i�<�g[���@=q�0�6?���H=d83=X�]��T��n��<��J=EC�<ZF�<Р���S=p�<�1:�#�����C��<�~k���0��[=�ϰ<.�=�.�<��v�B��4��QZ=�+F�&�R=$i��i��Ok���?=�i=�Ց#=[D�:2=��^�b�=�ż�����=65�<.�G�16<�x
;/=M��<n"�<[�=!�`��wW�e�m=8ߔ�O��<��	=�JI<�_<��m=$�n�[�{=HX��t�#�2��;_�=a>=�'?=���<�c��	v�<uX=��<[b�;�U6=(�b�"�6�B�< Gm<<�l�矼[�==v�;��Q�p<H��<�ۼ<��?� �B����=�o�<��P=JN�t�=��.�^L�;y�D��$=�/Mk����<�(���I�U�:�����=�{�J5j=/X'�1�7��;�� G<a�<>z+<�nc��H%���C�ָ��q��0���\;%^�����ǡ��c�w�.�
b<=� ܼ܌�<��=V-P��Ҽ��<�r#� $N�]�R<@U��n�ݻ�T/�oG0��߀;�<{n�:����m�*X��,&����V�@����d=�C=�=�M <� J�b��<�y�<������8�x��-Y�;靸<��\=jJ,=RK=���<���F껼ɩ�}������p�j<X���|�k<H֨���<�8q=�M_�����'z<6�y��b��k=�>=(���?���	�ԼT��{=2�<�F�<�F�<1[e�Ό�+�ڹ�{��Ӽ�\=|=��W���<j^`=�P\��][=�.���ͺ�4ϻ�wg����<�Pg�0��<��<iu�:��9=9X�;],;�[�E�+%��ٻ��A��:[�;v�\=�n7=��#�+�)��J�W�.�)�J��P��,0�<��D<-�':��=�&=��;Y~!=�i�}p�*�v<���<ɚ��O�<�E��̒<4���VAz;{[�<#+)=��ļG�<���<ҍ==L��<�滏�=�S�G���D�=-�@��]��"=J=@�ƪL����=��(� �B=�&��M�=D�S��;�G)��rR�6L"�D'=S:,�Pד��i��ϲk�/�� �V=���B}��כ<n"�?=�<��$<5��<�"<=˼�+���M���(=�<����c����?���ۼ	.!=�0�<�J��<Oa��P�=��J��ꀻ��;�_h�{�/�-�D�R�=}^c�U�w<2(Y���_=����f=��<�AM=˖=qZ���V: V=����G[�cq��2<f���! J=2]H=�):=��)��;�:l��\=7��<D�H��-�v��<@ =�{���נ.�������<���i�%�l�%��ǎ�ŀ�;4�;����o#�<�K=DJ��z�n����K�J�dW�=b?� #<罀���<#�=VM¼���<�nh�|=�fC<���:���!0�"D2��~��dH��"=C~��S=rC-�h<�4;4c�<0d��x��<b��<�	�<��-=�<�o��"�:����<��Z�F=�ͼ1~�<�f���=Qě<�C=]>���4E=ڜ\���-=k/=)
��P�%�������Ӽ��$��WE=��=�'�F�h=�u=��1�^�ۼs=��<b\g�_F�<[���ߗ<k��gr_�T�	<"�����<gy<���8��q�<��D<��Լ�m)�U�H<��`=�!4��X�����w	伹���.e�<)�=�&�@<��8ˍA=1�,��	=ҽ㼉έ<f��������"N�mHH=br���ȼ�Z�:�?_<�4==�c�<�y��`
>=�"�z��$�ͻ��\�\�&�$�<�����ҋn�Y9�<��=�=��d��; ';�>V<�n=KO���׼�X��]/=�l)����<.�*�!�_=��d=`�`=��c=#8��p�I;('���R�k=�&-=X{f<r�= �9�䨥<˙o� �g�g���SC9��m���=qs�<��;���=� 3�k�H�P�	��,�<ӣ�<I�M� =���l�<��߻!�����<(�=
�M�f�;%Õ<![��7ȑ�._]=t[Z�O�+�;�I=�s��V��r�,m�<�m��N�T���=|]�֥;R҉<� ?<��m���=�BR�	Y��<�л���� =(��>X�]�B=�2���s�<]�@�{�J=���q�<���FY���`�<���@�����4�(l뻧�����%=��3=�N�u�i�=F���lB�n���=�	�\[M=/�ջ�=<q�0=s��<�Vd=�-4=d�>=���k;=X��,ݞ<Z'��Q#ϼo���
=>M���=��u ��	�ؼ�;l=��o<+}�{5Լ��	<�_��'�
�h����<�M.���=H�ߺ��м�n,=�K�<�4�<$d=�hR:�D����r_=�[�`=Ȣ�z�5=j�<��b=/��	KǼ8�=M�A�H����b�==<�<�=X���t�:�<��8�%�T�n������<_V�<�Z=�<8=�D�Q:��<g�<(�=`rR<��8=2���r��;�CX�(p�<ez^���껵z*��O����9:L��<_96��S2��8�<E�!=�Q��Db)�?j=�@���<��)=�Ey<S��;��W�m�_;�n<{�[=ǡ;(�=[�
����~��<��,��Q���K==�CQ<AS�;�� <��h�[�.���W=9�|<O�=����}��<<�v�q'��4lּJ�3����=��e;��t��z����<��g=r�)= ߇;�#�<��<�X�<�;>�"A�Hy�<�u�<�@
=��H=�kC=�=�<��[��$�;�S�����< EB=7�+=�3��#=<��`=����(�R�=�g"��bü�~=��+��"&=�}�;���Qta��B�<Z2�\j=lQ <�lm�=�L��K=P� �۔S=��ǻ�#������|f=�ZP=͌/=R��<Pi�:�U=���<-?j<�!���(=,G��0xx=��:	�D��́<����H�ʘ����"<���V@=Ȉ=*��<��2<�Y���<��i=�fY���ʼ���g*��ԣ���><�a<j�n>";�HS��;�߭�3=-[<9耼�?=ϲ?��c�tV=�5<qK:��$�L�`�m�H���=�����v=���<�O��͏��c�����<�!�+����#������_��ԏr=_]���kD�~�A��O�<ZV�{�Y=�r$�6�<��u��|#=L�Y<j�9=ݨ���A���=~$<�K��9�V"=M�>=N���ͼ�i=��̼(ܮ�-�<8�<��<��¼��[�.�l�=�kżM�=��y���st<d��Zd;P�=b@�<l�<��	��=&��T='��A�X=oq�=�_���O=�4=�Pj=�<Ho0=4�<0`O=gp@=��v�sI-�8��c�;{�A�;�G�=�*4U�mh���ֻ5{�xD�6��B��;J�8=��K�P�[���=d�3�Hm=&��<���ך�AK2=������h�6F[�Y�z=E�<�EB=A�+�F�<���<� ���l"���?�G��=��$���d==G�}O ���X=<b=��M<�N!=��,<�#Ѽ��=�p,�`=D0[<'4�_�d�P�9=+Y#=ؖ����%����<�e<��=�c<}CL=+�?<:Vn=��5=�=,��9}}b=Ek=c��;�(I=��X���><�\e�tA���<�A|=˄�<$E�<��=��kȼ'z<�<q}<����^E-��<D~=�ļ]�2���<-C=*C�<�?j���;�{_=�:���%=�9�����<O�=�F2��=����~�5`R<O$=/x=k�<�8�:��SD� �O=􄶼H�뼱���3����6��=4F=W*<S~�rf8=ga=�<��/=��3=��h�l�.=S�������mi=�|#�JP@=�l�<r��<�`���:=�과,?3=[���!O�*�:V*�;:T�� ���	=��&#3=T݂<��9��Q<�A>��?=DX ;���:<Y~��� <1�(���2���j��^ɼ��=��=���<a�e��]����F�Z�ż�-�<V�f=xZ7���\<����MaF= �q<�(+�j���AH�\�@��%<zE�<9}}��3�|���=���;6��<�~ֻOx=�,�<��O=R�8<Z�N�� ׻��:��2���M=p�0= �o<���<��+=)��9���EE��/�<W���Fc=1ϳ�����aE6=?!"�<��3=%S�<}��<s����e�)�����6~��y�<_Wż��;� ���=鏁<���<��<E�*=�S=��*�gj#���N�}J�D��=�/�<f�ʺ����=�rZ�sQ����<���:g=A�9=֩�<�0��λ\Y=��A��<�ȭ<�`t=�n�9d���>�\�)�$=��h:M$;$n;�>�<p4:����9�32=��L=��
;�G=|^��Vo��~6��OK=������<,�l�X	=bWߺl��<:&<:��<�W+<rK�\&=O���/ȼ��b;�9<�P=��<�EH��/=HaQ=�L.=����=�fg=<`����=�z�<��G=ۧT��:k:��0��$�<H悽������J=�uټ,����3H�JNܼPbY��.�;���+��=3=�ٻ�w��,`<9��<uO;PS����<��h�	�ꕨ�]�*�2�ּ���6@�# 8<�S=2c+��� ;�}=9T�@�3<�<E�3=��D;>C(������<<��f=
K�;=�λF�6��ɼ2+��J�e/��ۓ:��;M�/=�<����ټ�?<� ,�g"0�Q��ݼ?=~8׼"�<8O���#F=��=��-=IR&=��F�/��<�L�<"]W�ˢT�j�=z`�<��1<ǿ�sO>=i_���0�*ﱼ �)�7�ּ�j5=��ݼ�S�<�&%���"�5����0�]�=��j�QSg�+�<��=�?j���[=yC=g�Ѽ�ƺ��*���E=ۭ��T�l=#��;Q�Y=���<�<I=Ѻ�>��h��y�������~=��ջ���!��/�%���l=T�;��-��ŽV�H�<`h���s	=�M=͙K��Ҿ<�����!���d��-=�)=�kO�Vx= �L�4׻H��<t�׼M�d��,9h���2u=�0=Zǈ�%;��~�E�TJE<���:�K��Kɼ��?=�_A<�b[���)�)�J=���=\��z ��v=>�\=�<��p��
�*#�v��̎�<�M�=�E:=c��
��;�0����= =O;��P=/T6=�v=�lK=�o��P�W��w(=��Ep�:8%���8<U�2��/����:�@��9��N<�*����<�ҡ;��<��$=��b=C�<,=,�=]ۻ�����K=���S�J<��}��Q伐�=צU��u<:2�;��*=M���ɷ<��f=R='�<���<��/�����=1��\n�J�����;�����s=�2=y���aԼ��	<38��;�����b=�-�a<"�=<SǾ<��d�N��-Q=t���=Q9�]_�+֯<���<���s =��-=9S��e^<���ܱ�<Ԙü}bT� �?9�3=��
U����<js<�<��'8�󊳺�@B=�p�<�!=t��<=�<�Y�< �<w*l�ϊ�+��:Fd-=i����A�<Yk=]����՝:�|h=tl�<�A��̅=�{=4��� ?"�z�<t����HJ=�5�<E�-�f�]=5�m�#_x=�	�ѳ:<�+=z�=A@f<O���Oݫ<�y=v�<���<�J�)��<b�L=��X=�*�<n��<�g�<5*�<o���|����;�z�c�<t!-=���<���<ݰJ=�7<7���-�==��	�-!ϼ��K=�g(=:��<S�I��3~���<"={�g��A�<��Z=�mD��io=���\�=^ʛ�Q�����b<�t?=�Q�<�x/=���cP�<�3=Y�E=�X=�'��	t�<�f�<�u���N�;L�;~�b�5��!1F�S�5=���;�ݼ>�&=�V=z�;1=�o뫺���Z�<���<Q�=͢�<�ŷ;ڃͻH ɼ�S;)�=}D�2rN�ֆ=m+=K�3�`�"=+�8=��ܼ��7t~8=d@K��}$=_=!��<gi^�O1%��<���u��%=ÂT<A�=���<Pb�c�j�A�)�����	vZ��!u�]=<H����P=Vtt=
�*<2�<G�=.�R=�a<>O�)*�;F��<��L��v3=�R/;ڔ�=���;rX|�s�&�ݵ;t�O=��1�&��<�T����=;)�[��D��<@u�<}^��4X�O�F=�x����
x����O��C$=q~w�-��<�`a�5j=��@=��l=�FU=�=���̃�<�������=��K=�m���} ��"k��6a�n�K�-`�����7$�r��9��J�+�K����<�쇽�
�<�p�q')<���=S�+�������=aB���<��@���d=R�� =|�}��h;�vx;U��<�ϒ<�j�=�\X����Z�M=�'<��=���2\���D��:X"=����H��;aC=s	0���T�-��<]���hO����k���л�����<���<�U�<"(�YSP=9D)����:�{w�eC�{oL=���<>6@=��=�"=o���r�Ѽ�Z��o엽ؠ���9��"��O�<}=�H��`����pY�j�o�Ҥ=R����<�)U��B�<�)=�S��)��N����	뼓�g<W���/s<�B�<]H�
q;8Z=�C4<A5V�)����lv�<1C����t�==�=��<�.����w�QDE�ܾM=�E�UB���</Z�7�Ƽ$��gq=�_μEd�< B�<{H~=�TH�k�8���=��D�)5=)�B<�5>;�k�<��I-׼�#N=j� �T=�44�n&<�~��=��H:����2c=`=��=��<���eAF�n��;��ۼ�������>N�<�dJ�*.*=��$=�)=Z4X<N� �/=�R=�������H�<^�^���'�������q���#�o���Q_:�*�<SN<��X�9="�� SE�{�G<���<�Fo�5�=�/�<R5H=��<��q�8=�ZN�S����� ��CC�Zl�<�T/��u��3�'I黗>@<[��<S�ؼ� T�ę�K=����ؗ�S������F�:<PVj��5=g�$���Y��ƼoT#�!'�0b��X=�;�\=9�=�u�*= ���=M)h<�=H�+���J=o[�<��d<���<�=J�wH&�ϗ/=���<�[�q?ͼ+^�<A�f=o�Լ��0���������<�3�����
����'!o<��@�����ݼ�9=(�7�ۄm=�	�<3Fv=�$Z<M��� 6 =�<���<�gD=�����P����<⊊�X�݋�ǀ���(��=a�D��P�<[��;��&=���:@=��]��a�<�@Q��M��6=$��<�|n��H��-T=�3
�B��<�"�<dj|���"=��8ʻB��,}�<���<Y��<Ih���5�!�7=J3i�
G���O���U=H�<�?0����<8l���f=��<���z=tz(�������I��<����� g�I[,=6
�P���)�e<�Y,=Os&<���<����� ��'�6[��p���~�>�<�H�;���<Z&�G�����
��0���<��<"'=�+=��{<�]�or�<VmQ=q�7�%�<� ���(�2	L<�1�|��<�qJ�m_L=*��bT<%��<u#�:�p�;6���lm��;#�}�Z��uv=r�� ����4���;'�Y�p+�<��x<3H'�T��v=� ���2=�¨<h =rҰ<��<l
��]="y/=�l���m����!<f$��y<�<m:�<��N���=�=S��<�A�Klk��`*=5b=d�T=�.���R�=����-���V6|�]"]�kt���R=;���Xm=��=V_(=��
���K�t��`;��f�O�M9:�<�HZ�L
����Y��Ϯ<Zh���2���s<>j?�%r)=s����=�<�=M ?�.g�j�=B��9��8��=�5�� U����
�==k*:=�_=h#!���#����<��<��u�ғ_=�<��GX!=P�ռ�=�?�<�c�<C{�;�==>x��ϭ<�&a=��;Q�l;�I̻X�H�g���q>��Հ���|=��<�'��a4<|3?��=<B�R��&�'�+=j�=ʵ�9*�s����< �W<M��)z���=Ԛ�:�߰��q����;U`�_E>���[;�ڧ<�=�~'=D � �,�Ė�;�忼O�D���;�2M=�	`���Y�')<��.8�<N�Y9�U�������f<ь�9�WU=������=;2��	{���i�D}\<��=�ky;����Z=������;����j;��Ļр�C��:�i��弤�Y���U=�K=����5:�[�Q�=�v=�G�����8�0�����X?��H�<W/e��;��F=�b=���OS��Kp=헼V={�R_P���X;�QV<�߼��?<�끻D<?İ<=NL����'�&h='n2=�GA=��4�1@�;�%F=��;'��<Rd2�
H���=ʰ�<ߏ:<���ID���Rw�U��<�R)=��<~������;_�y���==��~=�ۘ<o��<eXU=���<&� �z)�<P�L=�e*�|=���:��=ð�;P�=�H-��낉�:j]=D�Ҽ�	D=k)���ɼ��j����<5F=�o��q".=�pV<��8��w	��d<�@�<
���R��R�<�]I=Z�3=O�==��ƺ�~+�����p�<:�Y��B�<5����e"<��d��?'=�9d=0�.�:�.=��<u��<�پ���V����<����̟�����Q@ۼ�� =�»Xc���&=6�&=�)7���o={'��:�"<�VȺk� =�UJ=�b�<���J=*S<��v�Y{Q���8��Ӕ<.���"f���?<��$��G����<�%=}�G� ��<lrh<K�/=��=�Zv=:�=�Z���W=Vn�#�����n�b
=B�"�Zz��b�<5�������b���"d�����zR=*��<�}.��aY�����BR=Y�����?���,=1 ̼�(�<�Q;���	=��#i��FW��g�����	��G<a�4���=c[�<��:(؃;]��<wἜ��<�i=t�?<��?��
���<�5�������B=�\�<aI&���׼ᦺ<<S�<\�<K,�<zH�<�⼉/��C=�eb���޼zj��{���<���;��j���K��EX�v+�d�Ƽ7*	=`<Hc�;�=���6:D)�`#=�U��pP�;��<#����e����n�<I���1���=y�<��=�-=��@=��.�{��<7�:zJ���7���J;\:b��zo��*<��d:��W�=Q=�	�</�|:�� =Zh=*W=.ls�s�=�]<�;=4W#�nR<�~=�1==GH];wm=y�4=���<��ּ�=�:y=��(=�[�l:{=��������3=RK=�m
=���r+Q��^��3Zʼ�ZV�dL)<�~�<Tv�<ѐ�|�8=����*�=܆�<���<�-��)��<�n���ڻ�p�<�
��;@���z�<gʅ:��X��*��C���1=&r��
��<�= Od<�@����<l��U>�HRͼ��i6=�7=��<�D4��:<��s91�l=���<�v$�\ �<�=�n��� =!�o;Rl;��= ~'��8$=��;��<;|�<*�.=w�4=8������<~	h=���<�<��=��׼INh��X'�vr���１냽��<��ϼx]��XQ="1n��{�<uYQ�Ӄs<�1<��a�&;�7*=G���G=Ⱦ(�Ά�<��8�����/��.=RC�<�==�$/=߳A=G4���=�g�0r�<h�@=va��g�����F��^9���p=BJ�c1A��N=N�/�j�����r{����<-�
<'e0�݋��$�.����<4�?��8d=f��<:7��?%=��N=
�e;T�5�51�=��Z=� ���z=�,�<[�;��<qc&=�T=H��<#��<�Ԃ; ;Z���<	O3=�j��Ε�,ԋ<������7�<�X=tIW=3a�$A'=��1��#=���r!b�=�z=n=��:�A�O���}<��+�h<*Ψ�|Z��R?��Fa�ck ���3�G#�<6ޭ���Լ6=��bh=Z�V=�58=�>c��@R�c �<�wG�M/�<�E/=А)�o�'=}�94�%���=���m���k=#2B���<P�q��7�8q�<�z�<���<C*��0O���R��mټ����#=%E3��#=�����=ׂ=�.ټ��#�]�C�gh+��O=W��=S=���#�ػ8�e=�w�<���<�t�<iN+<�e��Ʉ<Qr6���D������Ϥ<��=��.=A�u=�U9<Ƶ
��Y���o��[�<� =����o7���S=A(���D7��D�pNH=��o<���<�W+��'a�Ċ�ܢ<1�P��ND=�N<o=>�:�P�<�#�=�J(���i=��5=���:h[Q��-~�m�5�Ǒ�:�m5��"�ZN=[�����
=�0�:�,T<NϢ���M=�,�8ض==�3
��kD<9�<K$<6s�a�a��N�F�JE=�.����Yo�<E�+��b3=��;=�9�;1�9�J�<"����0�Ӻq�}�T��a�=����Eh;=!U%�c����>=�?�PF+�[R�����v)=���<���lx:~�S���)�K�����ɕJ�L��+����<�����}�*=�J����V=���BD=�[ݼP�$<mR=�r<��&=�����<A�ʼݷh=�9�<!>κ{���@�<)� <G�������v(�<�g�
�!���J��}c��lI=�޿�G��;[�(=T�<�ܼ��5=���;��R���;½L=>8=���z���뼨]�;/��<`U9=�;�����<K��:�w�;����4�Q^\=��Z���<�5�����)k��8/���;�k���Լ����J9�� ἙN��`�y<{h=��N=&�q<�!1�\��[����X=uc8�o���/%=�Q{<�n= �y�7�l�:=\�;��D�Z����y�<�H@=��<E�%�����ۉ��Њ�
yP������N6=�䢻���<�=M�q��<px���,<w�<n�A=��9�mz=�h�C=�=�;��/=r��^�^�6
��4�Z���^=`f_�4��<��V�a��<~fJ�v=+w"=.��<��<���<�⮼�<��<�0<����X�<D �E�Z=^@��d=��Y�1�F:�=�\3�ws�;��F��Bh<� �m�7��v=�%�<�"(�Sw�<�d�;���<��F��]Ի7��KJj��m,=��-�32��;G�&���\��-o<y��<t(ڼ�n�<��G=�8�fҜ��"���<LM(=�I2��)F��}w�W�*��Li=�C��uS�Uqx��;�?�<��@=��;��&=H>=.�;,���<Me�<��������G;���S�4=�Q=�8=��<�#�<�B�����`Q��,=zk�L	�hE���Њ:l{����<W3���� <�*�uüu�`9��><��N=D��:�c��o��U��<p�
<���<&�<j�<=�z�1u3�09<�-�< ��\9ϼ1�@<F{8�?$�4��;83�<���;y'@=�ԋ���=�nS=��aA9�R�v�a��Bu;E&�%���[=�*�=�5ּjk5��<
���q=o�=j��{�<�F=w2�����0.�,.h���ϼ�S2=��;b�;;�>,���e�pD �m,K�7=���ǻ�<�<D��F��N�������g;�S;�z-��^��X=�ؼ�F�~Į<)1t=�g�<�2�<�����<�c��yhs=1�=�) <|+�<nL$;4�`=�!�<��C=��&<�PH���8=i�:5�%�1� w=�k=&ʺsNw=��r=��<P��<��=��L�H�=��<�W�<D=���-��<1wz�PKc=�Wڼ<F=G<ȼZ�=��<ԁ�h�p�`��$;�3���:��:�/=J�����	=x0�<c�ȼh�<�'�̉���<=�3L:{<=�'3��\ļ]툼�[E��P�$�=�ψ<�7=�U;�I�<�>#=Y^k=��<�؍��!�}�ؼ�#�<3.��{]�	��K��<;(@�G�<:mg�1�Ļ`p��p�Q���2=@i#<�u�34��߼�7��B=�b�k|=�����F�!:���<	���X2=�;j�=�p=�<�y=ل�d2.�� =}���^����=��A�:\�֓j���F=72g=��5=��V���=L[�z*��bG��)�<�����t�ӻ��<>�k= j�<_�����<JD����kh�_<�gih=,=�1����<�P<�p�<dH��Q�g=Ѳ<W]x=�?���;�Ԋ;�=K=�qH=!������\�yf��A =��<�Z$=tg<�'�>���Х'�U�H=�}��׃=1�<�.@=�]�<Q�;i�I�s�X�*	����Q=g{g����:-� �Rt��84h�����0'=\�H����'�O��<~0�<�* =���;wɉ�F�}<�_�U=�;��=&Mk<\v�<���<Z�<q�<x���Y�S<���<����)��ɼ9"=0�Q�<��<:>��_�u�Q� 嬼JK<s��<"�	=r��;]"ڼ�Y���<(n���^��<��p����<�8=��f=v�D=뻷�<�W�R)��bp켆�#��`<=�����z=�d2��x0=�11��cd=���`Qh=�=>��mx�<��<v�u=��B�P�8=��=9@,����<Sҧ;ۚ���ټ�d��V;=�֢�׍��m�K���Ӽ0��<{�E���$����<V�;8|	=cM�p�=�'<��u=���;e4�#�)<W��<��<���<�p^�ր����;e��<Ef�*A=X^c=�F�i�U�F!"<ynO�L]�� *�<�7���ܼz����]�;� �<&�<�_�sP��S;�/Z';�G<�V�=[ϵ<�楼�)=�4�<ǥU�e���<�T�<�*�C<�<
/j�
9������T=��;�΋=3�;�^�<;l>=$�F<g��� =��-=Q��<��J�L���v�<k呼-����K=6=��<�0=}�<�}��cg�<�Ś<�_,=�f��%7�1�'�k׼L�F=U�
��c%=���;Pb<�,=��Y=�W=ڨ=R�ݼ����_��=�G����j�k=$��LҼ�	)�<��	�=6O={
�HI��ݞ��R~�岝��[���P�<�=�nW�a�gvL<5�< ��һ�<�Gt��S����}��߂A=�==�]��<�n=5;�<�G׼�Zv��U�:D �b�X�t��<!��<Qeg��m��'�;��U�D�+���6�=��Y_=���<��<6�;��;���E��<K���S</V��f��az
��F߻"���B��o�<S^9�Zi<��߻JaZ= L=#=*�;�8=Ît;U<v3��J���̼��<ܴM�T#]�7
�;z�@=ɯ*�L8��%6�:�sD�`����N)����g;=�:��v=u�;=,���)p���<섘<uÔ�	,=��B=�D=.�7��,?���=U7k���2ʑ<J =g�<�ܦ<F@��(=K�^=E�ż��:��l_=�B�_�⼮�X�s)Q=۟w�t%=4F�<ѠA=ܘ8��o��в��a%<y�=���r];R�5�n)=��#=����@��ۉ;���_/S�%_X=��񻖠���E���<NB�=�f��9y�;[YQ�F񵼓�T�ֲq<K���f�<*v<X��ݲܼ�~q=c��<�q=�+�!-;��)=���<5�������c<iG�<�ɍ�C-/=� ����������=��/=Iѽ��$�F�4�3S!��,=~��D�L<`Bk��-�K<Ҳü�hͼ��<��ϼC!�<�T��P$=�#=j@=u�H����<DB�z����<Ǖ��xۺ�UQ�,���̽Ȼ>�4<��!��+=��Z�A=�� �=�s&�<��<Ѧ =)<<=@��ɹ�<fճ;i�׼�ܼ�8�<.���v=F=QG�:�E=B�<��T=���(D=�>�D)�<�8=�G=1��g-=��?=�\,=�Ñ=����L<�@(<�V��/-=10v��!�<
b(��{μQ2;oL�;�79={&C;P����Ѻp�L��ht=��g��J)=&z�<�kt���:a�;�ؕ��c�����^b��W=jBg< �=�jL��쨺��=m�;��S�w�=~3=��)�[b=�^�<�
)���v��<E\=�n��쯶<�/=�^��,�AU�I�<F�H���_<�J<�i��p�<�l�T=�"=��<��R�������S`��S==�Y;�.�����ᕼ��R=��
��o=���<H�2�KG��"`��:��_�;x�<���<�( ��Z'=C�#=]�Z�c�;`��<p}�<���N,�-}��-�n�;wou=3ez;�l��xI4�v��<�� ��#m<Fk*��C�;�4���/=v%���ڻaHa=YC=<*�<�1�b�T<��2=�9/=�V=	�Z=����<<��8�j6�frW�����
��3l<�[۩<S��<�����8�TI�<8VU=��D����4<A�=����a�� :<2=ep�4"�<���<I�zwB<�3���]���A�`o<�S;��=�H=�QS=���<zhL=��,=H�<���<S�c��8��!��?�Ǽ�s,�A������|�3==�iH=�ҷ��z���<�R=~����ڼ<<�,:=#�<?�<L�n<�<�O
=��ۼ(�g��=H�?��-��:�L(�	�J=���.E�u�z<�BW�X)��r�J�=��{<��O����=�=��H|)�;Q=r�X�.vA<�;x�+��S
;���@�;�'�<�T�����db��ߓ��=+o3=p�ټ���<?��<����7��<G�+<(Ɔ��gi��
	=/�Z�?��*<��<m׼�&Y<L�J=}������.Gl=��m=�V<�H���-=�n��E��@P����_�;p���<H�
=X�H����}p<��=z�����$g��7O=�B1�o=B��<T�S�"���=N����m�l�=;�j�3<��Xo��@�)<�yV��{�<J� =a�<W��=�B/��={��<�����<��;]R;���<[Z�Uݍ<�z����sV���Md���-<x�׼���7�<�9��,=h�l��*�<�HǼ�(<�Sa���3}
={ =_��;����Ip��Op~����g=�$��p{=��1=s��<t�<=����^�q =�pO�o�ʼ<M]��2�h~�6j���d
=M^�z~7=�5=��)=�Ϻ��cǼ��;2r&�[�U��<L���\E7��/�d��;��=�{ <��'�U�<3�=�
�<gzP�ހ6=��=l$<��[=�sn���@=�\O�̆:��<Sڭ���:=�<�(v���<Q;ʻ&qG<�0=���l�E�~=�=e��9�҄=ïn�&�G=����"�R��SM=�LV=��M=P�4�%��K�D�)k�<]�)��x�<��@����<�GL=0,=3P7=�z�<1H̼�3ؼ_�#�<��3=#�G<�.=�����<n7���N=�����S�����0���%s�8�.��GU;_i2<� ���M=$sļ���=�:=g�X�t�<�\�;h�<�ռj�H��#��LQ<�s�)#	�R�	O�<֋Q�;�����!��}8��P<&~g<i�'���H=�_�<��4�U@���o@=�X�9@SC�2s*��a<�m����<��;�k����;j,;�\"`<��/<��=�d�;�F���������9�I��9"=K�=��p�����Q:=�DA=Y�:����4�`=�KW���7=!�<o��;_;��5/� N�<S_����I=��~<r�C�i���� �2�=��3J�����T=�X�խ%=���<OL���I<Nt"����N��<�/=�2�<G�=�ZG�ʋ����EI;�6�2}i�R3Q�.�.=���;/=͔����=�f4��F��L�<��lr0�,�=G����r��G�����l�c��B�<b��<�K�:��*<B!&�&=,�!={R=k<���\=�J`���<�4�</��QY>��B=3�W��R�s�;=6�r��)�<��p�r`ڼ�=ˤ�l/���T�-���g=�d=5�7�����6=��<���<P4�[�!<5Y��*��<%Z+<��!��'=��T�z�;�;�;!��<�݋��) �m��<J�d<1��<��S�8� =�}===�U�[<l4�<ϼ��W=�J�/ѻ�ż��?��ꚼ}����=��i��1��V�v�|�=QW��dA�3Q�F�=��/<�c�����g�<��/<n�^�)���v;<�N�D��C��O��S�:�*��q_޼�t=G/�;E���e��G�=[����^W;!��=�<=e��<,���+ռoGn<fÒ���^��Ÿ;%R"=u1=�VT=�(�<�xR�=����� W=��a���<p�#=�+=��=>�=�S;��S=ና��)=Llb=BK<(.0=�S�=�jA=��<� N=�S8=0I=��=7ת;�(��a&����o�żE�:
���mb=�l�����O-����;:{�<o��<U��8=��<�V}<'n�wG<�1�<�л�P?=7�� ��lO�}�H=Sh���E�<�����MJ���+��5<=_Ю��ڙ:**:<|�.;�gк���<)�>=N$�l�<:�_='!=�</���#=4�(=w�P=R=��U;v��AxD��-�<�o�;�
?�)��w�W<z�ӻ�1E=T =�ü�90���&�BU+=���<�00=A���(<�d��F='��<{h=�k8���<
��#$��L�b=�?�<"�����}<֝)<%�i=;]¼ �S�y>=�4^�M#2=l�A�=V���쁽SA�Q�5=���'ټ�Լ��<hJH=h����<����;�:���a��M4��{��rȀ�U����V��0�z =)\ڻ`2=�=N�<O�<��Z��-���M�
��<&����q�Q�o<[o�;1,=aJM=�f�;X�h=�tP=A[=�i8=���S�=dP��d���<�]I=��=�- ���<��=��=�X��I$�x�[��k��ڐ<����w��}��0;�z&=��9��־<�̥< ߣ;^a��w�M���e<��5= '���Î���d="IM��x�<�*=6�F=�Yd�s����Q�?�(=��hsk���T��u3=�VP=y����Q0=�^)<o	�<��j�����#�b�~���Qʼ�@�<CS�<�M�
�;���۬�<��%����`,<4�<��=��*=pR�*�=�RԹ$�@=���$����&����=�e(=��^�Z����л�J<��=���<��<�<�߭�o�[�tU�p$=M���Ҡ�5⼹����.=D���[,=�-��h�=5��i�t�Sߨ;(�ּ���}p�Ԉ	�$W��N��<2�ݺ�=���^�g��,ؼ���<�rG��O[=vMX�7�,=x��<	;�+���Ѿ�<�e�;�w'��aѼ��$=��<�U���<����W�0� =���J���㭺�6=��<4�%�T�;]�<�/"<oQ=~���an=���r�=��b���<�=q�
Å<P����K-�?O7��MR�Iy�<���]j<�='?=mU(�Т��d=D�ܼ1�;|j��b���)ټ%��֑=���<��	�5+�<0O1�OVP���E;�����$�<� k�b�,�z�Q<�y�<�P�<X�<�S<�D�<o�#=�����pB=��3�[=<����d=H�8���e�(�Y�Q%|=g�a���
=Y =a�=8U��H���Q=	�=<U�(�n���U9=/���E�<�=��b=��(�e��<iμ���[��n�;��C;3�t��|�dq�<��D=Q�;=ԑ�<Nt9�5�G=���<GἾ�s=����V��;V��;�W(< ���漱��&��<��)<�G�<��1��n8�͉��]M�u�:���=|�<РZ��:=c��<cP�2 =�#H�?��<8�|:�k�<���΂*<���;}0x�7��5=��8<��<X���im;�!=�r=�]�9�E��a��% =��@������]���e��h��|�jt�FN���:M=)\��;=�A;����x��5U�<�z�Ƣ��qq�<B- =������	�!B<4A��W�J;�}o<���)��<�k=��%���`����ܫx����y伴�=��ӁO�'CZ��e@<`q���<^��<�X����(����<���L,��z�U=�Ċ�]E�<�a@=X3Z�����Tl�"�<[	�<�iN=��<y�=u)$=q�^�Q��<1�K�����$��mw�����<����S���+�ɒN��n���K=�O;=���8�<�+�7�b�M��<+s;�!V<�e�=V���Z�<(wl<v�=6⻍�0��;�� U=��=
�I��f�<aW�kv$�4"=���?�t<�g*�}j4=��]��Cy<�1=d���Ҙ<O�?��S�;�NE�~͝�ޗ<=P`O=�=��R=�ؔ�DTǼ�+���A<r^1=��<$��H6=�NA=:��#a��c==ج�<���<�*(=����s�ͼ� =��8�+C�2�����j��+��ߢü�o(=�%=�o+=��"��?׼��F������]=��b�~z�<WS�7�<$ �W�I�˽<Nr�<��?=e�����:�FӼ��9��5=n�8���<9�t���;�s=I�~ =��Y���k='�%=͂�;���=�	��24�2?N:�&��WM`=�v ���I��Ǻ�h���=J��;Gh���=�=6�i<͆:�1���b=��<��(�u���e��?�9=�Y���/�nZ㼻D��W�Z��n�<�|��"·��vU=���:}Х<Pŧ��G�;`[�=iQ��LL����<�o =�:�;%M=�w�<�r9�"C�� =��8<�w-�2Dp;m.<JNo=��8���=>O�<���}��L3=v_�'N_�F���=����z<; !�&���i*P��1=*����Q=�߼�b=�B=�W=�&������So<����%���{<�x����������;�;U�:K�8��N�<R��<�ӈ�,/�<b*޻++������r��]d��E=��[=5��&N=5�)�&=��R=��A=^+;��c=C�U��[:�ɯ�< 6�<�o=�ټ��� �������L�"6 <Hً��
g��;@=�qo�U����a�;7=���O��;/����o1=���λ��6����<�u[�~zd;\A"���#=�p@��B=TT�;=Nռ�tC=E��;/��<mƄ��d*�V9I���=�j4�)曼L�c�v�t;IE����6
6=t����={"o=��F�>�<�E���.��=2ڢ<�h�B����`�<���vY<=g���e!=DӘ�WT<����#�";u��<Z�&�ŷ��B�����;<`k���h=�q�;��2�!J%<���<ʓ�;���<�=GS�� $�<���:$*L=c�X��y�@�o��d5<���<��Ἓ�9-aZ=镘=7��=B<�-=k��<щJ��]�\Ev<4Q��2�=KO�;�Aټ4��;c�=A'={Ql������#=�ch;�d=d��<��<=p=�W��h��;��<<��F�%q@����/'<��<7	'�xBb==%<��<�$˺<�P=����ck�<��x��%�<}��<M0�[4.���8=J<�<,�<�J=}�J=��=�<�O�=�=A�/=��=��;C�R=��=O�U��9�:Bm=e(<�tO<J䘼u<�c�8z�=��9���;���H�<�9�<C�κ=Oʼ]-O��)2��՗�-�K=��ۼ\���r�kq�<�K�߯�;�f�;��=�>7<H�;=g�^��^%��Z'�,����`��֔;��:=9q<b=�>�q_>�6�C�<�v�är�T�;D�=��S��Z�Qfȼ����2Y=^�ȼf���X^���2<�dۼ.*��=�=�I<�Q���[�<umN������ѼA�:�^ �P��<���Igػ�Y޼��9��6:���V�EN��w�a����<���=�����_�x�,<��=>=�)<�ZD=�^;�׀��?=���v4�<�5��.�T�;+����Q�4 ��:>�'���Q@�<�E�8�(��)����;F伷��<(�<�<�5�<��=��M��\T=D�<�4���|^���:=��<�L'=��e��O=�8<l���i�*���ۼ�Dh=�)�<S�`��������4 =ۊ=� 1=HAR<U�;��4�&^)=��ự�t:�O�<�D�;?!/�������vP�U>�;�r�<ߞp��Ô<U;�#�=nɣ<�l�<\��<'���D�d�ͼ����[E�,𱼞�<�<u��<O�i=p�L=H�%=�8E���&<��2���:�D5<�SE��o�<oν<�� �
A�;�d=�᲻���<�ҧ:��f=��[���0�46� a�<hܼ�h׼�>[���i=f�=k����P=���<[��<#=���0�_ݹ�MuV��o��?��;X�%=��3=�<G���<7Ha��:�;��)=ݴ==���<S/�;U��<���L�w;)�ߺ�"�t(=��!��@ ��D�;>/�<��=/���� ��9�f�5ُ=�&�<�n=Q���T$=�˅�������<�WX�4�Y=��<b/F=WM==�$k�ysݹ1'�<h1��7�=v+<�K��̻� �[<�Uݻ<"�;��<ı�<*<�0����ͼ�{='\z<���F<�>=�p�<�V�DUV��3=�,]=���6=D¯�!L4� ��<Ƹ�:@����{ˢ�O�7�>�<��N=vS�<n����U��2ռSe�<OPm=B<-˻���<x�=F��?��YK�?�$�l?=S�=5=�B��x=ǧ<��*�莊��n�<��i=���<`x�<δ=�Xa����<�7N<�];=׆/����<��
��f�õļ˘���0=�m�<��<Ў�<`��<���A�ܸ@�&��ͅ�o��!Y2=�<����<�1����_�D��^:<I�<Q�x��u=���'=�>���8�G���g��U���=$WӼ�QM=�/��\��A�@��;\�Q�HR�<�y<L�{<"dѼ@0�<�ǂ<�I,��,�����1��=��x�R���q�<���:1Q5�/CB��$�iX={�N���l��]=��<�D�����Ӽa�S=q�+=�c�;�RS=^gB����P�<��M��]���o�d�<��<C�~<W��k�4���Z=��<<?����*(<����K�����;�=}3���z<qh������YaG�e�e�Oڼ�I����K��e.�����)=uU�;,��;�=ZP =���<�+���h�t�=����<�[�O�xM�¢�<{��;M7�2�H�b<�6Ѽ��F=<��<��=�׼!��=�*i�2`=xA<�CE���
��� ���H=�t��j=��8zB���u�Cµ<e=����Ji�<��;}���j�a=*�x�.��G���A�3̼߻C��v��=X�!���;p+%�p�o���D==˃=��5=J��%�������b�7=�$1��Q�+��:�� =�qV���Z=ԣ����<9��x����ݼD�=ݐ0=L9.�!�=������<�`��J=�Sh=f�ż]"��P���J=�{�;��c=9�;lC$=H��;M'<?��<H4�;�^�< 5=������]����9=�5H�[Zj���;n�D���x<I=Aqe��,�p+=�M⼬�*=�V�<�7=-S�ޚ<]��<	|�F:n<?�������!��1<D�?��NҼ�-���:=�?B���=�M�\�]<�/�� r=��;=��<�q��SJ�<2.=�W$:���<�M=����6���t��'=���<�7�����
�Q=�U���=;� � �����oeC�Ut=�q׼�-�<�}����P=@SK<��D��J=�G�����;+�A=�*����<AHh��h�;/aS=�,�ʘ<f���z�;�Va=B��1�U�I�a=E�;3�=qr��kZ=�+�<(�u�L�k�P�.=�!L=k�#����<G_P�ԏ��H:m�ݟx��9=�i[�;=��n<m%�<c�t�'�;<���M�(=�J�;���m�D=�����ɻ.D$��j==+76�<Q=�o=�E=���<��'=e��;�+��d^=Ie���<Ů*�#@��|��!�<�<�5�ͭm����<�3 =��.�f&��ΦB�Y���/�2d�;F��0�	<�?�v�p�BgO�K�[=�
�;{"=X�0=e%|�u�H���=�U#=h`=��Ń��������~���(�#<3F?=)y=�JU���%����<v!��0��h�<�⳼J�=.>��|�f���)���� �ݻ��i��
�F�=T&<�p���/���^�<J�ְ����Q=���sB�F��<7��Pf�<����!���� d�_2<<�sO�����,�}<�{޼��-�>�:�g�:Jd� �<�fB=���<n� �e�Y=RPS=i��<��<SUN���=M�m:�-��e=�D���=��N=V��c s;��7=O�f�y/��=�}ֻEM<���<r:8��>���*=N_k�I���(��
�E�o�I5!<d[��j@���=��Rja<i�=Z�`=�t=��˼�s��V�l���M�<��<�;3��=�	c=餩�瘟:!5M���~�+��=�|%=�7j=��<�����5<��;aҫ�b�;V�\��A=rb�9�����O��?;�$ 5=h�9=G�;��T���F=��P�P��N��F��ό����F=P���0�<�c:���
,��RB%�姣�j�a���;H�C�M�D<���;�ȱ<�l��{�Y=�4ݼ��@=nB�NBh�۝2=<=v=�-��=G*�{���z6=���;�.�Nz��h�>���<y{k=3!�<5$��|�Z�j=~\=a�x���b<t��<3�=�%=�I<
c����<mM\= ˎ=�
j��~P�v>1=���\�;��š�N�F����<�&g=�ڑ<U�3���=�ʇ=��u<�l�;@^=�zi��ټX�ȼ���;� -�� �/���-����4<]_��w�<�긼֌
=QQ]<B�m;GK�b*�(�N���=����pK
<<��N]��s%�wIE=Ӑt<w`�<a�м�,F���^��e�1�I����1�w�&�j<�4D��E�<8�/�t�L���;�L=Z)=�o���H7��R��m{\���	=C�<��L�+�0�dJӻ(4/��!��<.:%���Pf���<S�M=����#=�YU��-�g%=���<��4��@��Rb=7�=<���<��*=��E=|���������Q�W,�\0!����<Pu�=��ü����?�<}��;��<�<�<v��>�;�<
z=C��<B�A<e�@<G�m�����s<?k=���;9��RU׼_7v��LC��B=�f�<��D�� =��="�3,ۼ��i�k�:��J�^τ=�~�����w� Q2=],2����Yмe�<�=�T�;�\E=U�<9$f�0�~��g������i=^��[��@8f�~b+�^;7=�+:�
=[?=R0,=��=�/=s�J�`��<N���jmؼ{W�:åܼ@�*=M�;`��0�/=�=�!�<0�=b��;�_�<�|v=X�=߼���J���7=���<��	�9��Y�g=N�3��\	���$�<��S]����u;(��9����B�N=�����,|�x���@=�D���<��z<-R=t`;���KG2=P��R\�;
�='|��/?v=�ɻ���͸<�z�]"\=�D=\�<��2=a�<N�/<>9�<�2<~�|��7=�̨<ó"="G�<(UV�x�f���j�� ��9�<�-�<�$;e~P=�u��H�є\=�;=�j�����h�<�)\='�$<��;�v��/�������<P�ɼn�&<l'�*�0<���<Kt,��Η<�F�<���<+�<��<~v����<�?���e<�:��7�;���.��;�;S��<fǩ<Є�<�g�<��D=��)=�@r:L8�<U�A;85=�;�i�W����<�6=����d�m<t�g=j-$�5��<�N	=�V輻�|�Q�P���� &
=g�h=d��R�%={��]j�<�{=x��<4,=\�ӻ5D�0�似�c;VjO��	q=���<��$��5.=���$�W<tՂ="2�<� ��<��N��T�3O>�c���i=�\"�k�5=c%=p��$�<"���Z<��	=�����B=�k;�(=:;�<����Ji<����Sd�A�K<�Rb����47�<:�(<U;�'Լ]K��/��]y�<{$'���=�a;ˣ�N��<��<�[=:51� �H����-y�<�;^=¢�<��;��L=��g��3=h�c�tA�Qq-��h�<�˻�f�A������?k��.$�W�G=�:=ϔB�Ab<g���F=+�<J�*=<te���v<�С:}p=O��<�/��=;=z����J<���<�:&=������� �+�I���Ǒ�<dy=��Q<�un=gia<�re=&QQ=���2�<v@��P�������#";�k<��h�I�0=0
�<X��< l<�y�<�h�<� =x����=`��</=:>����<�,=�&�������F=�<7��*�<�O��[�c�弭g%�=��9��9�˩_=%=t���/�n=��7��
���<�4�%)H<f�=?Xv=�ْ�8|ݺV��<04����<�D����������6=�*����ks�<�4�<��=�����1=��&=1T�:�#�<�tX:�7H��ӗ�}��;l�<`]c�`�Ǽ�_+��O<=A���N�s��<�iV=0:�<�Hx<�$����e<���<W(_;W[d;A\�:Pt6�`�<��<���<B==�>����P<	�Q:�l6�:��bE��G4<�!�^��<��һ��E=��<-b~���=�8-���U���,�;�#=�=�V?�Wb$<�C�+�<5�<zHR�»0=Me<��������'��=$,�<��[��t޼)�^=�?m�R�F=1׻ӽB��B���@��,=��=S(=A�=�	_���0����<�c�Yg�<��%=��Ѽ�.=�s�� �؉;=�l�<��E:��=�)����������U<"�����<pl���=c%Y=��c:�=@�l��<������'����'N<0�=�x�	���P��3߼��<c�C�@�����Ѽ�,=	珻Rpk<%����G=!�<="��<�;��V�<- 	<�~�<<�<�x�rW̻�ȼm�H<����5=�b�<�|����;��Y=�e�f4����<����5��s�=d�e=V�.��8?=��\=��<�m�;�"�b{�)[(�ɋ=�ZP=�t��t{<:%=����|X�lQ�<BQ(=��!=��\��<�Ą<nɹ�E=;�%�cDp=�ļ��<O�=������y=�ێ?�*5P�Є<#�X��w/=Y�;\��;ʝļ��Ǔ<�E9=y�w=�ӈ<9Ȗ<� T�!�v=�x�<�V=W&�<�	=�ӻwKʻ'�=�
�;���-�<s���u^K��{<�	��Xw=��@=��9<�`7<{ܑ<�Z�<a�m�;@�.<e!���=����\�.�:��>2<T��=ϢԼ�ݼ��B�d��n鲶�����V��c0�1���s�z=�eG��:s�;ZS;S,#��8���n="�׻�S��$ռ^�*�o�P=�Ve��1<9��<
�<[�2;�9����-�����jL~<J�=z.��X��-�<����J�2�7,���;<	�B�;��.��\F=�m�<D��=6�x<`�=�^����0=���<��<�PJ=�9>��+��z�ͻÑE����8:���=Y�Y���&=k�B�Q��<��<]�\=y�介�(=��1��^ǻ+�	=,S`=�=�o�*j_�Z�%�b��g<'-7=�� �o�,wA���x��=�����gW<u�aӡ<�	�Pe=�
U��<�"�:U8�+s�<@Ʃ��c;�a�;�S �_b��(&�<��b=o ��T��5�=�P�=ַ�<�T�O� �,��9|����f�c<�<<����=dP<�R(=�<��Z�d��?u=AqB������<=Cu=��D�h�-�/���{>�yU��k�<$h���2=��_=�o9=d���OY=
�/=��+��bS�-� =��)=���Ǫ<������<%3����{���<=?�<2F�<��{<,=���<�i4��<R=v�6�H�5� E"�p��h�K<I����&���;=��	=.�<D.<�0;�5r<��E���!����<��:��y<��>=n�j=�����<X���!�P`��4�<��d� y��k�<�a=�}��PT�<�<*�!�$��/�`|��Ѹ�<���<�'Ƽ��^��=�I<S=J&�d�<�������� =ƀ���39�H=C�&=B��;�f<�u-=�zt;�=-F)<�g<�.�=���Oa�؂u�,b���"����a=4�Ƽ��+��#=r=A^h���#��$��BE=��=`�=,�	�V�~<;#�=��I=��T���<Rŧ;ڤZ��la=�4�7[b	=��V=Q*=3*��#���燩�{VT�~�o<�A=��u���7=é=�D�<�=ߌ7=�J�<��;*�����V�,��p�w�j����<��~<U�y<�����;$����{<�((=�S�<����o���'=�
�TO�C�
��6~��lm���;����9��<`̼��2=�}�<�7�D���B�z�o��L
<�K<�?��
���h=D�d��׃<�����y}��B�UaG=�$=��9�'HR������=|��(xK=�����%ݼ��,<C�=.7C�)�=�g���[<��U=�<=��<9I�kVP=�&�<�<��b=&���!X9=�W�<��<ȁ
=��^�s��<�-]���;���]�<�:���j� �.�	��I=�~������9׹��<�l=C�޼I�<�}��"f��3٩�Ls�=:7=�F�	�<}�C<�aW<8�����D�M��1�K��6��/�:��=@"�<]�=⣼�8;�u=�/�<�1~��z<�B����<�ޥ<T�ú-[<�;aW�4���4=�q�:���=�
�<�:)�3��=�U=�s=�����!�$�ܻ�`��d����>��,=q�޼�2*��U=Бn��i�A%�·���x�L=|��<m_0��-;=�����;��8��6/=gŻ��D�A�����]����Qm߼zpL=੖;�;ɻly�|��<"ԫ��ʽ���<�8���A�<E�j����<ȵ1=���\R6�R�� ��<�9�<Vca=�����5�i#A������ͻ�<�>�λ���ü�a�<x�󼚟"�!�7=�s_�Z;�=S� ��-=y�À�<�=��G�,=�*�h=�%���4	��$黉ex��`Y=R]�=B}<�fV��� �0T=���<�WY=AW5<���+��<�X==Ǽ�<1�cB<���<�=!�<0i5=Wּ�k=�l��X8�<�}�I�)�x��Eg�F��<���<#��<�F=b��Vz��� =V�\=9��;<�� �sz<�P=�[c������*�<�`���[����<�r<��}<C/#=��W<i��;�}����W�,[=��<��=�p��O���<J�b=�M�=
��҂A=�����=+��<��(=�?��y��v@Q=3d�%�H���5<��W�'X�o�p=����Xt=�J�;FJ=c?��S�<T&�<Vm�S)�8�$9���������3����<!�<p4=���=��<Ol��,���jJ��4�.8=#P=�Y�ӡ��kbͻjs�=�������f��:Z�=:Ӽ�����XY�;
A<��<�N+=�1'=@=�1@=�=�,G<p�T=�m=��5�_���8N=�e�&g_���Z�c��:�P���;�"Q��7p=0��<͈,��b���<q(=�c/�L=?��<���6u<Ñ���<�-X��	�뼒=P<��'���0�F\<���<��<6�&<���Y��<_D|=�-�<6�A� �����<Q0!=GA�z��L;��<{R�����<{�軚%&:h�O����xI� �I=煨����/�8<x�=�+;|�=��H=�����fZ=�/Ｓ�U�ى ��'�;��<���ּ��.��'���B=Pa=�W=�5c=�'ϻ_�J�!=���<
2��e����Xѻh�6:_�<"Iv��L̼�[���<�=��(�P����6�x;F���8=�G�<���<�.9=<	;� ���y��S���
����;�8ȼ̴���m;�1Ҽ#�Ӽ�'W����;��p<,J�<��r���[<���<��<OA=��<�1X=Pś<�=�=щȼ�:���K�<���g�= 1y�K��PC�;x��:�9��� ��FG�;�c=n�����<<aτ<�RH=c����<���:��;��n;lJ=#l<~g>��8=�<κ��=�/M=�O{<��@=���
v���<c��=B=��{6�;��<YM=�;�}�����v_�	G�;�9��{=*# =VB�;��<3@��}N=�x;=n�C=�l�;s�N;�R�<O�=�]���;s��<8�4�F�h=�t�,�;m�Z����H������L��x�<׶�P^��`�ˋ�<R�<WBֺ��u=	�T�(q��	�=�S=�@x�#d�2�	ݻ�k�\<5Eg��^<�)�<]��<\�;6zQ;���<f�==�a��qλ��xq<8o��B��8��^˼�5�=5~8��e~���<�b=�n��<=6[=w�ӻ�Y�d���X��iVc;%*�<DA(=D�<e]-:z��<��9=f�K����<0h8=��H=?7�.���&��%�ܼ>��<p�9==�<��?���<��E=���\�](=𘕼�\���CF;ܾ���O$9�)�<5*���r(��1<��<�u;=�u����:�]!;���e�t��|;�OD<<�Y��=f��<݌+=a����i�;�ޒ��Ё���g�p���<đ^=o�<^y0=��*=���<d�<��
=k0�-�>;�i=D]�;�X=;2=wq�=��/;�1=�p=)
��HX9=RQL�$�=�Gz	��&=с������D�i&���)<��?=V�����%��Ǽ���ԃ��P=�46���<���ߦ=�k=�qʺyn�<��P=K�^�5����(��Yj��g�<���!<���_���^�<�=4f=?�=6��;��=.�k=QLۼ,���v;i}�<��=e���#�;k�b<p�����O`�(4=Ώ�<�a=�}c=C=�8�U=U��<���2�<�K=4�H<��r�*(S����;��e<��S����X<��=�M=3��<-��<���<�3Y=�����W<��R<#�I���:�'�9�21,��5<i�<!�<*�:=k{�*�)=
��{I*���t�.�~<��`L7=U�˻fG�ks(=fN弲���n���[�<�乼���k��; ��:��;�Ls�vS��?�;!�<>�<�m�)W=/@����n�*��<�>�<�����	=��ۼ*����x��:����ռ�*R�]j	=�'��Ȍ�e���`=�"��5	=f�<'�=��Ƽ��6��U^=�f���;/�C�s�N=p0�K`T���m�a���W� =�w:�)=8�5=��a����d㪼tXu��y�<���呻ON��A���l�=$���F�(�<���U��<�H輴l>�rg=ҍ��)�;�$��ml=񴽼��<[���Y��Mm�L���}��D=g
H=��6�J��<A�<si���#=�N��z�<ku�%Ĥ<��=�#O=���;�"%;�o=3F�<ٔ<���i��N
=�ĥ�|B�������<Z
<E���0;T�<��L=�~	<z5�<)��<��?���u��D=�x=U=*)��1�<���<X-"���`�=C1o���#=�a=�'=��=�%A���G���S<	��<>�?=��м���<p��<_)�����<��q;�
{�ݽ�<^�t�e��h��<���%��?>�c��;���{�<O�@���J8��~�<��%=Tfۻ�;=��R< ��<�S=�,I=�==�~k=öW<��f=4=qP��|ͻ]����;%� =�m��U"=}[.���Ѽ��a���(��/L:c��g��ho��Va<��6=B�%=�dM�W��ຕ��m�F����<;&x=���<�l<�=<o7���\�RZ�=����iq=
��;�3=��������<���=���.����<=����Jc�<v��Q��<�qf�/>���j�A��<d=v�ȼ9D��������x�l=������X=�'�����F��㧼�d5��뺼�9=�GC�J)P��.X=r�Y=�<Y�d=�|Q����b&���i�Yk=���<8�<*���hdU=:� =�z$�ڂ�X�S�l;S�c\:=�w�;�� =���aM＾O=�N켝�R��X[���c�j�$�9\�%0=�/S<�"��ҁ�<��l=7b<׈<� �����镺r #��z�<k.H=*=pW޼ :���<*\�;z������tLѼ/�<b�<��<�4=G�x<c��LU�<�FC��78��k =��<���<��%�����o���"�_�Լ�~H���L=Q��Fx6=��h�#u�<Y����=�$=G?=ר<��-����=pS�<�A�x�l�!�B=�Mn=�="WO=A�J<s��j�l;J�>=b�'GE=�.��mZ�F*)�
>@<�<4x]�c!�<�cB=4�P=�U�^��<'̼�A;�I=l;:=�5%�XU�<[�<��<D=K�=,e�ń<@U�R�< "�T�㼾F_=�AB=�-�=w��<	ƪ�rJ�<m�A��v�1lH<�7R�i`�����bP��=Ixq=���\(߼��(=+L;��Ἐ`<ip�¦��=O3�Z)�<�	񼟄>;�u=IM��xMD��J�<��<�;?�Vuἇv��^ :vf<�����CU�>R=��V<�f��-���:W�<��0=���<{���]Ju�-;X4=�˼��߼B컣�&�Z_=��>6����#��
����N� ���*=6��?�<��<^|<\�J;
�2��I1�`�S�0=�`�<^kK���3�Jb黦��<��~��<�-Q���g=?ż����-�>#Z���S�H�.=���I�=�M���'=Ϻ�<2�I�R>�<�(����v�لt�
�=R-=ҨK=}�F��-�<�^�<�b�{�=�����=Q�;��<�;<�/=�(� �-<	�;1�z�9�R=⃬�]�E<�p������4�<�ڕ<j� =�W�v��IK�;��3=��0�� L<Sj�<�l»Cճ���W=�$�<{4=@�ɼC=���^L�>���繃��? :<;���"���=Av��t�F=�R�q~S�kV����<5J���Y���T�<x+[=���<�b����Q<�ZP=��\9G�A<>�����<e9B�5��:!t<e�ؼj��<\P�<Q7�;k�<�K=�c.=�!$���v=9?���'=`�G<��<H�<Vμ0N�� 
=�<Z=���;�v�=�>��䟼z쳼^vE=��;���E��
�k��v:ͼ(�c�:yx������(l<�n=��Ҽw��<�2�]B(=2�-<2�=�K�Z=�?=R~��=ұ4=��ᐳ��^����<��<�L��a��<vIm:�P)=�U�<���<�>�<��	=�7��UQμ�u���mb���)��r9=�ur���w�  ?<�i=���=).��Qg;��Z�X�V�$o��I�?���T��
<��_&�;+=D筼S5���o<tZ]��qp�N�]�4A�<q�Y=�=	�;+�_����FV�v�i=�y��/[@=
�/���U�۞�<-
�<�=Z�^;������<)�=h�ƻ�g><���<�ٞ<8O�;0iv��L�Q*0=`�J���=���<9(����;N:l=1�<%s�~��&�'=�t
�,��B_=���	l�<ڷ ���:=w�@<x. =(G=Y�����<A�K�eV���NƼ�z!�jsR<FI��w<�7	<N����:���:�j��n��g:<����׼��׼22�߭�����K>=�l<!T�������c=�FR�N9�;�xj=c>@=��:+0���X2<(=
��<��7=����-����i<=�9Ɓ<��Ƽ歗�<�<zbq=��;��r<�H=�=X&=��1�y@|<4��<�ϛ<U��<\��l=>�<�9���:��9�<�<V��<	�3���<��ѼN�3��m^=�+��L�|�a�=k�<YI���b#��O<��<�%�<{��<�=D��<���<�@�iN�<u�s<0�O�!*-=��}<E�<��５?M�OټX�C���S�}$�<�/컓S���C�q����J<�n;˔�<m=f��ug��X�<p�<�:"=�a�<]����h=��߼�<���{���F<��;K9�����}�n=���<���X;�ϯ ��4=1�|<w�;���<��Q�A��;���j_=�o��z���Q<I�<}�-�i\�����k�/ٚ�w� =�a�<����$���#:p?(=�=6V2��.�<��L����<�,=�;ʞ���=��y==X��<�����|��j���Р�<����bS���j�TU�<�1�<�')�X��&8=;N�;D�@��Ҽ�μ��<��y��=��Y=�}�<�*��?�l@<�P�<@m`�όu���o<d2�<������<�}�<F�ԑǼ�t�<�EE��L�C�V���<G�����r;? �<66�<	<�ܵ����<�;=dR}�u����!��=ϼ�۸<V5�<�2�;y��|ޮ:;Q�j^'��������c<�� ��l:�D����}=����K=S�='�<��G������\<�Q(='���R��;�u�<�N���;D�Ż��V=��뻘���ڷںg�2�NL�V`S<a��<��P���N=t4$=3�V���=nc)�f`W=(�X�J����=�tb���<	L�;������nS=�=/{�;�B���Y�:�0=)��9�P=�<���;mK�'|�u��=�@H=f2b=ʢ�R�=;�%9�O�<�b��Z��]=2�?=��W=du~���N�|���2_�<29��B�=^� =��<eu�<�W�Ꭲ��;҃��?�+=���;$R���*F=���;_�d��=�J=�>�'��<��/=Ĉ-=b巼<:�<�{�VEA�P<�;	z1���Qp�=r!/<�R?��g;=���<�2��%����,=w��;����K��/=��'=ER=�iٹ�= =�{"� �O=:?#�8��O
�=>��<kuY=	��<�����t=%?�;w�4��bJ�aܻ������o<)����K���f=�F���μ@�=PY=���4iu<��}�a=a��+R^���+=���<��$��~���LJ�8�<Q�ϼ��P���ԼfY;���<���;a�U�wZ=7�O��
��g=���d_�nQ�(�N��\���\���m=�Z��d\&�>������E�zK�<;Ba���5=$S�I =�!�<�}⻮Yq=�꼖=�`���`�jm�P4=Â�������M=� �W]<1�5=#�M;X�#<T =F9=�B=��4<CJ>�P*#�S��;+�+=��,�!{�;�&��ԤG�^b7=.���\+���<_H=�Ѵ�?��ncG=	S�m��=�xe=Kv�<ぐ�ƟT<޵.==�h���[=��b=�x��B$��Q�����<�<EM�;t����K=�8<b�<�<���<R�9ӯw=�U=�D=7��<`�Y=0ɀ���A�`V� v%�I(9��E=��(=ɒR<њ9�����+.���;�:;�4��=�H�<��?��_E����;;~�<�(U;�Z,=�3���[p=�<�?=�6$=���<T`K���<�4м[�!�b&�s܎<�8�<$�_=h��<�T�<
ȼ9Ж<�G�m���%FP=r�X
��8��<�o�<�21����,=����y+��ʸ<��$=\
=��=sgû�<8��U<�F{=��<�BT=Џ�� ~ ��=mx�;�6_��% <,�<�=]�=��1�H�]�_�伋rz�X�$=t<�j��!��~Ga< Q�<�9i=�I���=�!< �A=�f��X�<2��׍l�{*���#�<|Q=�7��,�
=��&=��H<{��<Ɇ���yE<j�$;�#=p�%=)6K< ����:�C<��L=��ܹ��}�&���[=�-�<ϭ�<�^����$�W��<�ü�%X=k�@<Q�~�dNe�&��<0E�x��ª=5)�;�	H=ZGY��=�<[����8=��_��6��~�<\��<&c���R���[<QM�<z�~���H=;1ûT�[�L�M�ռg߮;AM��4KB���J�P�1=cyf=d� <��<u�9<�H�渝�Y��=�=����N=h��<W�����<~]�m���=b4�<Cq-=j�=UL�<b:I�5E�k`ѻ?�v�AXX��&���<g�/B^�Pp�;	B���9=z�=� ��=��b���G;��7��F=e0���4��<�̇��#a�C-�<��b�V�<T�x�Wu��=���"\c��CJ=����p缹�Q<��k��c	��U=q�r=��b=<���;B(1=�vK<o�|�o0�<�5-=s<NdC<��,=wa���q�^���X�0<[�9=)E��gԻH�:C�;�@Y�M�O<'�3=�:C=���$�=D&=�'�h��<�_A<��f��I8�~�o��I�����<0�1�R�=2P��U��P(o<�(=^9Z=��<	�j����X�b=?{Q=��	��)"=h#E�}�%��O�<��<�8G�yzz<����S<p�a���D<������<���<hG<-��P=��=$u����+��?@�ь=�<O=��,=���eX�<���ͦ<��h=>X=�ϴ���u%6<��ͼV�=�	r=%a��~V=Y(���r&�"<w�;���;�뼑_�]�=��3=%3/�B �<�(�<0�z�=_����K�T.������r�U�<�w��neۼxHX�Oz=�K=��<=<@�;�� �*�3���<4@<Y�����&`=?�Y=� ��r!q�㲈���6�K���=~5F=�~�<a�2�1�w��LF�T�g=$�Q=��d��_ɼ��T��w�<AS��xQ�f��!P���d=�8<���<\iļ���<��&���=���<����ȍ�;@$꼑br=x�E=d��<P���ņ��I �x��<��<=�8�<��1��<��_=<6<��`���d<�Iݼ!{0=8�k=;4��+�3�0l%�w��<����7<��`<�~�<ձ�<��6=Jx=dM���={��<�O��,��{4����m&�}Є��񩼲\
=eVo=��=Yp=��=�w�c���+���==P8��<ȼ叁<K60=`h*=��<?��pP�=i�<�|�;o�?�UX4�����?�A௼�~\;6L=)�|�MB ��z?�F.d��D�<�<J��H=f~�<^���"�.�=y!����=�W5=�S�9vH=�=d�<�U;=�w?��"��<�t��O��<V�=
�k���<��_��G=�|�<=��a^Y<w
P��9=���<X��<2�<�g:=�≽m�A��=�+�<���<��U���$= �+�3�;�aY�E���e�-�W1�p=<YB</�A�\���:�<N��<�1Q=�������p���)�Pp�;Ka-=�;�t�:�+=}]w=�$_<Vi;�<�kG��	=6ʼ�m���=8W�]�e��.�<LOb�O3��K�*��;w�:�=�5=ȳn��\g=���<�cV�O�J��VI=!_\���a�Z3�-컹0��mݼ�D&=��=��m���=S���fΧ<��i��T��`:Sx�<�P��&^=��[���߼��X<��ɼ��e�顉�w�i�6|o=J�z=�y�<�����<<�5=j�"�nkN=����*�4lS���=gI�E�=~�,=�D%��ެ��TԻ�G���ɔ=��=�~^��=5�<#�B�x��<�|�˼�n+=��
����<����	��)d�����a�:���@�Z��<BL&<�g3�4�e�X3=��z;O����_�!����c���k�<25\�J�J=�����e�<(�ؼ�A	���Q<|�C=�}�<4U;��l=��I�%�C=�u����=�r;nY��i���P_<��<#cz=��<\b�<I��<[���=��j�%�3=�x�<��/=�B4=�J�Y�1=�E=�ku������3����<+�t���<%b0=!����>��]���;#2���g�*:5=#���ҏ��0��;[(����<�3�����:�҃=��U�[�=�b���~��D�<&�k=mW=�D��Q��}�#�y7
=���<OHe=n��Ų�:q��;FX���&�C��5���v,��A=J=	�]�K蜼�Qn�7�%=Ն:=�^�����<��<U�<i�ѼΙ�< m�J����r�<��<���<T��P���=�/���b=@�K��UY=�=�m=��<=[邼�4	��lͼ4
����<�we<�O��q�<x(�<w	X���<�3ȼՎ��[�;�Y���N!=W⼘H)=�F����=���8.<ӒJ=���<H2j<V���X�`��2�<S����G�����=��<2靼�S�:���<nҋ���&=4�[<m0�<�I�lɾ�ؑ|��C�<@��<���<�R�� �<�=G��<�2�
��<�ǂ�LR =�	�;͜c�]&=�;K=4(m=r/��9�o���3˼A}�<(
�<�4�O<�8I��O��cg7=G''�l��<�qz<�u+��\=I!�Ը@���A=S�H={�;�[���9=�;�A}=~0;�jy�;ެ=�>�m�̺\����>�+*r���F=X�$��}�<���Bc����<S��<��;�G4�AP��r��K<�����`?4=�i<su^=��A��.?=�(������|Ѽ���<���<�C�:G=P�+<�҂==|������<�!o�4p�^N��O��<i�)=zs=�ȩ<�`>�$o���<]Y�;�Mj��=I�b=rѠ��p��;:<�Q����Y<�4����E?����'`==@K��^p�@�.<Q��l~n=�]h�){=�_=s�=�~���:=�$;�:S=����L�IY�7xG=Ǆ=IF����,���
����q�*��Ӽ�c=����Ԭ�����5��5�����;@4<�o��v�<�7�������Y=���<)2=3n=���<TZۻ���<�h���=��;�S����&�<>��/����C����<W�F<Up=�=���H==o�c�F_�<O�;?v�<��=W'Y�Җ2=��S=*R���q]W����D�<G�ݼ��2=���;IF+��1� :¼��%=��A=�& ��Z��`M=y��<?_<8}B=z����=�t�<>~M<�a��G�;r��<���;!�=�!G�qE=��<�"=軼bnh������{*��4=WZ���d:<�=��6=ܖH=3k1��O�=<�,�\{=5mټ$����N��o<�zZ=X�<�=�o��gg�փ�<E�Y#�(��z	;A��<fƶ<J��sC=$+:�� I��e�Y����:z�vrH����<���<����.=��)�?{	=��<���i��B=���tZ�;Vɼ4�/=��+��F��L�a����:�M��d�x;lC$��{�<�
м&I5<���<a�m=���:�u�<XZ`�Z�<�:=�sۼ�2o�h5���ݻtHȼ��<�N4�ؔ= k)�lyV;)?#;pP=-�<R�=���<J�b=!w�<�༻u����QS��y4=��P�d!T<o�<M6��V�:,A=��<��y<ysI��X=,���x�=){�1=L'�'�8=�	�ٻF==M�u����<a=z���1=g<�+k:�T�W�����2=;��;8��,ռ	�<:d���b�Gb�<z U�B�=LIC�E��<u��ق<��r�4�<��]������<���<��!=��@=�A�E:Yj;���@SѼ��	��ɼ�ɼ�f<={����;���<H�=��2<����=�S8�<�ʼYI)�%�=�>=�9_�T�T=T�^=��==D�����#�:��R��<�J�(∽ '=��	���=��7=��<v��;���3�r<R0B=�+<�y�<[F������Е�RW#�R[��_�<�GT=
����
<�f�<{.���żnм��=�=�� =�b\��BE=A�2��.����M=GKZ����;�����BE<��N�G/k= �ʻ��&��8���	�?1=�B:=�S�<���8!�<HG�<�0/=V+��(e��u�<��H���f�:�P=a6i��;�<��z��<<'<8V�;W���#=
(<B�=?�<���ḙ<�6 <O�J�5da�;x���*�s��\x���Ի�gk=��/���ּ�ּ�E����"=b0!�jPE=}�L=���g�[=$��;ȸ<�>L�V�J=�d%�'�=�������9���.�<~�=u2�<�>B=r�=�E�U�\�m���]kѼ�Rͼ�i�;��+�@%=<W�<�}=��9=�����<�:A���c�;��s�<v�μ�\��a=�	r=��!<�E5���v��1�;?¾�铂<�2=��;<��ּ�IT=V�=T�伤�`=����1tr��e���G=U�,=��%<�4�;��q�|pV=��e�t��=�<o�=��<�~=7���M&���ּJ=6�*��ч=9D�� �<�<�
�<%�������=Wm�[xm��s=��=IA)�"S��U=EeU=4�x=��P=}S��<V�<=��໐��<��û��|=M\��&���=��[<9��=���;��2=w���ǅ<D�����= ,+���
=&V�C�:��{�WQ��ֺ$�s����l7�<�U�=K�A=K=��f�Y���5=�u\<WFL���<��Ǆ��a~��=�=뼵p=�O=���;��>�G�U���{���q�����<���<���<`�f=4�\=�� ���ȼ��Rgj��]=U�=����ֺI=}0��A���=y�X=DC<�d=������<=�Ѽ�7;�>\�!�k<.2w<�L%��������~��<��/<��Tn3�mV$=�O ���:ձ=�t<N�$=x(G���=c%=mx�������P�ϼԱ@=-U=hV�<���</�!<�=��<�V��s.< �.��1<1T;�*H=Ɓv��� =��}�-Y˼o�"=5.����_��;A�B���d�Dܫ;�w=�-�<RBM�o{��_8��T�=�}<�m˼�T==�l4�(�j�O|]<�����U�<���A��*J����Q=�yF=�l�\7s=�
=Kh�=� 9��(=�\;vr�<��>=p� �E	�<Q�L��2��#�<V�-�޻��==�<><4=��<;�\���l��@���==x�����=��-=_��|�����=��<�4�`W��;=�:�M�5=aWp=Ș =ף�<���$2=XW�<���=�:��%�<���<J�=�K�<Cu<+"��s="o��:��`��<��J�1E^=�_��;Ӽ7�=b��<V��8ya=��%<��);�`=s<$����<<@8=L;�A���F�� F=U�˼�q���˼�}�<P�*�7[i�2mȺ��ۼ����݆ɼc"����V�%����C=f�;='9��@C���ټ 5�;>��<�'�+"ͻ361=F�85�=��^����_nP���W��1S��W�_�%=w��<o�)��l�;��2<��A��%;=��<��W��_=�Xp��Zq<�/;�ˌּ�̄<-�ݻ��<��/��"� �T���;�!���f�<L�)=�66�82���?=��M��<d�=3��< �<���<_%�Y�<��<WJ������&�=]2=��
=M�#=DF,��A6�y(K�`��<�;�J��f�c95=�e �.���d����<!��<;�;� ��<*��5�	=���_�&��~�����<6�q�H�l<�=u:�&=�E6��ػ�D껺l,��P=[e9=��Z���6u��.!�;��<m]�<�\<�$�;HN����+=b�A<���:W�C�ّ�;��D<��y={�� �/�m=��3�y�C=�QE�3�3���;�y>=ug4��E���/�?n9=�.�<�'=F�<�����*��d��Iu�k�o=yl=�� �#�;=��<�Q�no�<͒;SN=��\�<V�-�F�=��S<�D=k�&�@́��pE���`=�0=�%P<���?�B8*�+��-2=�¼@B=�1Q=ހ6��^=�7=<^=��.���$�����a�;�`=��(=��5< �n:���B�缆�< �v=���:��0��� ���@=D��xI=P�лEK��Nu<�M�< !��l�`I{�d�5���.�i�<��Y�瞙����0
�#��u�ؼ�C;=� �������z��ɰC=~�b=�6I���q<�q"�����垢<a�-;��0�����"=��y=�~<d��i�~�W3<?č:�c�<;2�^�]<�4#�a)9=2C�u��^�={"��==Ǉg���;%Mj=�a����8;Y��Τ���=3t=�x_=�-��=}><V�,��Cڻ�@�C�ٻ�O��}��[�;��d=:U�<���U.7=V��C|7ϮB�>4<�,2��iB��!$����;����"e2<>"I='^F�������+�*=�^���}��C7���`�B�e�z#$��A�<�ؗ<��O����B��<N}K�A�ؼ�!�U����g]=y@,�I ���l;��X���ؼhp��adN��I��r}ռ�z\�����{Y��kB���	=���<�[�<�%���^��'��Um=<`M<��ټ��"<�6=
��%�BU���%=I=�@=���<��=�^7�@/�h)�<k����Q���ּ|� �0Ս��%z�<�S�y3=v�<���<��W��"<���<|>=��<>�<==���
W=+�]���q��
[�I|T<t���U=N��{<_����;��=��e<��.��;!Sٺg�[�w��<,�ɼJĥ���<�q=��7=S��;-ɤ��=U�'=��%���/=�ا��<�&��`A=P�w�;�@=�ub=I�}<�mܼ���<߇I=�,E���<�)5�&�����<T�	=��=�x�;��
�l�n=mp8=y�<��C��h,=�t�<�l�;���:�[=, ��'{=<�N�7�3�:=H���%����/$���1���=�Eo;�E�����8���d�BJ =�y=�9=��<���<�7z;.��<��&<l����<k�K�wU�M!7���d<_����d���$<�P7����'��i8X�H��<�y&��c/�r`�஡<�Q�<-�U=�b_�Z<���GＱv(=�� ��=}�
�oܝ��k_=\gh;t�����<�U��9�m<�8q��ִ<��s����<�۫�8#Լ��A=�_C<�q6�K�d<��A;��:�o�<�E|<�13�Z�=�=@! =ȵ$����<t�;q	<g���e7=D�=� <�pQ=��=v �=?:<�==����+ɦ�Ď�=������K&=9N��)Ԫ<�3=�'�<5H����1�^��5	5���<�j��%�;�W1��I=b��Iv��t�<L}P��<rH=޼ļ���<��<K��5i�< �%=��;=|$�uR�<���9�!����T<��=
LI�љ�Ur�<r�R=���l�_�Ap�<���;G���NF=�e���GӼ���<B��i��C<�g;�i�:Ɇ���[{=���;�n��⾼��;�M9�-��;!J�x���5�P=x	=�����2=̲�<E>�>�<��Y=���;Q��5��َ<���<��k=5�;���W��>ײ;*x	��>=�^�<�2ɼ�7=6R?��m<��!=�KE��l=r.���Y=6�ռL�.=�v���k�5x���<�_X�:�=�L�<qk
�+Ñ�<�ؼP�qB�:���q?�N��^a�`
<k��<�B���N=3�s��=�̼��=�m�$�#<���<W�� ƞ<�q��M0���/��=�W���0��� 2=G8X�<Bu<W���= =e�μ�\���R��hq<t�=��E�)�k<;�+=^���Z1=����;�E�<�``��M=�})��t����Q��D=��<���:��/;��;��<���<�Ѣ���=�Q=�X�+PP=��"�y^�<ʮ��*����E=��<aWʼ���<U�%<�1���F�ޅܼD�;3>��b@�L>�����=��]<dU;�k==��;��<�q�<�=L�$�v�h�dɻTDʻ0)/=UM��p<;�Z�(�DC�<�N'���/=1V����<H�"='E�:.�=C�G�$;9<td�<�ż�L����J�>=
P���ƻ�l�["3��]�<�_��"���c�<�3�	���\=�i�=f�:��g=Q�=S�c��R$=t���l������G<���/O1��zN=���۝�

=2�`��D��L<�I"��}K�u��ݔ<;��;q1^=�q�tJ�<��=΁H��_�K�л���8�=0�<��L�"L	<S%<~�a=���<,��\�<�Xr=}R*�R+i<�c�yO��x:�C~)=z�<"Y)=9f|=H2=`ӼBQ弌����=���b��>��f`��;<�+��_�<�~D���y�wVԼ��r%��W�K:=�TI��0=��+���)<�$;H�<xj�;�x����<S�<A�꺒� �� �<L�n<�G5�i�<���;� @=�7�<�CN=w�}�D=+���S��;ʈd��3���K=�v;Hk��i���ƻK't=�ʼ[�S6��JǼ�2ܼA=}��;P���C�ܠ<b-w<���<=ß����<��c=J�7=��x��ޣ�aK��.��ջ<��Z<?�,=F�u�ME`�~�I�S��<�L<�Я;U�}�H�!�d�`��vr��F�&��;Z=�{ ��'%���ż̎m���1=��<��<�!<hI=-S缑�U=!�I���a���<[�1� ��z>�r�~�&��	f1<�9=�u<њ<��Ǽ(%=�x�<��M���T=��;w�;q��<J�!=�����oY��%2=�>=WBV����;mb�{񏼴>�OS�<���v\=,n`�$��<0~�<s��Ըu�]�S<�e�I�2��I1=���j����5<�vU<��:=��Ǽ����wP���{l=ˑＴ䢼�������Hϼ�9��O�[�'�F�W<��̼���<��G�`�Z=�@=68=��h��"F�U�L�Vݛ�jP����!=�䠺V:/�d��K�*��0X=ޚ>��)u�yX���!�;-��購�����F=_�0=d���Iϼ��<o�(�ʷ�<	O�<�k���Q��q=�<�����6���<I��2�^=~�<J�h<��)���K��eJ|�(�̼J��;m=���;�En<ې����i��f�o��D%�����l��2G<Z�����<�����==X���v	V=4!�<15h<��\: �$=�żv�ʼ��"�.��<��I�s��ڍ��HME=��f�*��'%2��ȯ����=	B'=�>K�"9���=�h���Cɼ��<r=K
r�M���T���L0ּJ9p;p:�1�9�)W�"c9�nCK<�u��R �qԼⷔ<܉;=��!�z)=9;
<
d=m�<�y�<�����_�f3E���6�,�����;����m�+�u�<.��AU<t>�;:�=2T;�.^=����� PN=��D=�<A�j"u�~�<#?q< ��3g�S���U������=���<���P=1
лq*;o���;=l8=�jּ) ��)�*=�v��P�#��o�<�Z�0'?��b�<�K[�) D��+=�N_��v��]47�p�<�pO=�p<g��L��0��<��;=�Ό�B��<񭖻��<�ͼ�NR�
��<smf;&�:n�=��	=��_=�N�����k����I��R=KN�E�=(n��,,�$^��W=Lb"=�yC=┼�t�;�3^�wW}������,�kR�<�ƣ�)�<7�8�*��<z�*=�M�9-\����:�i-=��┼�H)��@$��
<���O*��&���b�Yxl<�S���F�x��<��V=V�F<1�=�S=�Y���<�%��!H\:wWg���
��\=���<�rE��x:=R+=A^��\�<��+=c��<޹����T�\�2�}�ҼF�=ޏ:��]<���F@=�M�;EC5=^bؼɮ��?�W=��5�Y��<�<}�1=��p=�c�<�<1��<K�M���;�Z�<�)=ӆI=���<�~%<lV�;�����g�;P[�:V.;�{�=��<(9\=�G=8D=/��<����O&=���/'��H
���dF5�@3=��:�ѕ��M=P�p�6�c���Y�<���^q=�F�<��%�^����;Pj'<]=&W=M0=�9��Ʉ<���<ڠH=����*����>",=���<g���z�J=�د����;�Ȋ<��<�H���0�<z������8.=����w4��nѼ�"ʼ��W=�������7�M#=��ԼK��' �9��<;핆����2"=���<SP���%+<aW���_������ܧ*�Pa3�eT=����J=��r�q�2=A����T�K�H���<�ꉽ��g;��,=������;�m�;��<��J;;��W�v���<̞o��+=>�=�R*�<��g����4�?2�+ B=��<��=�D ��OC=䘓<p���|�¼��%���~s<�	f=odi=X�;��������
ϼ�y=�pk<s%��8=����=^��6U<L�F=eM=
F�<a��#u=ɀ<hY��
8�V| ;�?ƼmW	:jF�:ic=��=<ړ=I1�<u2���#r=Z�.<�j�����}��=��˺�k��c0= s;���<�+�<!�����<9���z���"=$'!;/�E=|�޼����ӳ��f�E�b=q �x00��]=|J��c=���;%�=�	=�N]������;��<�"=��<��� w����<k�-��h���Ȼ��<��r<c=���<{ �=�i6=�$M�5Q�4X<w{������c���";���<4�i<���95mt=���Ï=����Fۼ�؃<Rc=����o�ؼb���p�(�/��j;��ś;��'��p���<���<��"������:=�;�-��W=.��<4��;vX�wK<�b,=||�����
d�;bR��	�=�tV���C��y���:�Μ����=Zh�<Y�J=�<�<��+=�[�W*�<:R����3��<�KI��¼Io�=��<Ri�<�#���}<��0=FEi�?�ü��r<p�|�</��<w=��	=�+&=?��<��p:i���^�X�b0I������8��N�����=+��<���<��4=��F;1�-�KX7=�)=i =A�<5Q����Z�^=VQo��3�;�J�<��,<΃�<�j'=�p� =�� =�u�<�U^�ƛ���<�����p���[��׻�	�:l�<k�=Al=��@��sE��O������^� ���%�'�B��g�� ��'Qa<���<He#����;��D=J�/�_<"=+����Yi���=���=��>=B��X!Q=m=t��%�D���=�H=��6=+w4=���$;=U{�<�]V�Z
j��h�;��{��/�+�/=K�<;J�d=��=������@=I7;=���<��b<(��;�o�@^����< �=v`=�^j�����<�&<s�˼�ڡ��*�;E.��?�Q=T>�<<>�+�6o
��NW�hz��<�с=���Ͼ-�G=&��<�o�<KK=f���J;P��м�;5d==�O��Svv���}<9���#�*[6<8Q�<;q�<����(���;�=<v�<XC=^�y<`<K�d�>�<T�0=W�.<�G=;�<i��&8=�ԍ<_c��'1<I�'���+�
s��t8��`<@Wȼ�L�;V�F=�z;��P�z7?=�2:�9h�:�==	Z���S�sB�;(��<X�j;I�<�OR<O���r�<�<��i=��=�,���ߺ��<��3=���� =
�ݼ����b;.�ļ��U=$�:�J��e^D=*QϼO=��u=��<5���%0=LJ)�����W�U=��F��ײ�0�;@d�A,��bn<+qz<rՎ<�Id=v13=geY�J�;`�<����@#=E�;�*���<'��˘O=,,�<[�U=�=���N=F�<�_�w<{�==`q���С<�t�< ϼa�E=�=;�o����f1&=�R黶��AK��l�=��߼�NA����-�� v�o6�<�EG<��%<��)=t�����$�<1��}I=% s�A��#�f�y�%=��"�P��:e|��d��m|-��D=��;�!0��wK=�M�<"4,�=�;V��<P�m�R�5=Y��;�!ü�$=�}Y<:t=��+�L�<:�=d�=�W� ��Ѕ��|'��M=�M3�y��</�$:	/'�a����9�,�ۼ�� =�Է;�k�6����o�q��j=H��<�z=�(
=�
=ۺr�*�&=S0�;�=ƹ��{�AJ��b� =�p�=�'�ڒ%=��<^W�<�,k����<�QC<
g[�
�"=�Z����:h�i=2x㼓�P��y;���<�ʲ;iS�MK=Ǫ*=D=�_R��'����:{=Q��<�S*=<0W�	S���˼[t��͔�;�]=���$D�\�D���c��d�k7�;:�	=�?�I4�x� ��	�w?1�"(<�����S�| l�Ba��}d�t�=QI�0G.�9N���q�c�G<sMx<j^�<-=C�w<��ڼҺD�'��<��U�t���м)�C=��Ȼs�?�2$��="A�ܙI��Ns=�|P�%#��k꼐4-�7�>��I��ߵ�:j�;@(<=7��<�;S=�;3�'5|=b����B=�W����<*���7�"=��O�7� ��[�D�.=7C�;��f:2��;i�T���G���N<g�$���^:T�}<	=�N<I��<�p�<�ü�|-=SC
=�"s:�\ �$]=-Mm��m=��<<|,=���aI;�nD�\9�;��<���j�R�TyW; 6��%=�nH;���mм��
}ļ_X=��<3~D<=mW�<�Ӽbw��nkX=�Q<��ݻLP���,��X�<��B=���u�=�X�<R�==�� =X��!=[<�m;�]q<�Z�<35��i�	=�����1=�"}=�J=Ӂ<=﹪��ǒ<����=��=�B^<���˚�<~	�Z~z<%�i� ��
dv�n�=V�<n�<X=7#z<��<��缋�<�:���L<��4=�1��Q=3�=)f6=\�B�h�=�]�<h��<-�"�"�=�I�=�]Z<�>��53��
�<S��<�V�<��D���i<�7��G��Y���z�<��=�Z�<�0�<�&=L�\=cڕ<?~*=9��<ڠ�<�`G=N|�)��<O8�<��<�S꼹�g=�{F=�S�9gH���R=�PK=4:�����L(�9%�-=��A�:Y�]Ƌ;j8H=S�GX��\�S=h]��z<=�5i=z�G�㼆���킽:+��}a������$=R���x�N=%ё� ż#�;��r��Y׼��,=�����=a:�:�Oj=������<.�=��F=�2������:�<h�=&����8Xx�Wrx�N!߼�v�<	h�<$�h��2!='CH=��)��YO�Ҹ
=R��;��c=ك��h6o<:B����<f.V�����ZX�~�=��_=��»��N<�/=�4=��v<�#o���=�+K�)�!�2�żE<��\=@h��r=��8�q/2�M�<Un���W��?4O�t.W7��
�����Dn��=X&�;.1<rL/���=ٱ��NbY=?=�z�<v�C�)F<=[+̼��[���<��D�D�+=s��<N#��D�";��=�@׼Vg���~a�ȧ*�w|�;��[D{�J?�p�=�+�<�֠��`�3�ռCB�<���<��!�O���s�����w<���<].ۼ�7k<_�ȼ(R\�)��6r���?;=�?��:B��<I=[co<��2=�s�;B-��v1<c�!��m�;�~�;��ͼv�O=�F�<�#��]�`;�z=�Ǵ��=U\=�A�<�m4��\���ER=�[t�e�����vi=zO[=C�a��a����<<�*="�=���L=�����<�`9=K,�:!�7�~<o ��V櫺􊮺-�ּ����,Y =�L<�)k�
L<�H7;��k��]j=��=���x�׼�.�<.��;�<�7���<8���E7=h.b=�;���=��Ѽ<;a�p�j�96��螽_F�:;������0�A=��=�=KFJ��}�*d����j�л}�kżѹ��C�ִb�E��;#��<�U=��Z��VC=�o=�����3=�<�����v={�1=D��<�
�<�1�;���۵<������:�SD=��=1���Gl�;�Q�"�=1{�=Ӏ��=]s=�i�������;,Z¼��=���<�m��\=�V3:N��;[.��O�<l==!�<6� t-<:�=�9��G���P�)�m�i���s�,��?�1�>B<:7�������;�}O��%K��L*���뼑nܺh}�<W��<Der���=�Vx����=bfܼ�Z�<b�\=�s�<���a;���-=� 1=�Q��{<A�=�,�<U�N<Q6��Qj<�&=��<t&=�7�;
�<�I<�<M=��U=��H=m�t<����"=��<(D(�}��^�6r�<�����e��5�l=t����Ȁ:��ɼ���������<ػ<��켍;$�H��%=�G;�d���]�@�u��2�<ɚ��j�ܼ�i@=*x<��X=�|K=��:�籞<�U�\����(�;�.Z���<���<�u�)��4{���G<�Ӻ�w;jr �opn=�ߜ;��F��0g����t~�<h+F���=am�� A=j�;�h<ˠ�<o�����ɉ��ܐ<D!::�9��!���»<��S=a�<>:a<�`�;�� �.9~<�� <��6��4���껹Y�NS5=k�4=5'=��aX�/��<0�(��k1=���<��'�R4�<�����<�r=0J]<KN5�~<`�t�I=A�b�R��<'��<cI@=b;=��<��c8����<+[��A�������hC<�B=1f������^���2<gO����P�@��.�R���ϼCK�x�=���<�!���/<FSL=�&'��l���+�<BJ���<[�C�*�j�g#G�^�L�"&<�Q|=� _���N;�+�<��Ǽ:Y=��b�|�9��+W=�D�;�$�FP|=�g�<W5
=�'���@�]�=x$!���7<��;v�;=�Q=a[==s5�=�S��<=׻�q������_�)�<�<�}0�ü�k p���l=��)��]�<�;�<1�=�`�ս�<�}�;��O=��fb���4=Д�����Af�<^s	�n)=�1
��㵼��$��=��=C\�;��^���_=��S=b~��iIm�:x=�om<��WhD<W<���1��Z��s����<�?=�t�Tb�<T�8<s�B<�fɻ+�=YA�<罌<�YѼ�j���D�\�m���;:��2Լ;<=aI=�7<=`6�<z����]�=]���@=1�Z��A��|A=ӭ���޼�A��s!�:jI<_w��=o�M=�k=�.���Ζ<Mv[��`�<(AN;��i=�����<�a�<`|=j�c�.=+��2FP<]�:c =��<7�����1�/�żB��<�����-���LX�Z��<w�:�`<,�Լ��弘96���<"�o=��	��l=��6=�̼tH=w�<�J=�p�(�;Ļ�<�aF=��n=����`����k1��~�<�����ʻn:=�rE=Ў=0=��̼
o��C"<Z��|���ɱ]�I3m��lͼw�<��=(ʫ���2�pȏ��ˬ��"+��4d=�I\=t�;|�?=Z�V���F=�b��(��嬌��=����ܿ<��=�%"�j)"=��;��T=e���*�<�5���<`�O�MI�ب=J��<��s���K�E,��$�l.F=|���Q�=��<�>�⺃i���e���I��M�:�r����=�$��*WA=~���!=
��8<�<ݙ}���+�{\='Y4��=�?@= �=n$�Ou�Z>��� =���<;L�<.k���q�<A�H��=@�A=]-�Ʀ�<�u��6�";,�"=��U��Z=��#�w�#�	&x=�� ={�}�)Tg=E�t<!�<-�s���:<�~��܁<,~E<�"<�x<K����<4�H��#!�0�a������޼�U�=�U<�*���?x=�sS=��=�x�<�6I=Z��<[(C��Z�h�`<f	��OK�h�6�+�d�;�A"���<�N=��㼀Q=�҅��%�����;��8��'����L�2=���tݼƼ<}޼;q*=���<�G�<CH��Jo\<�gy<�f����;��/���=p���z-�6��:�<ݼ���<�꼓G�<m����h~Z��1=\�#��6.<��}�H��J�<-&h<�ힼm�ܻ���:;!=�!��������<4��b�������3<<`V��\,�YN%�s�{;��.�2�4=�pt=TRI����<�~k��]G;�2z=c��]f=}��uRؼ�(<;��	=1�Pa��w=� =x7Q='��!�?�y��<rm�<��r�dv׼��z�.=����V=(=��0����<ѝ<^/�:���d�*OU=4j����L�o	��;��)o=D,	=,�L�7劼�By<V8p<��<<��<_Q��9f=�4;=cH=4K�<cm�H$/�"���8=yn�<�:K=��;�V9���@=�*��H}�<}����Y���A��É�e
?;�^<��D=v�T=�h�k�q<>#�<�����Y"�\D=i-�<�v�=-a2�|�L���=*�<$'<<�Q��dR=e�M=N�=؁,�Mi\;��<����͠J<��ۼ��g;��=h�=̾��췫�ZJ=��ջX��J�5=��<�Q�<Z�&������*/��F�]3�<�V2<O��\W�:v�=�=��a=G�R<��;C\���KV<��*<,\��V߼��#=]U�<�W�:�4"������X��{�BWy=��+L�q���n�Z�<�A�Ma��r�c�	�"� ����Ay�w���??<�ͷ�dvA=�*k��N �b%���u�����4X===��!����<�Z<)IM���ճg=�l=ci��<�_����<��a<�j?=zf��4=/�<�K<J�[;���<y�1��R=of���`���A���"���=F��~ڮ�������<��P���;<���E.��) =L�V<��N�U?����n��<>2��-�5�كɻ�}���G^�$A>��$ӺK��q�;�%&��/"=ǾA��#�=�P=�r'�ȭ�ҮH�DGa=��cY���'B=�p$=��g�|�<��1�l���4(��<�:=��G=$D�<8(0=��6��!뼓{����6��K�m7���;��U��A�<z�=��=��4�<üsb��*u_=���<C
���3o;�#=t{3��x<�������<AR=��
=��o�d
�$��;�o=h��������q�<3	9=�= =�#���<~g<��=Bq�<?O=s�=��=
'�K�W��.�J����ǈ=��=�~ż�)=�T6=a�,�\HL;P�E=V��fp(���m�Ԁ;�4<$~2���a�M�^<���\|�"��<94�N�=�}>=�*���$�d=�)���&=�Sg�q[=�,6=9)�<�8.<�=�?=9�����O=GT��Y�`uN��l��,>��S;�W@L<�;�[��5�a�<�S%�� �+2���C�����Y�:���Y�;�:��$7=ܾ�G�/=G]м����)0=�=E�;u-=��Y�l��if��Z|�8�9=*<�q����i��Q�;�ZY���\�<�9=隑;<݉��v5�%dX=�j�zd=�ڼ�U��\k�Rm;ט���Y�T�B�&LB=�Fe=��<�K�;z�v�k�0�/�9<�^�%M,���N��y��
SL;)�_ټ�<��4��?%\��݀<R��s�=�{<���>�;�<�<g��;�-E�=�h=��0={��D^�G�<4A��u]E=��a=�/7<�i����<$k4�-\l=ʔ�;2�[�y����)�<PI���C���N�;1��֙<�H=������S=�[=t�P<OL�������#�������䧀;?�=��<%R<Ro����&�LQ��IH�����,�\<:���P�Ы�V���󬺋��<#�ͼ����<J��<�+�;�!=?_<^k�<��N�i�`�2ly�j܄<h�V&=��7�#��S�)=2;z=���} =�#W=�q=2F�_��<	��<\�.<N�S=�6��Vl���J�``�<�+L����<4��<�<\V�<^!<�,�<�Z�<|,��\p=�N���1�< nW�%j�<駦�hr�<5Լ�OQ��s)�$@=E}޼(�A<���I��:�'@=.5=2�;�iV��� �`|���Є�@/3� D5=|���~� <F�5k=WR�Qo=ߐ����U��G�<�''=��A�<��<������AZ�<���<�=
�ƻ�c<ԁ�<�V�</����<�cd��.0���X7=�T0�8�J��1�<��ݼ�!�p�=5@T=C�<�5�;�߽��_=��e=c�X��&-�3a�;�xF�tؽ<�@�<���<B���K� A�<w/�<Վü�����Z�k�	=��s=�u<�24j�M"ݼh��r�;�R�6�g��cu�< Z��:���<��F���ټ��<E�<�*���C =�M�<��<��E�P���6p�N���^��=2���N=�w�;��9�:=����*�C'��S�ɺ�EżA�H=(�=��̕;�i�\�;=��n=�c�I@;�!ܻZG5�\ �A�<�=Hx��bD��0��1=|�"�ma�<9%a=8˖<�P�;f�?�x�~��#U�V}]=�@&��F��&ʼ<��q<M�%��:=�C���̂=y�׻�J:��y�<�H��Ζs�\O��Ao<Y���`��{<�ǻC�=��G=�j=���"=z�r�"b+<�)T�U�<�B����ky��ެ��h�=��=L�1~��=ߛ�<�^=nu¼�����-M=�̼�	x�#�+=ؕ=�t���l�{�G���x=�x���f=]_=HV�=\:=<ʮ���!<�'<0�(=�w��n#=�*�<���m>=��-��P�o3��!>C��iW=�D����<�n�=���O�#=��ɼp�P=���UR�Á��=�f�,��/��V=�"=88�#p7=��%=̪���r<�L=t���4��}"ݼ;��;�=���W#d��m3�?�J��F	�Y(;�a����<��:e*S=D<=蝯< ץ�ۛ$��=��D=pͪ����p��{�Y=���;+��b7�ۚ"�b�X<b2�<�uy;��5;4�]�W������<����_&r=v�*=;b�<��
����QU;��).<�L��ͼZDo��?[<l/B���:6nE=w,=�� <�?����<]l)��8�;M{ռ�!=z�*�+}Q=�<e�2=���<pz%��]]���ͼ�H��,]�<���;����<]�@;����7*=��"=��=�*~L���h=�	�<��0�4N;pżt�<�=���K���2�<��к�)]<��"=�̊=�H��2	�k�
=��-<�7X���=3�8=�x1=H%����<O{�<�7;=�-�;7CF��'��>=�����q�n�<kAE=k��<�B�<�iJ=%5=�� �\S<GxJ=�\(=�)4�:��(�N�it��b;�Nһ�~.=A��fV켊�<�=g���p���UX=r`�<�q"=G
\�[�:�X��Cr��A+<�6h�$�ż,u�����<%�޼3'Ϲ`���Hڻ�>�唼�ۛ<�+�V�8�C������ۼ)y5���0=����$/.=�/|=��;��U��==^�<*�<
\<���~�����Rٻ��=��<Y���f5=�`Z���׻�)O��.]=5��<��c���=�)��I���J=m�[=��=kk�r#�0�ϼS��<�Ӑ:`��B.�<Ӻ(�/�<R�	Ne=��2?���x=��!<a��\==��y=�6��^=6�=���;5r��eZ����
=��`���;�Ｑ���E���+�#��Z=ZKV�@x=��H<���<��Z�5��p=�m2�����Հ�^0=�푺<*_��U��<��<�����:҇N��6=.{=��<�cۻx���V�<\�9>����g';�+N�$ބ<l��<��3��Z�1櫺��6 5=eY}�8h8�eR��S���C<r�<�WW�W�l�8���-�c��f]���<8Cz��S�<S)=S�(��`K=)%�pI�';}�{<�<���+F���ռ�x�=�΅<,߻���mV9=;�o���H��"o<��==A��<(�޼���8 ��"�>��B1�9\4=�c,���<?`t��
6�x�2=œ�;3d���Q׼��,l�;_��<X;�$;=���=�(v�?|�#!==l =�@�<�`u���˼��Ǽ\�</hR��Lv<2����,(�M�<��<[��<�[����Ƽ_M�9��;��<x�<�!�1�XR;'��<F�_��<@���R7�]+�p�����/���@����;�� �(i=`�<A@�5�I<q)=�@d=+8���O=d;ڼ���c¼�(5���;k�<�L���<�1=�2;�"���!9<b�z�
�=,.�;�
�<�.o��`�<��(=7y載:��a=�<�yI�����A�$��1�ܧ=�j�K��B�<٥E=�r=���ن3=�6=װ����C�u<�V:="b�<; e=��<�=�h$��#/�����ˣ<�1���޻r"<S[=�x=�\�;��<�)t<J�[;�u<�'I�Yt�����H�L<bDW=�`�<���<ះ<L�0������D޼��f��F.=�n=���;���;e�*=��=R�==�mo<��
�7��)�+=3+={�w��w�߂��+*3������k���p�-�{�I��@qR=XzJ��c#=^��<��/=st��x���@��a7g<� =<Ų<�꼼,�;��d=��мf�k�Vs{� 񏼻zg<CY�T$<#Q<8��<=���ʼ	Ѽ8�v;���<t2Z;���!';OC�m��<r������=eZ�T��nݎ�i����1�<���ae=��;ݪ�}F�蓪��������"�e��<��.��g��/˿�ku<���<p���u��90=���B�W�X�]�h��$�T�U0�OJ�������<x�D��JI=4����� u=���<5�<�o��8��2 ��0����<϶���M�W!�]��<ں ��%𼉪=�o�[=�v\��M�9��"=�Ou�s"�<�=��!�v��=��ἃ�=��ʼ/=�O��5J<]YR=,o�_��;׼�gM���J�+�<=H`=?~<T�S���(�s�=���<��'�+�@�%$�;�&=%ѭ<�0=jڽ���=���sc�Eh�<�lj=��j�~�O=��<DM��j��	�Լ��J<���<\#�{LN<ʆH���g����<s�<��=�T���<�_�<c�7=v��;��������(���9�#��<�x;<5�ݻ�s�=�c<�ޮ<��<�<i�$�̂Q�:���H�����z=�����RB����<��`=aễ��;d���P=�~h<��M=HZ�9b�H�l�G��$[=�F=�%�<��7��4<s�8��<�I=`ⅼ�-�{ d=�z�<��T=���<��7��Yo�r�<���F�s=tAd=�!�<Zü�2K�k�»�C��'���Xl�<:����*���O=��0=v�b�0z'=�\;�]�<�,�<�;0=Z��{j=	�ܼt`	=�^A=a�)=�#����/=߇_���,=z&=���:�V=��n��X=2�)�0cw��d��T�<������<_(R��7H<�n��]}+�P=�o8=Xy���Y�5�=P�#=��輕����x��˺<U�1=��<A�	�	r���;�(��9=л�<$l<!(����q=r�*���(��h#��޼K����B�6�=�O�<�p�ׅ-=���pg'=�r��	���� =��;�h=�7<Ò޼�)�=���*��6Œ�S&P���>;�%^=�g=�	#��+��Ϥ�!Qz�av;��2=�ؐ<*�)�m�W���i�C���G�m으���<K|*��l���<����b���=�)۶<��<�2�	φ=�FU���=0=�h��}���뼶����F;��^�pD�q�L<?�=�~l��<R�<p�e=�I�ړ��50=�ڹ��L��<�OK=J:v�D�ʼ�h$�3�O=��;�F��!���Wռ�N=<�?<�B��,k@=�(=ES��z'=@;<pr=0��<i1�<9�i<Wm���D���6=��s=�7Y=	���2�Moc=�G����<+漅"=T�r�>#�;җ<jTa�Ҭ�<��1���<3��<W��<��;<)#���񻳎u=�t<=��<���=L��<�=_T0=M���
d<u��̼�>�<���<�)ݼ��<a
T;��<ǚ�=�>W=�J�\Y��1(<�=��<��	��q=�����pk=��9;-ȥ<^�M=�9��<4�o�H=p���9&���p<��k���P���0��db���׼f�>=�XU<�����7�0=8o��<���ky�4��;�#��G�=�3�ϐ	��bZ���=�2L=yWټR�;=P׊<5t<�⾻љ<b�;�Q=��=��h;�C� ��#���F=m���<�%Z;�.=�S
<��ռO��<�=O�#̬<�W�X�<1�=���۝=��μ���1��<T=k<@��)�<`������5<�ͤ<�H\�*�=��l=l=���=���<�:�;�T�Jy=ba?=2�<��=�]=Ӝ�;-�ټ8�i�aT=4���IO�zjU=�.=��4�Od����=��=��G)M=U8'��}'<7V˼�=ټO�H;�<��M;%d=V���(H�<�Xk�ꅼ�%b=��D=+1���(=[t=�,�G����#==�W���	=�p�<�J�<�R>=�^;vc!���:�G=����/����=�@�<���;tm�<�_��|s��<=u+�a�H�Qr6<�l<��V=`����Pe<���<L������4%=`�`=��N��+=��2�Ca�bD,���s=�=P��;�o�;+%��6��<�X<�b�������`��l��=d7ռ�������<���;��q<�W����A=�8#���J=����D�-=�ȓ��'B=2����)���fb��WQ=��y�`= !�5�=u��pܼ�݁=:A�TX�j��G�0��x<F59�k<���<��L��=H�^�@k2��N�;���5�?���m�{"��F<�r�<�����ʼJ�e���>�MY��Q��f�$����;��<���;]}�
�q�ռ�?Q������0=/Ò�cv�6W�� ���2�n;F� �v��:
�;�e�=3H<�m�<6F���&E<�e�;ܼ_<��<y �sY#=r��ޔ��������2�K"��=%=�ۓ���４�Q9�K��Y7�4T��\/��g�<�=�u��"�I=��3=�"1������� ����K�=<D�<4=
���}yJ=n�==}�b<ˏ7�AS���	F��+�Y<�
=*�Uo����"�-�U��m;�=}��=��?<�9N��t>��V-=�u��D=��4�e�Y�ئ\�\UX�2�b<񊲼��=�^�<��A<
d���Fq=�J���[�<������H�^�B	⼊a��}k�<�Լ�L�Md�<Un���~=��
�BSջ'[һ@�K=Ky=�_>���!=1��<�y.=E�;�37���=�c�;��<>/4=�8Z�Ό�<����!_;����ה?<3�b��W-=���<g	J�N�v<�r���+��ټ���<ԗk��T�������	��<+�;�5H�z]1��{���$=V��<I�G=���s,�f�<������=
Ԑ��I�<Ӂ�<�B�9��<�z=֪뼚�&����<���8V��%E�鰘<Jq�����< d��v�&���ػ�Q��9E�'�<%�<ZT^=��<�a=RBg�;��<�j�"=�=�G�}�Ӽ��=9`;��)��XN==v,=W����9S��_y4=��V�R����@;`����[��	�:<�̚<������;^��T	=�MD�j,=hX<���#��=�P���n+���0�Ǧ�<�n�Q�A<�'=��A=Α`�|m1=��:��V=�#l=�2<��Q=A��<3�6���)=%�\=���fW=���<p]�
�<� ��d����Q=-�;�(Y=#ټ>��g�9=�=q���P��["=�;�C�-�ӝm�meH=B�=_q0=W�ļ��M=aټ+�;��%��1༧����:��h��<��U=Lꝺ�,�;���!!����D=�U=쐂;M�o=5/���%�<�r�<ļ6=��Z?�<��S= �����ջ�S��7_=�%O�m�:X�=W��L�R��R��<�s<*��=`~��F�Ֆ�;v;�v0<Ux=| ��+���;K�`=��j���n���O�
�4=��<2姼M8:�\j���9J�T����TW<�Eb=n�=#�=��;��+=ư_=�� =��F�^��D����.;`f<a�����<jU�GQ<��\=}@<H�������"�v$<���<�L@�.�伍f�<�?c<*�c�'���G4��u=�r��(�Xh ��G
=�=<<5Ӄ��G�>�;�a�jj6�O=�J2����<��9��<��6=hG��M���A���t)�A[�;��\����<x%�$ <�=?<G���3����;�+=�~�B�G= 11� X>��4=�2
=�	|����伿���~=��^=���<���<�dU=8�-=�m%�:�q;��%��k���C��:5�I<#�O��x8�qy1��:��:c>��'���=��%�o��7-���d<?BZ=eי:�Ǽ��9��[�$�<��2=�3;=��O=�gܼ(;�l6=�c���V�<+����`�#1"=�
���y-�ztW;����ʻ�#F<�UK<�s��}�;��<���������,��MƻSDK��=�I|��{^=��n;�S�s=t�0��]�z�C�0�#=��,�t�������D<W�C�-t(=G�_������<T
K<�=�+=��<�ZG=7��;m/%=2����;G�A7�[(c=���<�ӻ<0��zs�<��'<�c���ϭ<���<O��<���e]=m�R�Fe=&�4��	#�����[э�� �<��~;JK0��t<=�R=_vD�]>C�~!0�	��<�4f=�8Z=:��<l��o ڼ��<$�@���<�_=%�<��Ǽ#�
=\\;�[=�%$<�3= '�CK���9U� �<�c�v�|�i��<�\%������<�_�;�n=6��[LH<ql*:'4�<Q�d=�Q;=,�|<9�Ѹ:=�9��s��<DK���L��CO=r�;1)&=}�,��[�<E
=��<�h_�#������O[�afV��ln�v���}㻣�<�<;@���3�BW ��Q������j�<9�=�+@<T!~���<�)<�6IC=]�Q=5	q:��4=5lY=��L=�Ec����<�2���-=�ۼ�_�20��4�m:��SW���"���<����|'�j��<�.=.�=Q�2�iШ�f'<巳� "�a
�<8.E=���;V6u<?����y=��=�Ƽ�W&=��<��(�s���W⼥�[�w}�<�0��q�F��=#���qS�<l��<���<g�=��<T�v�O1�<�\=���<��l<�T2��1"=��-���G���,=�!��ؼ��=!�=��==|F6�C���%2<x�Z<vvF��R���I=ҭʼ!�＜��U��Q=(�4=b�c<v[����7�_ �:�=���;3�]=�^7�c������"~��ƃ=޹�a�<`(=ic,;�d��Jj��D=<�H��-�<�P?=��c���,����<� ����<��$=����a��'B<�Q�ؼ�8Fؼ�	}���==_?����=�K<�`ϼL�&<O*�<:�|<��y��~�<=�K=�M=g�q��<�;e�<(��<o�<rO]���޼u�=��<c�7�xب�T��<���<���<��D=�z�q8-��e�<ޤ�;�R������<�8:2oL� yR<��7=�<kHݼ?ʼw\=GټL�=-�):���<ge�3�ȼ�]��lZ=��W=�z�;�/�<��H�`��i?)��[)�Q$�<�@<��Uj�4�&�#b{=X�*=�gp��<G;�/���!��uK=�I�<�	><�<@���#缕I�<�*�<�v5<��(�G�L�h�<~h����=:�<���<k?}�N����;7�`�2�<���x<�'=�\>=/V=D��;ڢ0=O�=�OX=�=L��DB<���<^W=��=�E��?V=�Q=�H�N�(=og]�2l�<�м�8�;ѿ>:Q�;��H���;�j�;";�>AK�"G?��뮻��R=�*�<�mݼ�/<���<vB<Omt�&�=P��=sN=�q<k�<�8�OB���	=�ƼQ[�%N9=�Y=�4��>%=�'Q���<�sJ���;$�s���K=���<��s�KqV���6�I+</�
�_	#=��<ɋ9<�0+=�!��x����Q�ܤ=5�$���-��I�1�N���޼�$�<�=�m�<�>��d�<����9=/=�\ּ���<1�(=0�<���<����8=#5=�I���!��k�<){6=(<���,����<=��4;�dc�Lʳ<\�R����:K�����f;b/N�p)P=�J˻� �;�#��!��%|i9]L�.z�<�-�mV�9dH=@!/=s�<��Y���w��=�<��< ��ڛ<�W��+�/��<���<j	j��:+�[�<�/����=�$�)+z<q�*��!��M=;�.=�C=	վ<��o=��%=��A=�W=��d�[E�<�K�</�=|������<�.P�6g;RL=wި< ��<�	=0,:�X2f=�B�;%3�<��Y=��¼�Ӽ}O����>=�E.���~=�'���g�<s���0���f�<�<E� ���a��Ǭ90?�<D�<v(ҼDxH��򅼸�9;^Z�<r�I<b_��4���ҼZ[a��C='=�%��m������zԼ�v����<�W�$�U�=�9�w�f<�VF��iH=؅Y<)�D�5�<��>����<w�#=�_f=������=���<,�4�\
��n�V���<w�b��P�<�Ἲ��@=EF<��r=�/x<���%�=X�0�KJ=�<K<ʂG�D��^":Sݾ<-M�<%^��]�;��5=F<v��$ �?�%����<�'=R�<�al���W;2�Z��;=SUK����O�:&y��FE�;��;la'�[}#=��>=F�=jb�<��<;���6T�<�A1=�j==N=�i=d��+���ϼu�ݼD�ϩ�GȂ��	a=F�<���<r�X=~C=��: =�gJ=`�s<��s��d=�t=|�B<ʦ�<x��;B�<d"#=/bI�'� ���>�7�"����<ѩM=�w��D#=v�=3|a<����+C�ʼ�<�!=�`м�R���<>1<]!;��Q^=�{)��t=��<�g{1=��<�>�<�7B���Q�K��;��<V��<�J[�D�0�ya=YR��,=����b�ü��<'�<]u�<��M�$�U=� =�M＼�V=���.@/=bxȼ#���<2=R���K[=Z@�<�[�<'�!�;k��j=�k�<F��
�)2�,��;�뛼��;���<���<��
�0���\@�[�(<�nh;�+�;PZż:a��C�<eL�}L=@�R��iY=hPr��<<9��=��9�-=���<�a�ų,=}f��\{����<_�<2+;I����9<�'<,��;zۼ+��<�]ܼ6�%=#$���0=��7��D�h=/z�<l,#�n5�<��b< �=cb=@�=���M��7=�m#�0���^���`;<H�=� �c��<op��E)뼜�H�=�#=�,=*��O�E=�à;N�;&ၽ|QV�J#A<�-=;f<<�=�4��g=���<uV���mN�� =�i<;)<S��<5<9=G��~\p=K
&�Vrp�̜m���2<��T�-�=$�=��m=W+=4�l�� ���H��\=��<l�'�Z��)�<Z.k=N}��5'��W�<B%����n���%=��V�#P7��0U���}�!�<�}<��<��.�yq�<#�ܼ�;�b�=t��C��� �/;b�=���<pv=<��<������=ɹ/=�������%��J�Ǚ<&�=�<�q���<��-<�f��%�q�cH����ڼ0=��<�u7��_�<
�<}�J�Ab=6���Uc�a�C�c8<�k��;aJ�K9=�<Q����R�-==ȶ�<�E=ƞ�<J8<5A�(Q��R'�\����0=>Y��E~=�Y�j��,f3=�bռ���<t�T=+�=���<��<x6��ܥ����</�i=EJV�&Sf<L
;�#�&<,"�<�z�=�g����O������V��,��ߐ�:�=�*N=D��<J�5;�f<� /<���<��W��4���jV�T����t<kP�;&�&*2�O�޻A��;�����o��=�A)����<5P�<[�>�D�`�>w=���<.�X����<��=bY���~;5LĻZ�O<FB2<
�=$1�:�
G���< �#<�Ɠ;�9��.*=�&:<��o��Q��S=�`�=�3;z	m��I�<WJ^=3{�<5=V���D��<�6z=ps<��"��� �kq��K��K���=ş7=�3m=w��<.'�;�g9����<0YR�^�%���A<�;A�����5�:=堑=��\=D�
=���;$h=�BQ���=\����t=L�ż��p�<���<���mFP�5�_��~�$?����;ʀ	= y�;$8�:�=ۻI�<���a=�!*�n1<��3<��<�xk�/N��識X�+��~p<��:�5���,�z9�!���gI��lc��A���=��i<=�3�T�=��9=��y=�!3�l8^<�� <1�7=�M���<-z����p��_�-"��1U=8}�<Y���p�;W�=oY�>�3<���l6��`��0��=�C=[E��j=	�<*��;T�N���;��""㻫zм����#X8�A]�<|#G=��M�N�%=oZ��ȕ=�z켴?z=�D=��<�V��|�R<��<*ga�^")<�����j<|�(=��ڻ��:��ټF�L� ?�h��<��;�/-=�~=25Ҽ���;�,>=���<�0>�7=�)|J=�}X��d�fV7��|R=�Kb��be���e;�x��+fX��T�<�G&�͊�<F�b=/�\;�q9=���<==��U��X�<�I=���=�B�0�S=�V�pɣ<��=Bᇽ��w��V���ؼ(��0&^��^�����z�H;��=�Y���b;��#=7ҹ���=�ew=P\�;Vm<d�=��,=��_��I�����<6�a<&^"<�*�ۼ���"�=1S�<ΐ¼������j<�hJ=6:�<����8�7��3=%h�ۑ=�5��2=ԂQ���1=�[_��z6=B��<���<O==|b*==;5=aN�����w�O=T�~���8��%I��߯�n���w���O4=�Rݼ��<;$�P�#�k<>O��f��<��=�r<1������c�FaQ<M�X���M��ᨻ;�Z���e<@�j<T^!��v=N{w����F�M=C��<hV���<�h�<,Q��_	��w\�a|��ῐ<,d	<���i�^���]<��<���u���,�����!۞=
�=�p<�~��p�=ûu=M4;��1����<�� ���d����<�N-�7���dnx�t�`�:.<	�Ӽ(lt=l�n=���<jmz=z�<�ݸ��,<�ھ<�F���F���H�<��=�[h=��;�1,�">����<?R�<) =K������<ej�=�N��[W=ݞ��Ç<�Vq=Z.�<��[�W�U���<�D�<zȸ<r4 =��?��xX;Zt<U2�<��<����<��;��2�>�ՁC=�x��/����:p�,=gD������@n�� ��>A<j*=y=���<��L<�SA�w��-X�j�=�B*=�ma�=��P=�|���U	=�콻5��<���8Q���(1��VH=��;G��!�<j-&<��,=�-=x�L=I�9npm���9����<��<��A��'��c������
�=X,2=�P<3� ���;�"��m��<'�Ҽ"�?�ѳ4������<,#�<��2�\=[�_< �#=w�}N�BD=�1�:��h���e<��+=N~9���;�22��6��iKϼ��S='fc;���<D;=�a1<sżA�]=��6�Y�'=蹃�1��<�����w�#@=�H����i<cHb��%J��A@=���<��/�^�*��&��ЬE=�DA��G�<S�;�:�4= �<^�ǆ�<��Y���弭D2=�B�<�󁽆#�Ԗ��*���"c�<��e�2��;�fI�V����"<de��p$��=�_;m$M��C���=;=��
�Q�4=\t:�ؕĻ�r�R�z����u�?m =XD�|�=���m�἞8V=f�<t=�iM=1�%�i<�<C�;���\<��f��<��~�<��Q=k8���)��ރ<iG�;��;��ݻ �x=�}"=ò4=�`7<Z�:=d�r=^�B=�tA�"�.�C��<R� �a.�۸g=���c�R=R���Y�;���׳���޼&��<(���sBp�Ȋ���W;<��=oB#��j<�Mk=T6K<�=d�T��d/��v =�,�c��<�U;��6�Y��RT-�z��;]�7=�f��
T�?\��g}�iTe��ݼ��2����Bk@�aw�< }��	�:�#������h�(=�El=�j���TG�����C�D�G�Ő0<��h��Nf�p��<c	@�s��<:nv�^?�; Y5=�1U=�PG��*W���ܼ��H�=��A=��e=6^X��O׼jE=cc�<�+�<u@=.��-D�l�弣�%=�R���<&�b=�I���$���<��<�[��!�����Q�С�<j�^���L�y�^�U��hZ*;��滏��<��5x�+^�RR�<�~=ܻ�:��<�z<��A=�u⼮qH=Ǹa=�7=# |<H��<_͏=j��=�<�S�/r�D��;b�?=����4fI�ir=H��;����n=2�R=��[<�]�`�=-�<K����Y=n*�<W�G=�^�=<4[9y�=�(t�n'��H0=p�'=e_=ob=�>a��=>�<Vݙ�ư
<�K'�n!��Å<��=}�y=�Y)=a$ ��w=�����+=����=>|7�NU6�ـ*=�t���V���b=yi�<-2=8̛�F�H=�k�; ������vx<����<i�L=!O���=��R�+O=���V�E���|;N����};�7)���\���Ϻm!(<�A0<^��"�����;=A�=*+�=j����7�<�d=�+	�����)="5N<��D=T0J=
B= ��4=xe=+�/<��[�۾J���=��ٻ?�<;7�u��qK��������q�<�r����߽���`=#�9jV_=�����j�h=�p�U���o���O=D�ۉ}�����D%�;>;fÊ�L����xF=�==3��?��<Ia==��g��<�� ;�����':K==R�;�����<�O=�uK��Q���2=��>�=�L<1^���*:ӫ6;�� ���@�*�Y<��=267=�XE=��<*2����n�>=�ҩy����<�?<]F�����<<�x(��4��<�ھ;���:㍩���H����<³��'i=PyV<'s:��1���G<8��4s;��a�E�弙<4����ɻ��^w��'{=y��<������#;�.������[2=_�<��<ě�<��>�<��<�ef=
C�ᖼp����L����@��;�ȼk�=?7�<
W=a� =�=���<��(<��<zUV�Iy�< ��<Z���t��߻�Cf�%Fw=^$="}��}���)
��1���N�Y ��5=���<I3�&�'=�2%�#_���$=>8������\=�4�������L�u4=µ�:q:I=�4<iX���-��I�<e4u=&.�<��{;��Q�Er�H*�:��кODA��9��
�����5�[\���xۭ<,a>=�	=8␼�(�RvA�w����`d=Gǽ<-d�<�G<m7G=i�0��=�a7=��;v~L���`�<�� �ˎ�����&"1='1��S����Ʈ�<���<h�C��ڶ<
#S=>�ڼԭ<7<G���C�<I��#ʊ<A�<�7��r9<2��<*=I6Y=b#�H�=�Dp���B��p�;�ܺ���6��;�~M=�P���C=-8�n%����<M/0�� �~�$��u�<�rW�e�,^7:l/=�]=P}d=�yV��O[=6�l���������9�=v;ü�j��F=���U�=��K<�ռڰq=]Ѳ;�����'��.���=.G��4�I=�)=T��˿<3q�p��;<�ٻ��T<��<yʈ�wͧ�ƒ2�ҏ=�/H�f��;Q�A<�3�<Ny�=��U�Ի|Z�<�sd�]��<Bː;��=2=V<K�$=��'������=m�����`��0eX�a��8�<�N澼�Ox<ú�<L�d�$��ɚ�<D�4��5����޼ү�/	;�u|����։d=p�a<8hӼ	J3��P�9�7�v�'��z#=a�<��U��G+=u�z��<);Otp�r�2�"#`���X���/=��a=0|	=��������P��s$B=0����3<j !<�l�;i����.�<��D�_n<<��L�}H�'H����=\(8< �I=~����xK=S=��-=I�~�l&�<�e���=;�c��MY���=�"=Gܔ<>P�<���<��=6�E=QKq<�hw�Tq�<6�j<��1<"5C���N=�3s=e<:������;��g=�%���;����c�!�/E���2�f'��D2r�u7=é���<��=J.�����<��Ǽ>x>����9
��=�N=jf�<������4�����5�Q0��fX�@��<��5=YI_�$�9=��D=��'��0�e�c�{���H�!�+��d�;M�<4�`;>+=�V�<Hn�j�A���<�|�_��<�*�a��W�mo�='P&=y5�}�<w汼W	�ȉ�e��<���빼d��<y=�E�<H�;��ݼ�g��׼x�=%���dX�*vü/2U<��0=� �t��:�[<2�/�<..��P�n �=[�=AB =^:��H��J=S�(=��<��<z�=��j=��j=BB�<i��M��<�~<��$�+��<vs,�Sm%=	&;�"���U=�G<3�9�z�D�_�'���<���1*;��=e$x�QoW="=��<s^e��v=H�F�2n�� =�J<u�S<�C=��$<CX�<@j_;�ј;;#̼5�J��Ǔ=����ǻ��+��#�sS���\=�
<=lX.�l���S.�<�n=a2<�yh<��;��b���aa�<��f�p�<<��8�;��̼��<bL�;D�2��s�=�#�<�9F�X'���Q=G|�c~q�-=�ɼ�6�<(��<����o�;�z`='�b���>=:�l���1=�T=o�i=G�c����)�CL���<g=zD缙,y<�3X�31���.<�N�<�� =��<z�=��A=,oN<�<gs>��4v����l=��<e =h�l�*�����=e<S=qk���Ր<^n=�'=�xW���<49�mTI=5����(=�1�����~0=���<RI�<s#P��)=��=֨
��k=�5���T<��r=�`��I�C�s��^��<��-=�����%=�=�Q��<)�{�=;=�~�w�z<��;��1��$N<�3��dC=OZ��wɼ��B=7�8���<�&���=�=������I�I�����<Z@=|���%����i�^=�󳼬e�<��C��-�'_���k=��约�x�Q��n$�y�=�j=��c���4=}�<�k0;_֌<$~6=��;rLQ��~=.j¼1b�S�=$���N��/V==�+�v>��-�_��"1=u˼��,=|R =�'�<�;o<�����`&<�Kk��Rh<�;f-_�$>��_EM��q;�0��<0mU�U=^�Q=$ם<�0��f�<�M=��I�9�&�f�����Ҽ#~=0���0�<vn4��&�<�(��&;<��<8�K=幕<��;=�G�]� =��o��C�<���<uܭ�u}�uSo=�p5�4J=�{�;z#=�R�0�D=�f�Txn�w�Q�LA|��=��=�f�PYo<X�=��<��<�J@=s����+��k=�;�w=r���q�	�JH=��^� �����<�'==��ϼ"	�+#L�W�#����s?@='�o=Z�=�y���<�������g���x=t"��.��;�K=��_;�<�I����<�<僵��Ci=t��<�RV<�;S=8�ۼ�35�7˛��������:��<�$���<[C(<<�1=�M@����d�&�
!q;16;t,O<frS<!��5�<���w�[�<M28=
�N��T�<�ڬ�i�
��`�����:Ş:�cT�}����{�������N=G$_����;��ܼ��!�����`��|��<0 {<�ti=`K�<M��<��<*f3=�1Q=o�9���<�@=�.���	�<�F�<͌�<�K�;"��<BЅ�g=��<O�+<o#���P�;N�+���n�<!��<TΊ��F�m��<XR�����E�x�\��b=sy<��0�e��;��={fp<m�r<�%<��\���:��)�Κy<�A���=[E�I�T�`]=}V3��GN=��;q%�=0,�<�zP={)���!���r= �V����<�����논w-Y=���;k�-����;؀g�iը<�}�<�&��gj<���;�-�T.�u9��Njm�?9���c6=����;���0��0?�ˍ=>��<N!m<Ί<�悼 `��~0�'�Ｉ�T=�� =7ݕ<L'=(�i���<��᪄�d����/��Q�} :=��<i'i<�D=��r<V��F�e��HE�)м�SX=PU=MC��c=��_��'-=,����B4=-F=((�`���Y/�<��<3��<����|�H��T��<��ϼ$���\�<�ؼ=z7=%�=���<��S�k�/�M���}E��*�p;��<��=�Ll=P�=� 1=)@�>��<��6=]j� h5=��9��k=U:ӵ<���;��~'ϼ��<��<�9y=�=^�"���)��h�<���h	="Ȩ�]m�<��<Ԍ��|�!�s���G���];>��?߼j�=�>���[=J�<���D�^:����y�<��<�n���I$�P�X=6bI=�҆=�A=�p������h��=�g=��9�+؎��69������ p<�JL;�K��,��<��8<{&�şd;�Q=�|�/TT=6r�<*�
�9�:7�+=h�2=k�-��.=l)=ib��R=�Rz:����6�kG(=�	�<Ty�/l�<�=.=�~�<��XbS=͜�ϕ���]�rVD=�y<p9�i��,q�]��Ř<�bڼXm=2�:��ռ��ջ�3o����|8=��m����&�<�㖼˵�;�=���<��K=��"=�E����J�c-m���[�V:�;�߇��0X�B�W]����o�7<b��	�\�'i�<<�0���<�D6��<�<s�:B���u�<b��1M=ah�;�<���<�G<
;=���<�J=OQ���8�t�f��K�[�o�Ht��tO<&ʮ����e[�<��μr�f���p��$`=f+N�$�-<R��<N4�g<��%�ס�<���<RNȼ: ?=�6��e==���<�8�<(hD��=��ۼu�f<�L�M�8=9c��`g<���� ����*0x��6=��O=����
��z8b���T��z<#�/=��\��Sx�/r�<���j���+=����� =��C�'~+�p�9���<<�8=�x&=2S�������=kb:���L���;�Y���R�6lż7bA��6��W'=����w+:��Ϻ��μ�g�<����/5��x�;���<ՠ�;��H����]=���r=::?�$�ʼ�G�<Z,8��O��#5�Zi=��V=�Gļ��4=��̼�|�;�<�<F9p��
0=s5Y<����\�Гf<h�|=���<C�<]*���	U=���<~�v=��<�t=!	̼�\X�'�<]a<<��<Ӥ]�^B�<ÍQ�iL?��A=մ���Dm�����4����Z=���<ؿ��'��<_l�<����<�A����.��a�=�3b:���=�a0�p�N=�:<�u�<�p�;)tp=ά�<WP]<2�b<�7=�]N�n����N��"�6%�<���su<���=��=�8=~B=q��<�7q=�5"=mh�MV(�~��B�I�X��:��c��z`=UlZ��<U�I�NB��ļ�p�<>Q<�T=���N;żd�=C0�i=����+<� <ښ��{}�<B a<����k�=pg�<��=�����C#=0�9f�2��绸''��"�<�깼�'�;��=�=V=qխ�WNA=��Ƽ�s����=w��<�!�P{�;��<P�;�d��Ի�U��Oɼ.[��m�;���<{&�;I�\<wPƼS[g��<�������o=u����6=�uo�Ϗ=Qi=���>
�'�_=���;�ٓ<1@*=n���]����v�<g�YK=i�)�;ބ��bS�E�P<�R��%iW�!�i�&޼��;��=rN!�����A9="M3�ZK<���b��;H.��S����
�#>��in&=M��(:$*=�ו��Z�;�xۼ�{�<�Y~<n�����.��;fk�<���bw����;=K�J��Lֺ2,N��ۧ<i���N���+=��9��C�;K�Ƽ�k=*��<� �;JrA�,�J������T��<<�E�2T�;��Y=l-�^i|�9�
C�0᩼���4�=�]f<��=�]<��4;��Z<[v�<�~<i��� L ��LT�Kl��=���<���P+1��6�<�E�;EҢ�Y&����Ø=xϝ���H<��O�";��X;t;���<\Ș�h�ѻ\��<["� `L=1����:�����ˇ	��V&��<�;G�<�����4=�/M:ﲊ�2܈<��X=�R\�<�����=D�O�Õ;���k�\=��n���<��=�<8� <0�3�l�-��
/���<�,�=>F<<9�x;��c�Z=��^;(d�<	>�<�;�C=��z<Cq��,<�pQ=u��<ċ8�Cd�=��Ļ�����:��+=tk����,=��������<U ��?<c�<<�>=q#\<��	��O.�SN=�F1��f���p�w�=��F=�q=#4h=�Y8<�6R=!o�<��=�=��n=�M=�_Q�
�iܼ���E�{=�%�<�b%�R�7=�<Yc=�s����<���<�e�<0��H��<��[��_S��>���}n=��K<k2X<�Kһnl�<5��<o���O* ���ϼv�˼�9`�i.=���a-���,<9��<�zN��3ۼ�&��}T=�V��g$�lú<4i>��w�<��Ct�_�5���Z�t�.ȳ�{.1��=]���q;p�?������H<�JQ<��g=+=A-T=��<EbN=�b�&�0=9��<�%=y^=��x��~�3�ڼAO��s+=�^</��<�ʂ���=
�5=� ��m=�X��FhŻ�	�;+�ļٖ�<��;@�@<�D��.	=�4�<_���'<L�<iX����*�B;"�޼��]�&�2=t3h���<T8�_<,<?�<]�}��SF<o'���=�&<�"���e�;�~=�bn=�D�-����8<�7�ug%<l�"��C�d)�v:0�E ��%��\=�A9=:-��P�.<G�?��<���6=�	V=�Lj=[�M��=�1{���x�<CO��?ǻ�v��}�	�(=�l=���<��=�(=a�B=^F��ܼs=�)n��1���A��My��~ � '׼t=�m`����i]��J�8�����J�K�y=�o���	�E뚻���<q `=Z-= H8=�E7=S����]�hj��y��Α�٨�-�.��.��$��-[��}P=NZ =�]�s;
=��-=n�n=ȲN=2U=*����k=�8Ƽ=Al<e2=����jv��?�=���I=央:�x��=4ļƭC=<�B��2<<$_V�i�:�,̼O���� ü,��� =�_��"i�we����T=tI���&=uN����.��H�<��+<ehd��1P�j1~=0�U=&?Y;G�2�2K�nD=u�%�%!
=�SH=�v�Z��<С{<;�v<����>v���'%=A�:=T�Y;[��<�+=�,P�N�!<܊2�N�V�l-n�~�7<�C�^h3�����{�f�=�0F=���<%+;2.�<SlI=7�m���p��t=����=j�λ�`�<ED伺yڻ��<L��F��<d7����=h����!=r�<��$= �E;��d<,�T=���<�4�"=K�)���G=~3�<�����P;F�)���G�	&g=Ź=xB]� JC�wG=���&=)�F���=�W:=;�T.<���e��<H�<�艼O�1����1�C�;HW=.�E�RI�<!s<�.��O<⛀�dm��\��&��<���<Y.����b���%��=����1v�T�ż�f�:�<���<�L=��;�����$��j�8�r�r��ߵ��C�<�>^;��:�B=�일��<�=�B��N� <��<v�<&�ͻe�;�(��D���jq<7�9� �@�� <�m*�:X������<3�9��-���&=*'�=�V���J=�'=07=�
�<�ͼ�L�7`ƀ�բx<!3��̼�!���<pD<�"<$!9��Yۼk� ����R<��I���=���GML=L�_��-=�]�<���<p�������� �R'=*��-�>=�7�<�U���[=	�<��;P9^=�d�<o<�;��S��Z�<3ww�*v?�Y����=�פ�U��<'e�p�/=�L���<5mҼ�b��G~�(�O<�a��9,=�-��>�����@�8�:̀���lM<�qԼ[�Լ�:��&=N�˻������ ����;����+��0�<C�></Ʌ�(���<�w���o�n��<�";=�=�k�޵�<�_2��Rx��<�;��Z<�� ���=�~O<�zN=d <�9.�^X=�-�_ʺE��,<pt����U<�t=[�X=���:Q{Ǽ�=.���N����L�<�Ӽ!�<�U�<Q�6�)\�;�x�<tk=l38��%p��P�z�L�چS=�3<�1��i�1bJ���==��Y=�"=�����`���Y=T��<�i�;�y�<D�𼵑Ѽ�5��"{<�eu�-R�<�� =dZ��e'=�[������q=W9=���j���<��'<;@h��.E=�T¼+�{<��=X��;Be=_�8��.=�P�<�3<��@<v��^j<�8;���<R�1=cz=�=8�h��� 7������.�<)��<VXX���ʼ��1���\\V���=�
f�|[<Ѥ�<���;𼖈)�,Fn���]�z�=��;@<�<� M</Y(��u%=�<�<�Ll=�Tb;��<'�Ҽշ8=Z�u=li%�
�;���<��ܼM��;2C/<��n|<\��&6-=�=Β1=��<Gw��4�(���j=J��8�9o;𐄽O�׼��.���b=<�1�=�I�<Q�<x��\����̷�����<ϔ1<�V������g�0�9��u�<֏;�}��u�<A� �	m=��-=����rH����<?T!=��ѼHk�4�0=���<(،;�r��v;6�	]�r��y��<��=�
��_�N��]�<:��=�_=��@=�F'=���<��f<I'�<��t��	'=�� ��2�<v�f�$=�%K<�$�C�N=L����7=����tك<�+�<�C9�v�[��r����D=]󾻈��=k�K=�M3��/V<���h偽)f =�k<�&�� x�;�]�<��	=5ʉ=��~�=2(W<����O6=�r��+��V��0D�:B�鼓�˼��*���a;T ��7%�<˚�<�j��|S�<�	��	B�4X��\��Xν����6�[�̤*=�ʅ<�^Q��!�{bb�)��;N����H=�[<��<F�u���+=���:��#������ۼ���3a��՞�q=�v���g�]��Gg�7������ƨ<M�E=Du���ި�y�8=\yj���R=wzN���U=��;��<�0=,���-:�ɑ;��e��;��<��<�E����3�˻���o1=]�<�i�ǖ2=�Y���J	=K.�<lcϼ��W=��k�	��ȗ<�ü�����=�j�Z��<b'�vv��9C=�����j=���<(��<��:�4y����<uB=�Y;��s��<����lc/<R1�<��:l"��l�;~=8�i��W�<rc����=�Q�< �b=��&�_<�5�%���[�g�:w�X=�[F�:���8Լ�+:�>�~�} &=fY$;ᝧ<&(��9��^6���m=�OC=��<��=�=��;�Є<�%=l�~���g>���@4<�3���;=x��<rj=��p;œ=T}W=�j��(��J��S<��0���]�j)=P =�?K��9�꠽ր��d�\=��w=l�;͸�C��<MfK=�.:�f(�Dd�پ��Z�>=U|+=f�=� �<և���3m�(f<͟(��<���r9�=;H�s�n<#w�<���'=����<�i�<J�~<떛<��˼��<ms{=��(=#Q<�u�<�7�g%0=Fni=Ok���N= h�t;#��6;�Cu%=��K��;�!A�g�V�w�#�0�[�ւ �oh�k�s=�1R�Q�7=s���:W=�o\�#���;5��F�&=��k=h,<tq	<�Ww=������7�9�pJ��ǵ#=1Y���Δ���{�w@�<+ހ�q� =S���s��9����}=�I=:���&�<����Y���<�h��Z5ἒ$�ϴ6=�d�=Q�I=����f#D=�W<,=^�ʓ���!K=H�y�uMż�[�<P)=�)����;Z�=m&f�f:�+��w% ��V��r�1�ף�=&W�>���e�T<)�~;���<eԔ<��b= =���;��=��3*����<����F�U�r=�o=SD�qI(=F���1h��U=`���@=e�����<�_[<��<(=<=�����֥;�n=5��Z�;�=��;�ֻ�4;��ټK�}��X?=�3��A&�<qm�9a6�������C����dS=�}��Y�<���ē/��F1��	e=�=Y����<�	[���ɺ��r<diB��_��V�
.�?����|=�Ё<)���宼*:V=ƞ��X=ɑ_�Zp���6=�v�-�N�� ����]=c7$�3�C�#�2�ۼ�e<(�c=��X=_�F��
�;��o�k =��)=�H%�
�=<Y����9g=
�L=�9�<&�t��?'�
�;��<��=��6=��8=s�=,:�!I�;q���rؼi��=�f�kd���Ѽ%a=D;�4�_P�<�5/=k�4���Ǽ�;���i�=��%�1J�G���!p=O�$����:�ݻ��8��\=b��:�H=��E�{�<wd3=4���f��<�m<����yܼ��C<����[/=�5�e#���ٻB8���}�J^�<�ܭ<z�=P�.=��J=���:Ǖw<��H=�ݼP@��
�<��g�7)3�r��<���;��Z=DrM=�޼��B�����';I��i��<���aL?�5�=�`A<��'<�|V=�0������=?b,��+���*=��=<Ȗ;�ɍ��0��K ������3�<�*��}�����C=��9���{ =�ZQ=�,�� ���-�����[�=\�=N�6=b��<�����o�;�r�<��|=/*U�7H�:7
@� W��y?=�6p��.=1�˻��`=-u[�SJ��厽QB<�!@=dCٻZJD;��+=���<}�?��5��oP�61R<� \�*O@=Ue5��M��4p��p��$K�̑�=�r�<���7S������BT��u��I5�@V2=O�B;	�=#�<�<��/�z1E���4���<D�7�$:�h=lN|���A����#\<�X�<_��0�W=X�лyb�<�ɿ<a	y=�����`Y;�:#=P����=����(���}X<�JO�s=>�)��������<�'�:fɼ�R�;G,+=ow=�M�<2�2<�O>��w�<(�4�~��<GJ̻�9�<A=N���ay�Q[0�U=��6=
�=F����B|�u|F=K�=D��<IbJ<8,�;�&����<g�=��<=gw���¼�Ř<.�&=u�s�M=qbO����<u�'�����<�<t��$g��=Q/�=�P=?yu=�<
=�C=��Ƽ������O����<�J�<b��S�g�`C/< ��b��a=f��^�;Kz⼊��0��<ȫۼ��6�)���3]^��D`<�`��� �<+�2=��='�H�x3�DIb����<R�c;�.s=���jX�;1��=nM�=��_;�dP�,�;<��u�ڬ���<C	&�0B�;����	A=X"i���=�
м��W��*:4�<��X��{%=a��<9U�;,��J2��W<]L��P6=�6༖_�
W�<�U=[?=�c<g5h<��\��V=���<��=PK<�vo���:ʩ(<�D���!�8��9^��=�V<o鉼�<�3&=��� �<<�T=d]��ټ=��<����༏Ú:�bt���`<e=���]�R����=ܹ
����<N�����\�j�����<��μP6������6��S �Z=��-=��(��%F��+��OB<4y�<�-=�!ٺ�G��/�,g:���<��V�w�;�N�;R�ɼu�F<5Y��ʉ�<R����\�mD��;R��<�`=�(=�6}���=��=�L=�.��=&/;��6M=?�o<�h< �$�<�8�<X*�<*�B<|<P;��=�K���\���Y��E�<?�E���d=��e=�36=�m�;��)�K�$��_=����<� ּu<�lf;�rr<������=�X�;��{<U\l=%k=�1A<qz<+�m���W�,=0YO<xx�<�|��<[Լ�i����<Z<���P��FF�*庡��<R�[<�K�<8Z:=#��9i������`)�Du�����`
���;ng=�屼B�.<��<\�
=	�,��N4�dJK=#�X<Z<A��:�f��Ed�����WZ=���;�f�=T��V�3�UL��F������i�;�ְ<��I��"��|�-���>�6y��\�,u��ǯ5�"��;E�,=����M.=�s�<��m�N3�`����T�,!=,�=�<&���<�>��r�D��S�^lp=��#�4�V=��2=�8=�s<q��������<�n!��g=�^^=�����h=���<��N��+=i��;O�¼�xl�=v3����=�=��CsU<f�T�g�==�aZ=c '<`��<<��< �;[�_�Ï�;@�<H�ۼg[�<��P���`�!
I=�^&=��;F%�G�`��`P=ە��K�<uL��B�kۺ��ּj��U�;q��<o�<�
ﺬKh��ǹ��<� :=�6o�W 7��Q�ĭȼ�Я<]�3�j�7=
����cD���;�&g���<�Rk��ie=�z<vmS=��6=l#�<ǸW��"e=Q��[�*=�ƙ<a�@=���<(�G�DG8=����FǼx1�K7<�4�<&�;�=�ō��(�I�*=�
�;g*+=�@�<0B�J�<��!9�޵;��=������?=T���wV�=�N�<�|T�z0�� =%����ڼ/D1��Y��Ն<#.���<���<R�<$�;�wU����$��+�<W���J��<E�*<\�ּ	�"<=t鼯�����J���-�5
==���������!O=$�����<�'�;O1�e�P=�{1=�c*������>=L��<��ռM(S=ʂ�<8�Y�|�=��o=�Q�<�o�<j��<�
�.~�l~���
���
��={���4-���ӻ,��ǋ=Uî���c<gF��1$=[	R<
���c!= ��C=0�6�b<:�=���<c,�;����u"�<�mI���H�)�=m��Ob�l��<lp=�+@=�>o<��=�2A={Җ�+/�����I�Y<=�F�vx5=/���"1<H蠼�=���űμ��=5��=��H�� =��꼑]��2<_[d������*�u<���<�	��&�g��]���%K=��=�I<^l����j���ٻf#����<뷳;G�.���=����}� =(��;��N=�&Ӻ��ټO�C��f5<�V���5U������6����<te�<Q=����x��<��=����%%�_�W=+4<�QT�1�����a�=c�q=�Hͼ��[=j��zLʻ����ǌ/=���=�<��3�;GL\=��=��F<���<��-����<��ü�=�BL=��<ʧ4=kG?�uֺ�J@�7�=ڜ��aּ���"��<n�}=_T����<�qZ<�߀;�F3<ڼN�����==���<F��<]��z����"=�pW���=S�+��F�z�2= ��~����-�q�I��>�Ӱ ���'�u�,���B�e턽:�ͼ(��<�K&�3���\f�6.=BP;=��<�tE=�����l96<�؁�X��<��D=]�<eH���=�5���=��2?<��u���w<;�==���*=�����<�`K��]�;���S^Q��˱��n=�4e=��J<����H�v;�-=�b�<OKu=��
=F4U�� �=���
`���=jH���H�!���N��<�ԭ�Jc:^��<φ&������N���I�o�1<�)^=��g�q=}�7=����k�Mkq�
�Gͼ|yS;� �����|������T���7�����0=�2J<]��<�	=~M�<G?�<�?��'l�u�k<Ci<;��;L�	<�v���]=� ��P�9���<�-��(�r�=�r�^�=v= �I��^U���)=Lۼ��X�轭<,���-=PWC� J<�/�<`��<�+:�4�S�$%�<�x��l�2����<�쯼ս����X=ƿK����s>=��=�$;
��<w4=nl=���<�o���<�k��%��F�<m=K:Q=l��<p߰�oi�N�S�(#X�I���l���c����;[�><�X; S���sa<F����8���"=!�I�s�q���\=�.=�h�p�e=��	�L����<j�)<��j=b}=���3�<�q�9���L��v6���4=
�<H`=BF�<q:��,�<)R��,�|�	<5�K�9�L:�[u<��2=A�I�VS:=�WE<*�S�����,=��T=m&=Hj�I��<I%U=�.�I�.=�4<R�
��=��S���!�ɲ!�n[='�+;S�=R3n=I|.����<��ڼؽT=Y�M=u�n�R�,==z����H��U��L|���H�f�
��p=ɲ��k��?��;�<�0�D�߼�o|=H޼�u���|�y�J�^�6��Ղ�t����<���!�Z�RbV��硺S\M�A<5,E=��b�P{B=<��7q�|<��0;Å�= �z;0,�<�ុ�mX��¼�.=u�^=>T�pJ)��~���4�o�G<5��<%U=���<�y��-=|h�<�7��J��<��F=��_=�a;�~ܮ<̢h=t�0���#=_��;�j�U{!=?4��њ���;�s={�;{=W=�\ɼ�5Ƽ�M���}����{<14�;�-�EGۻ2�<W�	�l�����&�X����*�$}�<�gs�fy�;�%L��cr��M*=����Mz=c��!K=&n=,�c�~>5<�?��~�����a��8ʼ�V<4!�j
�<*Nf��$꼳����<�1ջڀ�9.���2i=p��<�T2<Kl�Z�]��R5<VY�dL���M8=�Z$=ٵC���+=�����/�;���=pK�.��<ԟ�	�#�{�qƛ�T!z=��9<3��;0?{= �J�CS=�Y^�W�:�Bf=]�S�dl=*H�;�ef�y*�j�I3�<�Gr=V�<;�C�I�<�@�O6�:���B���_^#=:2��N=���;j����M�<~��NN�*,=�e�:'�X=uQH��!<�!O=�!<��<�
a�*���pU���49<'�r;-��<�����FP^=�4���޸�7��򷟼"Rڻ� ���N�<��s�ļ2T��=?�<%]M:�� =�H�
��λ��0�i���m^	<wM��ұ�<_�T=K��Ѵ(��e��Y�M6����c=hτ=$z<2��<R�X����m��<�x0��/<�a�;"�x����<�lѼ�,�l�J�48��oLA�V���J<t��P��<�)�=,	�0=L�c=�א;�:M]�<�#'�� �Ɇ�<�<�I=ebn=Si=׮�;w*=2 =cI4=��U�]g=�M�:[�2=Uĉ��ͪ;I�]=�.��"x<~�x��<6�B��;��4=�;=�ɀ���=��ؼ� =� h=8<�,�<MO���>=gե<����I�;s�M��7�;}�V�e7�<�L:0�U=��k�@i�<��:�rF�S=��;Ρ�<�Ҹ�^F�<_�.;M9�����n�X��Dw��%$=�#=Η�G�E=٧Z<�'0�k�<��I��}B=��y�lM�o���9=&��;����[⺼ !5�Y��<������`�
m=h�	��P=-Rn=�"=":��9H�4+5�L3=t^|=�=�Q;+���F_]<C���e����E�J�m=o��t��
=O��<r���x������9��O=9��?Ds�#1=
%=�i�<�["=�7�:`/=�-D��;�J���/]�?�	��Ԃ=�O=��
=4�[=�r�R�L�˽=�ؼ�7����^/G;��=����� =��$=d�,� =˕=�QE�$L�i{d���|<�S�1P2���v����<��<�F�<3�<�����c(;<�@��xݧ������e�.1����>=e@(�@�)�i���K<z%=�Â:�E=�R���H���0G=�D<�8C=��F����;4��<H�C�cV=��<}tQ�e`��/-��
�;һ'=V�7�s��k1���<X/R=X�`��}/=p�/=U ;���M���=�6i=ׂ����{<8�<[xO���Ƽ�DY�ɓ�<����ƯW�D�7<��[�}@9��c$�ZԼ�����b�#=z#�d��0%���=�|L=����N�;�4�u����r==#y<� �;j�Z��;�;�'`��y.<e�(�J��$�d�h�%f��W�u�R<��;��(Kb��kE=�>d�:<�;��<[xJ=��7�P=ե;�%_=��&=񮓼}�(=�Q��L<���<���<3I=|d<�9��6=�S>=GRV<��>q��^<sL=��p�]���M�<��~<r`=�`P����<�x�O+=uTQ=�s�w�A=V*2=`�ռ
O|=��N=�*����<���<{aA�FR�y������<+m�<��r=!�<lB=�3=~�:�xv=��;�6��o=�n���4=���<( �<+U�[�V=�@�8�"<�M���������<���<��=��<0{Y<n�=,��<_j�A��6P�~�(;�+��a�%:w�?=��Z�#�=�0^=wJ	=�T��raL�Pkw�!ܓ��C���<�S8=�9=)�_<�K<�<S<l�
<�\=�x�<�����l=�%��tJ=��D�W��<><�>=��F=)>[���r�¼a@;'��P;��V���F��A=i�����B= +7;�ⷼ�/�ATS;�D�R���������k��I�K�;�C�;No!�x$��?�G=�OZ����;��<�31<�˗<��ܻ�N=,-=�4u=��@���<���m��*輳���㫼��E;���;ɸ<vyP=e�M�îL='�7<��h�Ih'=ޱm<Y��<��|<�8p=�ڜ���<����p����<P�7��i�<��;�g=[���>=)+��m�w=ڮ�;!�r�Nz=��k��j$�j�3=b�y�fv0�΋]=3=��T�O<�s���K=[�B�� ��+=�jӻJ>��dP=mAҺ��:T�=ޛ�9q�+=�o<sgl=��9$�Ηp��<{Ǹ�Q�<��L���Ǽ���(���[<=�3g=�Fq��g�<c팽S�2<�μ<RLS���$a�;+~� 1��cN��|�4
�<��`�%�O����<�-��Z�;��}=��<Z9;=��;w=贉<5`����<����kH�f�߼��`=��c���/�@��G�����_I��ҕ:=v�<��K���ּ�ѻ�Ŀ4�B�;�r<��<�K=�;�ф=�ܦ�jĻ u�5�yL�<�z��U������#f=��<Մ缁z(=��<o�=:X�:tX=�������E<1`C=d�����<@a=���<�����):�f����S��m=>l���x���<�5��<��7�A����K=J=���<ăT=�d�:ܷ=������ût^�<]/
;*��<@�-��\?�����
��<��^�WG=�:"��<$K���<��=ds<YR�?�׼˒�)$�<��w:�eW�q��<}Ô:|��8�"=��r=w��Q�W=�\s=��;�|�{3�4����;��Y�~��<���<��_=p3A=P��<X�6= il�U:K��%�=�Mk�8�'="�<\�A�{4<`9�<
�@���	�H�"��|������<�
��x<=oq��;=u�"���Լ��O�"<C������x�<�y5���:s��<��<��=�*R=���<.\u<ڹ�<S	<�fܼ�"q���;7뺺���m"U�Ǖ>=e3�;�O<�|�</�=�ؠ����;����s��7:"�=b/��H�x༹���gG���"��j�;�N����4��<����aA=���<>z<�U=j7��}��D=֗=OI#;sn7=T7�C J=5�;~�~<�ź<�hc=��\��1���; ����K*�B<@ij����=�S;��\�g	�md=<7I=Tɼ^1�=���<�=�=�۲�˲3�_=&��;bh��r��;�?���@�(�/���Z�>?F=�&=�Mɼ��z���e��w߼��2=&=6�=���t^�p�"=��O��>ͼ��<5�<sX��=%Y=�Y����Æ��u��=�},�� ���$�\cf�|,���h���;EB=[F=ҧ���<)J��9�;�p�����<g=�<��;�֌<U���=@�v��M�iLۼ�
<ƪ�<���yg�]�}<��p�ۙ=E}-<] ���h=�@��	���t��� �$1=������a�:���<k�b=�ؼk듻�1%;W_z��z=�Kڼ��<�"�<6	�<-�=|)=n��;��:�n�=)��+�T�缶�W�9����i=��M��a=�|`��\�$�ں�=�<����O�e��[+�<��>���	=�ļMk��
켥k>=��=M�;EA�<�t�;�ŻI6��6�R85=��=�;��Bs��E�<c[_���m���S}�;�pM=���<̠<3�<�����'=NY*�PU������į<�U="�=�?<IPB�.e�:h��C:\����<�O�<k]G��o��;M<�[��%C=��k���"�\NQ����h_�q(Լ��;���Dz��z�3���<�*>=��,��T��<��]=�4Ӽ;N=����n�<��=7Vz�*V<i�1=�5!�\f�;&4<�6c�<�;��S��PN�6��:�-=��e�8��<2�D��P�<=.=�yK���ϻ�n=4ȼHe�����ۢ�;�8�<=�\=5�	�1�J��>�ܝ<��3��˿<|�r=��g�O:�@��=�G��z_��)�H�P�гs�r�(��p�|>�<��0)�b�(;A�M<�s�<���<F����<��<�;͢�<��H=/���y��� ��B�*���<�Z=꫁�d�G<$�����C=5x�<hs��˽<_,=#x$;ǒ�;w�<r�R=IB�
�1��V���̑���_��OY�<�H�<�x&=0�h;|\�<܆$=���7<;��<�JC<��a=����ڲܼ
Z�<Y���/,:ȼ��*=J/=$�弇й���%��	^�϶{�5t!=��;s�ӼN=�<p���h��ʒ�4!A�I���$�<%^μ�6��~`k=Ж��5�̜��LL��A�3@��(��WI�<���!9��%G+=>����ok���ᶼ���;p^�%a,=#t}<�h1����<��6=,U;pY�<��sÞ�=��<��L�d=K����np�<�b����p�=���=��g��e;<�I��=�.��;���;bμ�6�����zE�<R_M=Ix�WP�[	�?�=�.Ƽ{$Ｍ�<m�<=p����S=�y5��x�~��R�V=���l�ƼU��tY=ig����b=)��<��i��"=�--�P�[�}��<ں
<c
`;�b=������<%��?�=�L=��=v��9�ϼj�=�ܠ� ��[Ǽ���k�=b(=ζ����B;�|��#=��<�*�<y�j�p�=.��Һc=�����;=sR�<��<���<S��99Y���3�S�ػq�v�[`���=�6
�i�-<Z|�<�AL�Iv3���?<#hU=�/�<�6ȼ���<�������pc�<Y#�f(M<
�==�r�;b6�7L$<���K9��x6�|��d�4�4$=�>���*=[	�<���; a|=�T;�=F��<�D���ؤ<�Ѕ��Af;��="�@=�=�)$�Y�6=z�;�+=��;R��~�`=������:=$<���<�@B����GfP���<Z�=��8<JB�<��<C��^v<�K���.�������|�#=���JE�<vO�;ߐ�MM˻g�U����;�񝼜ʼ��[�M$<���<,"7�]˼Q�ܻ���<�z,�c�ڼ1=�J�<M(żX�<.7=�qO�K�_�k�<O,=���D�ƻ�l=�F@�<I�
=ѳ=��'���w�:���5y�+�==?�<�s
�(����'���l9l�0=	R)�=gN=��=I>Y<D�R���>=��+��<�,o�1�)=�6M��Cȼyσ=#Fa=�"y���a=v�k=��9��ŉ<)ڟ����J�C�"�<NJ��mh��J��<8�<��/�'�W�7�a�>=Α5=��R��ӆ�>Qq<��D=!iQ��u��<=&g<=��N=z}�<x3K��nw�%=T|�)�<�sl�֎�<��/;
m=�.���*;�Q=�`=��!=E ��&��=.=�^�h�ۼ]�=�����H�;u�P="���YN<I:=�BH=�m?��Ӗ�wj�<8�Z=��6� r-��
��7ݺ��a"=}U�;�㼸Yѻ�Ω<Q(� \���4����L=��}<vQw���
���&=���<��/��~	�����ߒ�F=��+=�D=X_�<����╼b�/=�y=�7��$"=��ʺiC�B#��c=e��-��<��)��!�<�"=��Y=�KO��xG=u�<��ۼp���x�Z�$��e��$�V=��W=�~�:yV=Wn$�9�#�w��<���Ap����;�_:���9<#��<� �;$��s�(<ɗ <W�|��E�;�>�;��K=�D��&#��yB�/�|<'Hv�$�Y�-(]=@@�x�=Uʕ<"�ǻ��=�|I�=�2=�j�;녦����<���@:��:=�[��ձ�<�H�H�	=y�n��w�=,��;���Z�ؘ=��*<�⼠L�:�gA��j<Ċ�<�Ym��1<L7=�f<;(���W=�<�E'�	ᆻ%���ֹF�e<��<9��<����|=�;��8��<Tm,�WlH��!=��G=	���o⼦��<�	Z<+�P���a���c��tU�sb;�%��6=ʰ=��;�KI��ż����>��A��<Әq=\	1<��P�i;9����e���=J��R�ȼ5�P�严��˼��-=�]��xoV��%2<;�к�9�<[���X�1���_�ϛ~�q�<v�1� e?=}4��I��x#��Z�;w�M=��h�ҏ�:ʐ���V���O=iF�<é���P�<x#��=0�����U��[�;�R==T�{:�^<��=��#=8&=�\��nC<�=o&=d���JNS�z�.��A=�9*�v�=rWD=v�o��}ܼ �T<kr�7[��n����U���T=db�%G߼o�9=�hu=��J�ޜ�q5ּ8��:���zY=G꘼ʥ�<>�A=h�<;�<C�S=��!�w�=��A=	�g3@=w�8=�4�=�$(=<9M=��=S���:e{����<�Z
;�A����<e�;��@��	���S=�a�<@4F<��W=��B=�dO�b�!=Mf��t��''�'�j=KX��j=��)�#$=ߢ���f=rt=��<Q����p�=
S��#�<o�E<��!�"�9�gκV+����<��p��\'�XJ���D����<\��<%�g��8=��T=�l&<v@�:�Fn��1�<�Ҽ�ަi��1B='��)=W`��=x9;q\�<9Ԅ�;���<�Ԛ��y�'s"=4{r=H�I=gL�&p���J����=�<����y7=�/�<�;��K�|m���L==��;�Kݼ6�9�L<=C=�;�T�M�����ʻ�I�ߠD����6�H�+U�<��M=�^4�Y�4<�U7<�&~=�s��p8<�u=�mP�n�S�l�=��5=�vʼw3���<�T�T�溍�e�� =�;_]<�r�"`�<����<I=����|�C��Y��ٺ�����;4 =S[<��n����;~�f��!�3��:�~O�ES��W��A=�<4��H=B�������]�<oq=�*�;�Ŗ<��R�}���G��<U�:=|<T��z�9������<�ң;�-;���<
���:�:Pb'=�J�<@��<������;9[�z��p+��4Ǽ��d���>#</�w��!<��:b񂼹^������Q;`F_�O� =��9�p�;qǉ��!U�/Xe<V����<s����X<�8=:�=w�;�2=S$��F��<�5=�F���w�< ��9�'�B�<&�q9P��ռ���<�O6�%7<�:\:='��;�6=��=��<�1;p�<	<_�b��<'��<́���E����<W����<^�h<�EF�����Ύ<�EB��_����<�#~�gM=���I/=���7�%=l�:����}V4<9� ��#�<�=�H<�<z�-=Y��<
ƺ_�
=f�4=�mO�@��<[�=/7�<�����(=�]*=�AA�B� ;�"�<�=�<���\��5�;��J�G�ۃT<��[=`-=��U���{<
ƅ�v�I��_=ʾ�<��t�=��|9�m�<@� �RS=�%E���=�-�5�T<���<i��;�뼠�<�1�<�!=��8=��
��͵�(|6�yB�><b(���w��8T�����LHy���/�Ec�<���;�O��HR=�$�<ځ%<��m���<�cz<�_�m�μ-�~;)��<��
���	���ܼ�P�<��<=D�.��+N=`bP<!.?="� ��$[���<�V<��:��=���<aWh=��=\Ҽ|5���"=��{�d�-���^;98�<V�<�#<�Q���<�,,��A7;��<b�=Sk�<�����9����<)�7�h&G���R�YA̼����?==X�f=o��;�|��#��to��AH=�;=у��p�<թ=��0�tQ!=K�Z=ƕ�<.EM=$����s=�C�<�y��<�59���<���: �9��y�<�Y�:ޜ�<�f5='#s�3A�<���<V'����=<34v���N�uI=xh`���<h�?=�3��6�<���<�z�^��m�~�;�(<N�<-���^T�:'�0E�"F]��pl=e�<��<�H��Q��Ղ$<��_�,�y<���<p�<��8	�/�U=vI��~?���a����<��<�(��x�:MC9=��<��M=�CN����GN%=��ֻÈ�=@}��;�<'1Ǽ`�ۼ����Q=�e=y!���l=��(=J�*��\
�%Q4���0~=Ђ=��4=@��,y;��^=�=��a=���!l��4�<#�KF&=��J���d��L�Tz<93��=��9��Z;��<���N=������26z<���<43='�8����n"<:iN=;��4�ػ���^g�<�p�<K�7�Vx��_r�<� c�|�p��Jf:l���ԟ��=�'��� ='=hF�<I<<��O=;�3��>=�O~<y� �K�]=/=�6P�*<�<�XX=�9Z=�bƻؒK�5�w���+=Y���+	=��?=��b�r"����+�����gB;�|=��<��b��W���`-<�a+=m���;_%��	G=��.�W6 ����:��<��e�ΰH�1��<��$�W��:;%+=��<nCP�`��<��.=��~;NXJ<���',������	���q�2=���J=Q!�<���d�5���:����d�=�];�K=�ü��L;��F��/|=���2��� �3<�@�<j(=pG���Q���7;5���4M;e��>��<ȁĻQ��6��;ŭ�����q}e��̋<3BJ���z=�?2=}��%y=��=�|�<�ϼ۪�փ� ���E��<��<^D�;��@��Ǽ~}�� �=�,���=َ=̤X��Q�<@��� =4��5�]<��G��2V��%��v��<�T��.$<u5Ѽ6�j��x=�����<��輪�<.�s<�/�s*����l��4r'<�(Z��F��"9=����A�<��+�/�\�����#6�鴺�:�`�={6=���=���;��<(���L!�]�<�%�e�ټ+�U�CQ�<_�=
�=��P�)�=����=ձʻ�e�<��g�S:�<A�*<Q-ܼ�0�^�E��j�<�/,�Dp��
G��&��$4;�3=���<���<��ɻ�!=�Q��*M�gҋ��D�< 2n�'\��w�Y�,=oP/�ӊ�<�b�5��U8�Ƃ�<)ݽ;?o� C�ͽ!=�Kȼ�=��!h�cot�I*.=�TP=��0��c_�����ޤ�Uk��*=��;s���w=��Y= �O��Y��w���X�<�h���K�<a¼��=mZt��f5=u1 <�if�8�_�?E=�b3=��S=]����/=괓�*=[.�;�{;�no�$=�vB<ch-=�ټ�T���?�<�SJ<�a�<�}%=�X�fiU��Ƽc�`����<���;�X���<,�=��K��yv:,��<8up=��=��
<�w	�Y�Г�W��
���!����<6��<���<�#=4��;Vu%<F��;=�T;B�
���<Rv���=!�<B:�Q��e+�b�1=w������9�<���<�4��#6�;\t����[=�MP�6P�C�*9�Z����h֤��g��
���	=GO<U*`<0+�:ý=G��u&=�m��~���b��=Xz�;���<�a)<��<uۀ<Ɍ"���
��<޼�o=j�W<:��<.=���p�%�rz�<��/<P��<X8=�v�<�*=B�A=i���_;
ކ�^�[=��9���==e2n�
=��=Q�v�H��A�@=��H���&���=���$��!p0�{��<��'��=W�����Q�[=��<��=����kX��<d�M=�)��ke<6���=hײ<|�Z=p7<(�ѻ� `��=�;cb�<Z��<�ʹ�=2�<;�/�0=�Y�[������,�=�,c��ڈ;C��ݴ3=�0�<Yֻ���v! =��6�aUv=X�<��H<M�/��#�Y}=�/(��h���%�e�&=~@���=i;��)�Z�9=P=LL=��	<��<F� =nԆ�Ns�P~�틙<�`J�Ǥ:���u��f�<	/=Z�=�Iǻ��F=���=lg��x1�u V<S����;@=KGϼh?�:+q6��<=V���|��>�;�&j��'[���<��K������p�<l��J>H�Z"�1��:0��;�,L�8�=�t��?k=��W�5W*=c"��=�|������l���f����`��isJ=��t=���<<���B���u�'�	�<��T=<㽻y���D�(��+/��W�<R�Լ
�S�$q3=���<���9g���<�N����etG��p��}�ʻ�A=j�P����;'0�*�<ǯP��F�A�G�����D=�缃�o:�����h���=��ڻ���M7T=L�Ȼ�=�<��b=�?=�>¼�G!�Z�p=����⯙;2[=����!����0�=Sݼ�$<�Ӽ�05;Y/C=H�.;��!���_����<-v�z�!�Uq�<��"��>I<]�����ҼL��;$r=�c��^��ҕ=ce�0����(<0 ��l`��=:���}#M���<VG��<{�<J�I��\��=_6�Rݼ�ԗ<�<&,<�N�<�i���<�����;��	�8�@�R�ռ���<��.���f=����Q�Pw��S
���;��t<�=��<�'f<��:�<��Q<df��Q�=@6��fm<K� ��q�+���hX<�b�;~���+�<�U<P,�<?=�.e=�8���n�<�O=�t�<��k���=H�������<`Xڹ��<��V<c�e�rg�0��<;�!=���� ��t#���';�����x�[��<�1�<]1I=~�*=T_=�!=��[��rM<��R=��=��0�0	P< D=R�~O=O�)��=����cV=�C�<��*=�&�<H~%���M�\>#<���v#�<�g��V=�A�ju��;X�z����;��9=C�D�1Qٻ������~�{�;ݱ;Y;5=��Z=��<T>��U���=����~X;\B=�Q\=�6̼���� �d��$x<��0=J�8=P�2=Sa	9�~&��Vv�GŅ����;��<J�w=��t;��@��[���	)=��:�#�"=��Ӽ�5 =�{�X��6�@�m>=��'�9<<W��<�/;�<<���<y��gX6=K4�<�c�[{�<��%=������#���.n^<��=�u�"
򼴁M<��<��1=_q�f�H<�k=Rd�<��}��~˼V:<[��9Rs�;��Ӽ8�����<'��<=�ż}�!��t=ן�b����GL�Oc=���vpA���)<��ּ���QuE=�<Q:=>���*�#�:��������;��=�:2��ص<��ܼB{C�a����=y��<�.o���=	:���vX=M�R���<�[5���j���4����<���U�;����Zr�<�e��9��Ga�<A�D�J��R�:��$=x��?�L*"=�0Լ�~�<�Y�=J'���N<�$�N�U��=��<���*��`{=d��;�o=N�=�r^; �H�*��<'P��k�"�O��9Q}<��~�|��;�>�5�<��T=4|=��<WL;=֟�;+�<�2=�ˊ<Q($=��G�"��=vƬ<;�d%��u<�j�;-ָ; {�;�=֏<
=]�.=���<��; Z;�1���8����<A�=[@;�*���3=�3�>΍;��w���< �&��	C�s �S���ά�����9��0�)Q=z����$=;����l�<K�<1/ټd�Z�x�9����K-=,���=�"	=<�==�+5=��7�1�t<�i =}4��`Z���<��n��y�#����;/���=m=D�;\R[�W��<��D�.J����_=b@�;u�==�P��)��j�F�&��<�r'=4[=�8��C�a�-ߠ<\>���<=�\+<'�h�e��#�(=Ċ��Q��<i�<��"=t�h��{/=��F<q!�<,
��R=�}���/=K*�<�F-=�^����`<��=���<�ݼ����N��i<;=�;��_=ơ�<�='��1E�7�����[=�I<�c�$��<�h¼��>��l�<���=$�������I��:����%�A�����*;�a5�P%�<��n=������D�<��0:J�R=��=�d�<�;�qc�m�<<�r=)�@�I��<�mл������;���:qv��2�<=d'�y���(<-�~�A��<�.�<ZG�w�<T=.
üY�<)�S=�9�<}�X�MZ������&=�B�;;����3�ט����D��U=��<s~��Ϻ/�����<�a�x��;_��:i%�<�r�<�<I��`Q(������=��l<'J��
�;պ=h����=�yQ=!�:�"���Q�<k+< � =_bļD퀼)pͼ��&<�<�9X=�0��B�B=@�h�_=�����=�~�=�tD=D�o=*�/<?:=��y;�O�[�Ƽ��%g=�:�4�x<{5<�i*=q4=��F�������<O����{q����� ���&[�V˼���z�����<�O�7�o�2�Q=SzO��l=��4<��L�> 4=�D����L�<��0�߼��~=�� =�>h:�O�<h�<M4��ƹ�jJ=��W=�l<��7��z�Έ�>Lk���?� `=�F�;$g[=6{<�<�<و=�V:�.�=Ju.�I�2=EC�<?=�,�;��S=m�3=E�Z��
�={���+��V<.�;�7�<,���8J<�w�<���?�=�W=���<��<�[���;��@=T�e=t���<��<�<%�=M��<l[:Q-H=~�#�
U=_"�<!ļ��
=a�aF��j�q=�����e��	w�KS��Jl�=��=?�P�in�<k0]<yo����Q�ּi�-=n	�<
�=x��<��� =�h<@Z˼ŖS�*.a�����QƉ<||=K� =��<��q<f#~��2�v���,j�'��<���N��<&�B=X*�<B�s�o@���Q<{��<��$��.
����<l�׼{3���=P��<%�M=�;'�o2�<��,8�2��֊��N�;������Z�۽<=�l"���<"Cq�KR�;h4+���F�:E=������9<���-=�4�o�;�q<�	��w�g���=�=U�<0z���"=W6����=������<���ac
=�)�	L\=1M;=X==d�Ƽ^e���_<ׅ���6�zp[���a����<#~ʼ�?�<�M�l� hN�3ϥ�UT5�����3_=~�#<��=���<�d��{��3Z����<��;�a	�-�j<Iz��zb=6�e<kx�9 ���T�׊�x,�;@O�zG��ڼ��3=��}=�>�<�"=d�'��=a��'=�K�<��O-����(=�B/=M=I<B� =�QԺ3�W=�B�<��1�z��`I��z2�����ܜ�r��eV,<5�U�J�=�w�]=��0��B=e����=pg�=��;���<�(�)� =�{o���f���=��<P=�g<�H�=��Y�����m&�Bj�$o���������O=�S�<�JN=�b��,�;�μK���Q0_��:���1�=#�3=�+�w�y<��Y�2��ת��i�<��:<|
=D��:��<oL�5������1�a��>���,:��YA���˼�;Gy�;/�i<��<2�(��<{�w�!�h �Cu4�.�Ѽq�;73=ғ,�D���Tp=a�~=hZ���db�H����*=.��<�1���WX=ힲ��ن�!<fw�<u�S��I=�X|B=��<a����缾�4=	9�@�=���<k��<�@=~C���<�o*=�*]��e�0����=��=�'���m=;�9�}d%<僪<�
=�=���{���%�oػA&T��7�<>�<���y�<i�����	e=p󼣵���<�7�<��W==�P�*	=P��;�NY=_P�DqL�h�i<P���^�D��{|��� =��w:�Q=�:�<}�������,=,�;��#��ƴ�<�[�_����Hμ�e=�1	=+��<xYu=n�)�7�<�2A=\�)=������3<�K=S6�.[4=����3��D�Ȼ�<~Fg���!���J<��7=�Գ�n%�< p�;׉[���K��Ne����(�GS1�_�<��;Y���%tX��ռ>���4�<�O�<3�<nU�<F�Q��<u�a����<�����77��z=\��;�=ew6�%�= ��<u�<�b�#/M=a<���J=��;�z�<�d=�&�3>��(��;��d=^s=ER1=;�<���<aË��o=V�<�@<IVĻ�o��^�<�=�\߻O+Q=Hf�<��{� �����;�71=02,=� �uԷ<��w=�y��f7����<V�H���M���k9�6=�t��� j=����T������,=��A���4=��b���f=�%f��+�ǒ$��y���<�
�<�@�<+=9-<�t��|6=��=L�_9�u<�==��=_z�<�n.=0_+���������sc<6e��,=�v=һ==VZ߼G�ٻ5�C����α4�6::*m��,��K�;�_�<vFi��м��:�B6=v�;�E�=�wT=��A�i�=82������ng<w�5���u�� ���F� ��<hl���=R��]���F4-=���OǇ�y[=S�=Q�;Ic,=-�<9����'��R�U01=�;T-I=��ºm&c�%�@�5?=�!���:m��1�;��i�kl�<1U���y������Լo܅=b�W��5
=�K�������<�ő1=�T��V��k�k4���:Q[��SJ=Dڼ��UټpV^�����p��=E1�<�a����Hށ��\���;:==Cr��T��+��"=�!�*��<�Z��$�\<xw0<�l=;�^�<{�����;T%��/=*3�<м;^{��NR�<~Ae�c��<�<�:�<H J�\�^<Pi�;2YؼB�=�2���;F 	<�.���zݻ�&e=#�==
�=o��<�|+=3?���8�D<��V=�"b=�
f�+#=�z�r��<��`���<�Q�< �����"=�<ٸC=�6b�DZI�U�8=�`
��d-<xq���r��XS=���^�����<'_=�k=z�=�~<p_��1+���8= ��'��<��=�c<i���c��°�ڹC�W��r{ۻ^a�oA0���:|�»P
5�P_�<�>c���o���B�[(�<��}�@�b=�Ǽa�r��>�;Ә>��=�t�:\-=@|X��Q=����0r�����U�Q=aW�;�E=�-�<��=f?�=/v��%=�E����<�xۻ�@p=��=)=N�x�s�����ݻ>I�<��P<2�Ѽ���#��K������Z���<a�����ӌ�<j[={+=�sj�Rޣ<J�μ� V�Ov�W�<�ſ<z�,=C@b=�@=_��!�<:'��s�<��=�⢼�o�;�MۻU-=(�޼'57��NE=xI�z�;<�+=�����|�@=Q�����=�V=�����8�9�m�6�=,��<.(3=��9� ta���=��u���+��=
c��J�<l���，*$����<��?��r$=^���7=Y���H?�<�=��﻾��P�j�׼X<�1;��<Q�"�
���j���M�h�ƻOl/�Z<s���e=�gQ�)�=��E��G=��J=����,=�$F<��K=O�:�x�����Q=ہ�UH=*/�x��@Y4��%6=p����%�R�,�s�>:���</�����<84�<ax�<-Xn=�C�<!�*<d<(���ڼ��̼S� �Ŝ	<ݵ{<k#;<N����<LH<U���^o"�(��<�$/��o8<�x�<���#'+�L��;��z;�4�<���<Ƕ���3=>�Q�InZ�X <ņ�"�!<ff�8�;�q�M�����A$=�9=:�<@x��uv=���;��<:�=�A=uO�;��>=��|;Լ�$=� ޼~�=�(��G��O�;��=�,i=�/=wq^;�4�:7�<	ٹ�c�=8�)����"̀<�֪;*�=ؿ_=o���=���<���<=N�=��<Z�<���$�ػ�3���<��=��l=H�w<���<���<~�	���r;�4=cӔ��/\=4h�<cb¼�0:���<����	�H�쀽��;�L^�V ��}��`i=A.��Hb�09,��W<4Xj=gHG��;!�a%n=�V= i���)=�ؼCS�r7C�3̚���U�d��<Q�"�5�ü�|i��+�-���?b�;��^<Y:�<{a.<XT=|W��f����;�$+���X=�A=>�
=�.��g,=]�I�}j=��H���=(����>t���׻�h+=�5��
=Oײ��;��o{��e׻T�=�Ox<�)�2 '�a�;��<!]=��,=�� =��;�Y��v��;8HS�3��<�����u�������݀=C�>�����4(!=D����
�T7�<J��&�M��M(��p<�����U�<�$5��]-��N=�������{~�<��,�%=0�޼���<��=�7=]��<}C�<r�K��G<���G�%�z=�	=�8<�nݺP��<�yU�nH޺�,9r�<��$=�d6=蜀���9��PH�a�C��F��5ы���E4��}-��G�<��o=��*<p Z=��ü�����>��hZ3=dV��6?=���;2_�sw�<@F��@��E��;�O=B������@k2;�s<m��<li�Y�A=إ�����%й`nۻH��#��<?� =P������<y�=�����<��\�FT��\��=��u���a=��8}d<֌���6�1Vż��@=J��۲@<�6�K�C�o�=Y˝<2�1=G�=��3�s���؊����<Y#=��E=������;fֱ��]��.�N� �L����c=�+6�����O���3�P	�<Y����%�����R�z�=~��Z?�<+ϼ���=���CK=��a=Cy�<^��������J����<X�<��<�Oͼ콅�҅=ȟ�X/���tͼx���p=|�׼2F����4��qt6�L錼�"{<�����=`�/=��f�@@#��}=d�v;�ߣ��+<���;�m�<�(G=)r=�Q�;7;�}�$=Q-�<C7=�M<�����qz�1���l���$�<D�=9�D����;�_���=�?�<nm�<��h=@}L�%�=�i��<��<&2���5�����l�:�>��w�R=��A=���<%�N��;�Ƽ�;6�=��s=ɲ3=/��;�@�<�;��}����:�cE��d��y`]<��f���m�=���<���<�>��6= G?�6�B=_[.�Pe�E�;���;�!<���:ڿ�<�|�;#K�������<?�?����<���`��������N=� �<�?�<6�9�tD=�����/L��{��D<@6$=$/�<�5= ��[["�p7<��g><������g��t� �	���;=u6=��*=�&=;[�<�{�<p����:=�}Q<o�=�@��Mc����<j�3=l=���H�A�<|=O��<���"=���;��<����¼�G�<�����+���heF=酝<�Z8=Ө#�h���Ic�X�L=a6O<^f�<���X6��R�i=� �M4��%�<*�a_3=y`3=�����3����<�[f=��ۼ�L� <K�t������ƥ=4�<�M �HԬ��@0��&$<���*��.��*wڼ�n?=���8J6="4;��=�J�<3�=��z����=����4�<�L��ʹ;pS���=�e=w�4<�3�;�I����&�XjI��Q<��=΄���<���<B��!�,s�����)���$�I�)=LD6<�T<gY�=�H4��Q�We9�p�&<jP =Q�f=y� =7��UsR= Jn<�s=o��J=SH�����;���<7�^<�
�2'��Y=��-��dN�t�Z=5��<�o=�z3�(���f�=��0�ϒ�;�X@=!,ټ��W��	q=��<��[��C�47B=��=1 ��>�=��(��F&;�}4<s�0�]S���=	m�:T�U��\��8�{�Gz�<��_�LsA�u�$=�F =�O{�zJ�<�9&��
���k:"�)��$vμ�^3=< :�6�=cT���8�+��À<Ф-<�;���k�WY�<dq#=�Bܼ/=n��h4��s@=�K�;Z5�;=G�=���<֡�<���Ö�뒓9��/�[=�ƌu�n�4��J�9ÛR����P�0�躶����=��<kL�<�m�<���;jЕ�.*ʼ��q����ϐ�u�f=��	����L����D=;�/r<vR?��G�a������<$�<�6=(Vy<T\@=����o��ꦼ#������<o�9-=�ф��h�<劫:<0�q�;�a_9o~q=�6<���<�z<z�:pG�<��>�&h���<�[����=��=Hu����1���R<�;��!7�zh��8�=ODE;�<[ @=��{<`};=�m��V�<F���f�2=,���{�Ϸ$=+�<����AT<)B=P��<D���k�o��������T}<)L����];g���å���<�<s]�<E�:Tz;�� ��&i=cw�<�n�<Ձ7=�԰�m�p��S^��yVK��p=�=_=߰(���%=l{�;퉍<��<,Yr=}E	��jn=fP��2Y�;��p�^�߼��������(����y��E0��VO�Q~�<)z����;��
�? <8�<�ǼΩ�<�m=�E�Ds3=���<�f��!���U�xſ��W���_�4�M��3��[��o��� =�V�m���h� l�<� 4=[�-��Ȃ<�^�Tx�<f9�5wU=��%��h����<�β�>�M��A��?��]_<=$8H=%t�]ꟺ t\���'�wX�<��<r.H�2=���:y��<���=�,�= <�E���;��.�^G�����A��<z��<S��P ��_T�iŴ��X��:���b�<�j�;�`O���!���м�\��ݑ9j�D=�'c�9�~<)�л&?���Լ�"[��P��&�D=)r���`��H=5����u����N��Y��3�<��=?�,=J'���H=�b=3.�<g�`<T��~< X-�!���Ew<�;�<ɈX=ں��.\=JP�c��*F=p6<
l̼M���7���v<%c\=b��̥;��J���=\=ߝs�]3����Z�BM=�+5�����F>;,B<vEټD�f;6��<���<�:I��l��
Z=��`�/Y�e ��=<ݫ����
��
9=�E=3H=>堼q�m=`�6=gc=�<C��0�S��B=����h��7a1���=��6�+�Լ��<���}��<u�<�J=� ���\="h����(=IP��u�)=�A<YQ���(������O�;�dE��_�9�ۏ��<wP=;�j�<��L�Ǭ=�a���eʼ+�+=p>~<;���_軎�;ܛݻ��<3���T�;�
;=��N���2�����?��;�L�<��<í躞���=[��{��ΖB=�A=��=��0<��F����<}홼�B8=p����4<09A=ԧ[=�r�<�:�<}�	=�_��=h���@U�A7<��&=���<�x$�H�t<���h�f	X�����46F�{!�<'垼�Ѷ��{=nGԼN�>��[><!W���=��:`p\��7��eK�V���ż@l��b�<1�>=MZ=p�<�Z!��X�<'��;v��C�=ƴ��\ܼ���m^=Oۻ�����n=��9dd���&��--���j��%ݼ��<�O�<=!Y���G��'�<�4�2k���/�"�J�x�ɻ�n��f"� sM=�}=��c=�fj=�P!=�̼ľ(��>�?�j=����l�ܻ�Ԛ9�WG��M㼥h�z�<b4��i`Y��z"��tE�[��;����v��<A�g=ķ>=T��</�ɼ
��<�	����H���r�u�=j:<5�
��!=��<��[=*��ۊ,� .=R�&���I=���<{/=)xn=��5<��5�<ڳ�;e�;'P����#���<GV�H�J<a=���<�#���=�aq1=m�<O�#�-����*=��<!Wp=��rm=�K
<ւd���e�l�<��<7�Bϻ��ݥ<{rM=S�=<v�1=��=
ٺ� =	���S=�*f;�J���^6��d=@u�<�u��/�<$߻<�cm=A��;� /=�+=��D= �=��6=��r�����k=��ȼ��Y=�>;7ɘ<i3_�U�����_�K[ ���<=�K�<A����<)!5���Ѽ�̀<e�&��}�P�����E���q=´=��R=�P����P<<R=��<b���!]0<�^4��]i�އ=k=��G�9�<�����?�����=P�r���X=\�Ӽ�0=n b��˰<��e���O�/$=YgB�~ػ���<bty<�����;'�*=�Z=���}�I="b=ߦ�;�O�<́�=�$f=�p�<��H��Ԁ����<��;ҕ �(w�<�����7=�7=�w!=��e=��=��D2;:�[������'�<.�a��t~=n<��0�s�;=��~�3=�4ɼl�"=8�8��?=6�;~+����<��9<奉<��o�P�r=CN���"{��S.=���<Yb=��:=l�l=
\k��z�RQ�X���]�u=�̚����"ꦼ���<�"U=V�="��:�锻/�=�$�����<�;�<+pT=L	�9W����f=����c1�<U�ټ�K���[=Q�ֻ�qA=�a="}��f��H�<Lʎ:.�ϻ�
=�9�`l�=�J�?�6��Y<֣��1��<�l:�ݝ��Ѩ;�����;��]��~żB^=���<�Ib���+���<蔙����;��<8|�C����h��o�0����iO� �Ǽv-/��7�� 3=ebּ#�!���W<ś���<�G�Ѣp<�8�=��֕=<E<���<���<Ly�<סp=?��<�y�a
�<`ݻ/'ۼ_:$:D���݀�%C�����4�< F4�E=��:�c(���G�:Bм��<�ϼ����뼼�@�+z���s= �;C���[;!��?@��!�SL=3T�������w���4��:����ƃ=\Ib�|���������a�/����ͼ��X=`%R�����Î��q��&s<Ո!� H<uD�<�+V=�ڡ�N���Q��}�< �\�.�q;��G��I}=�L�<�����C=3
���;h��F�<11�<gs`���?<�lZ�մ��J
��W�J�=�D��mۼj�C���</8���������V=u�=�&�<�v�L��Ɛ���~<lc �| v� �J�-�=~�J�)�<��Ǽ�{���==��<�:�����<[�+��e\n�&녹-�������漂`^�c�=Tb�<�*���)�[L=έN���A=�޼�޹GƧ<�ͧ<.�Y<�ĭ�9��<���<)a;��
��䘻x`=.W=���i�V<��X�����۬<o����q=��<-�<D���a�<0��L�+���B�=*�#�{�a���^(��&�;�<�xw� =ߌ���x^�/���R��z��Z�=˸�;�U�<��=w�9=4]�<��<=��<J1 �I��;+\B��:U��<�F�=��";E]_;���]�����<b=�I����;��Z��d=��;�\1;Ǌ ��!<�>�5�t<�)�:Tu�<��=�2�ZȺTS=X�#=q��<#VR<W ׼�Y�HƼK��9�<�T�0�Z<���<A��o`�'<��M�͖h���<�1�<����O��?=�&=�
!=V��<�k�<A�a�����-[��/�/=u+9=���<�C�j>�< 1=���<�B�n�L��5�=Ҹ�<%*����<��%��h=P� �\|�<rP��b���qA��,��R��?]<0@¼bޏ�y:�t߫<p|;��ȩ9"d==?mo��zi;�?	�4�Z�<�5o=m>�<�;�&�<�=��>��M�=A��2��`�)�u��;g�5=�	I�G�P9c��<t�_�=]~=���<o��鎻���<{�=t%B��<���<�jW=�f���o&=���9R8	�}���<��:a��9��=;�qe�����<!4��dd8�!ͺ�ʱw=hܙ�[=��R�+�h��_�=ը�=v�4=k�W���M;-�%���W<DY=9�n���<��,�$)b=ᶇ;�z<���<#'|��X�<��O<���B�< ^i��n�<ٖ�<��A���^l�9MZ��E	��e=9ڙ�M��=�& �k�2���
=D��<ȳq=�Z=��!=6�S�y<˚ϼq����V�<��E���@=��ڼ� /���E���T;��=�=r�<E�k��@ <�]=Me$=�R�� s���<=����֚=x���B�<~�F=j?p=�����G���s<�o;߁G��\����<�Z1=�k=o�=��g�no==����P�<0�<��	=LI1�:�#�sfH=V S���=��s��� �S����=��f�Ҧ)<FG=gl?=�¯��I�<��`�v`�c�ѻ��O<�H�<����'��$~<�%b=�9C;^�<-1μ��2=��4=�h��ݼ~� ������Ļ�<�a�y=}x,=�Q�<-M�Œ,��Zڼ�6\<�.Q��H<�Oq��qf�*=<�a=H��r)L=㇇�P����!���L���<���<F[J=��I=�9=���=M��1W�$J�7��<E�޼��&�u�0��/X:�,��u��</�S�ߊZ��p�:��<��5�Q6��Z�]x�<k�<~�<���**C=S(��z�g=��C=S�d=U8<�d�$�4�����;e�=����Ϧ���1��<21w�'��;�bA��Q����<!L��N��:��_=���Û=�i�<���Q=�b��<Il켏�Ih���<r�%�I�=C��=�߻W�T��x�<��C����<��<����9�:�Ŕ��Zc<�SY=S�<�a=G�L�W�!=u�<��-�3�:�~�L��<�5J���D<C�=�n�{�;�=h�Z=�yj���v�l��"<R�<5�2��e=	�8��B�=����f|���	�<yϹ�<",=���r_�<D=,�<��j�<Q���I+D=�hO��4���G���<��n�rxi��=7*�<IU;f=���/*�Rw��<��(�,��-����<���1�C�%=ν���_��Z�<��[�=3�=Jʼ�%=���<�V �)�z�]��<�I���(�vyb�2gμqC'=��W��)���
l���=�R.=�]ּ�̊<z`J�{=&�.=�}/=B����-�Ƿ�<�� �>=[��X���>=	_���=m,�<�:L�����<aی<nE�ff��L��9��;�}�"ͼ�cW��=U�;ZM� ��2�i�+��<����d(=g%=�<ќ���p=_Q�<�=2= ()<y��C�<5��<K��<��=�V�<�9��7���;A{�<4"�|���;I=U��<��;�=�n=�!&=B&����.�{�Ǽ���Kw�<�+>�i�=^7�;�G]=��Լ#�"�ȯ=�	�0��Bm<���<��G���F�aM2�U|<e��<p��;7C= oZ��f��&\=��z��G1<�x��^=z�����<�<r\=?��T=�W@�<��<�kv�yO�:�<fu�<��
�}��:=�'z�Kw=TP3<���<�@=�
�<��c��x�;��K����<��#�<���<�tJ=k�ü��G<�&=Ԣ��C5�t7�<��������OI� ��.ǎ��y]���N�T�}���:�3�;�*n���<�q����<=6��N@��M=�a-���<�V�^pr�./�<di�Q�=�.;�%�<g�4=�L�I�=�0����Լ0�==��n��.��	=��μ�^=1Wc=�u=XÁ=9��<�E5��++=#�=�dj<~��<��
��04��6�(d�<�=$��5�;��t<'e	=���<�-�ڌ����&="�=^����]<��ͼ�f�<��8<���<�#�NSH=�A�y�(<�Q_=:�-<,�;9�:��r=N���U=Y�)�h9=�����<��<D���
�6�A�L��<��e=0�[�+q����Y��<�'����:���SC=��<=�k<dGI=�-3<��5=�Sc�������H�B�;0Ka<�>ܼ5R+=�̼����<A���}&=��<V�:=&�ļ�Q�<�%�mZ���5�_���U&=�F���<��	�n9V��{�=�=Lr�կ{<@�*y����ټ�7�
�A=�i����?�M�+�r�����d��K==�
W��˗<q�+=���=ض�<�!n�>�E=�5¼���=0=�<qNo=ݷ�<��=���n^�<��<]��9�&���d<�}"=ڨ��:�c'��?��#�:��I=-ޜ��@�<E �� =���<�l�J[�`�b;��3=I� �~������;�@��r����i=�s=��=uw@�+�<iʼrv%=�7�+f=�F=+G��kXS<�
#<��5�`�Ҽ*�]Gw=~x1=�T�h#=��f��o	���'�1�qy�Y������P�<:�9�H���i�5��;����K=��o=�z���I;*���=[=��T��ƌ����0�P<a��� n_=ŕ��8�=C��=(<�<��<��<�[���<wǳ���<?�<�@&�z�<�'����^��ｼ�ċ�|�<:�</dt=�$B���+=�-��������Ի�X�;E�'��*�<��5��d�x��<&��<��<�����_=���<�U=��>��6"�-:���Ҽ=$=�ռ��@=a_m�D��<�l�<\��<���)9��UO��.�<#=J���;��<���m���8�"ș<L4y�v�<W�����)Y<2,r�Ǖ"��j=;0!=9�Z=<��=���Q+���=�H=x�<=��t�ז =]\e�tXI:�z�<n ����=.����{|�g�ú|n=�]������P=D�*=����<FP���/f0�b�{j�Ľ��^ =,\�=���<��	=��	�%��;@|h�l?�<#b��<�Q����Y��T�<Ww+�wJ+=W/==�a�D+=����&=r�I<�@=H;=��=��<E�=��,�*W����T=�/�@�A;��=�<=fQP;�T����{���4QӼ�o=3�v�@�>�'�<}�<�;�N�J}:=BS(�n������<�=<缕���w黪�9=���;�;;a�;�Uɼ7�����<#_	=�_
</�<�';���T=9�A=��=�ꀻ��0������<��p<�<�l���<��<h�.<�%��.�<�(
^=6p=j�Y��(�N�<��t<-v�g8�<Z÷���,=�G�<��p�q�=�Ϭ��v��}�<�<TW�3���U(� !<q�<�8����<��3=Zs.=xK|���	��q=\�={ ]���a���=�L�<�1¼��;�?����,R�q�g<pj�<-��<�o.=O6O�H���-F�@Ϻ���׼�E=O�<|�>� �<��V=,���Ya��=�<4k��j�����.=�M�<)��<�xh�Z��I���<�Ю<(�<.�����.��G�:D;�<��H�?E5�XF�: ��<��<6�;b�S=��<$�c��ǉ�]�"��/Ǽw�<�_��"�
����<�=�'�H��<Rg��o��Ogs=�Nh=̸<StL��;7\�<��߼HH�=�}�;�'<��<N�������%�=0�=ì=�
=�Y�=�<���»l�==-�+=~
R����<���<0�j=tG=�W;�^&�B�R<1ܼ'��<U�@�)/:�^=�[T��h<3�<�<�ϑ����E��L=�˰<9�9�L��h4޼�����}�E[{<��s<l��;��z<�s��H�H=u��;����8,=�`��9�!=j�H<��<Y��<ȶ*=6�p� �?�o��&�=��*<�&�<t�μ���X�N=S�<���<�o=��4=��Q=H�<|�=R�+;���;��%���;Y�����<���;|��<]�6=]���xȼ̝I=�DQ<b�=��!��Bk�L9�<*v=�#�)����������Y=��Y:	�T=n$@=(�;C�����q������i�T�~�=�t <J�F=Y5�7Vf<y��<s(�CI;(<�zɼs~;�C����D=e��K{�<q�t�ב=4\��4�<)T�ܰt�����#�0
�
�6<x�H=�BP<�Gs��ф�?�^�mɼK~ż���-�=����p����;��=|KR<�t�;�9�<�3K�����,9���1������<ѝƼi�w��[2=9h=��<�#��]c<{�\�I����b��=Eޅ<��л=��B<�ճ�$-=�&��C<��X��
<�*����&=b�Y�F	i�\$@����'�,��C�<�v��3�μ��Ｘ���1ļOj���h�#�k�C�����z�=��=m
���G�`�#=p��;]�;=\�'���@�D))=�pe<�=/��Q=[�o=+���	��=����#;w�S�� �<�h=��i=�	_=գA�j_X�xU�8�F��b`���@���<0=�.=��;�#���ǼQ�&=�G=-�_<��d�a�=�w< ���-;&#����H=�|߼@�<��G��0�<W	����aY��Q��<�g���&�˔E=�<�*	�<�b��F�Y��OB
=E[��a=����g��:ຫ�����``�ģ�<d��==O�<;0*<���<~��<��=c�o���Ӻp?-�6�4=!�ؼ	�t=��;�Y�}��cr��Y���p<_�J=;��Ka`�Q�0=�.=aY=��.=��Iwb�ǗP�4�a=n��<��<&뾼e�!5�<lzؼC�ݺ=�h���<-Qh�� ��̔;�VV�n{6�Y�����=� 	�,j*=�8+�
��� J��9�<��*���&=JEE�2X���E9Շ,=yZ=�P5=):9<r�L�����==�b	=-�!=�#��I��A�<^��<�N�;��.=YU=��C;�j��H��ئ�d�<Q4�<�_:V)����<�
���|.<K�C�a6~�s��@\������`�<�_I=�rY<���޴^��lF=�,a=�?��s��N��G�<:R,�=B=���<Pk�P�<\@<�cW=7м2�=(7m��<�<h������<�L���-���;�r��9<��\<`F�<���<B}<=Μ[<�|~=`-F��=̼¤H<�\?=ǦY=����_=�,E�k��	"���Z=-B�<a0s=�]!����;���<?T\�`ԛ=�lJ=x�+=	΄��[A��H�<I����;�=cf��G���V=_�?=oCL=tH=��=������<�.=�5��,F4��Mh<�B<-#<������<�T�<��C�qW�<��sq��? ���<+����r����Rü��<}3a<ӯ꼠7=�'M�1��E����j1=Y]���,�X��_�?=4dy�ioмV�"��p3=O��<eGf=�N�<lB�e�*���^=)qP�5�E����<Nt���i�W=�9=�y弍��ⱍ�&F=uUi���4=��:����(=.�筗�,�=�x���0�����s-<P\��_�G=��;��=�E=����1�K=$FH=��#<6j<��K<�Ӽav�<�mɼ�z�<�o<��=�HF!=��:��.�De?=��2=���U
�<vn	<�V_=��:K~���G=��,��n<��ټ?ɧ��(¼gwG���U=w���Q=@x��X<Q�~=.��^�#=���1�D<�m�;��K=�k�-=��?�����J�<��&f=T�Y<0����Y=��Hڭ<���z��F��"5�;��<��N=�1N�iߜ<���=j_˼���
0���,;�(��U�<J�%��N:c�<Eş��_�Qh���L�_�V��؝���������º�_4�)y�����;���<	|�5Ǥ<�>���X���=h|��M��;��V=�oW��\=���:��I�<�hk=O������<�e=9M�԰_=oX�Lo=�P�<��G�3�@=I��>!�<n�<cg�:��A=C�<e!�$�d=2?E=�#K��:�=��5=u��<V��;����*�[������E���~��o\��=1_^<�>F=��;_��r�}�54=-,���=K�;�0�=^�7�ه:�I�9Kk�<�C�<�&�<r���ܻ�&&���W�P�ʧ�<q����ȼ��<Υ=�����=Z����\~�~Wx���߻!.޼�UE��Џ��4�!g��<k_����L�qV���9���/=��ּ?j;�/�<J�%;��==�뼅5d<i-��N�F,=)Zo=g�$<�Њ��©<RcF<gY�<(��19� �=������:��B=,�A�'iT�1<=H=�9=/�D��FQ;��B�dp���k��1^�ޗ1�nR<Z=2?Z=�?�<��g;�x�$^����8�:w���R;[b=T�<�6�s�<:�K=���<�@�<�H�{&�<�����;Y
0<����`�<r���h"%���Q=Jr=ծ=xc�I���Y}��D@	<S?=��<�����<��=�Wռ��ּ�<��T�<��R	�<d錼�e�p�"��db���\��&��^R=�=M�J=����q������N=�{=�t��+����<x�J<�}�<9��:J1��%Rz�8X�<�N=f(=��<8�b<�>9�C͔<�p��d�0����<��.;�95�K�e=��1=2�$��U�l�d=	�I�˷0;|ǰ�y�;��u�;J =��R=G�2;n��7��<M�����/<l��<4�==�n����={4�E�=]�<YK��4��<��@� �r���<���n�<��������13��!===؄�D���h��A��jWh=��|=R�<���<B��<�$�[����ȼ��
��tF=�m=z0�<�&=��i�4X*=�~���I<ě�n��<�g��_I��qS<����u�<�!�(Yc=B�;�
=�w2=@�G�h]�<�|v�Z"�;G!�<r��� ��<[sq���!=��0<L���O ��]<��.=�"�<��i���:ɟҼ�e7�k]<��=F=�'����<����W�Z��<PZ�<v�һL�)��>���f����;�c�������y!=�Fs��m=�����<����n=Ѹ =)�#<	�c��6J<�t6=j��<��H�'���+���C=��S=�ϭ�:?=ph:�̧ؼ��<��i�*�<I�*���;�\	E=a�?�l���=$A=H�o�y�/=�A�z5v<��Z�����Ѽ��Ƽ�_ǻ�!F<�T�;��E�Z=-�2=22��߽<Ș��
G�<�<�����d��O�<�Z�<lԎ�/e=�l�x��;K<L���׼L��<A����=ߪ��p(˼{�<��<�p�=z���2>=�B�]�/=�;4=�j����<����[\r=�Z=&;�HV�< s���Wo=�����@�B��;�eB�7�˼;�Ἡ�S����<\�j����/9=�PH�{�4��M	<�՜�}�_�4#��<��ݼ �.�$��� ���<bH�B#�;V#��d�x� '>=���2m��P�9��g=���;�p���_}��J=+~�=�	�<��F��|T�Y�=%*.�XK�(';���#��P*�;��׼�×��G	��<�vV�-��<�����c�-;H�q��[����������7=k���hQF<]�޼�T=�tռ�,�I�5==��q�<�$=�#�l�������w����:=�F	��4~=��d�Ip���_=��ü��)< �H�����EV=~h�|&����L<=O=�(�=�3,�DK0�Y�T=x�-=<���^�D=�b���u��np��U�N0�<w"j��|=;k�;�&�P�S<��D��Ҽ�C=Iq��QJ=�}?���X���S�a`<;�<�d�<bq/��M<^9�<��P�)K㼊7t����"�8�=��<ݙ�^�U���=�ҫ�r~���,A��ܻ[���(��'�=���<5[�<Ed=�S�<f��<��L�t1��x�<:��[GѼ�k�<�h<Oy����P�N=3A���<�����A=)�4��<x����~*���,��� �<������="%�<ө=�b�����<�޲;�f�<��x<M�^�U����X�����~i�H�=��"�����2%=��u�D<GQe�&%-��rI��v��q <\a�¾!<뀼7�w<����!ļW����<8�=����3M�"��;=���;�k�=��=^Vm��2�}����	=�W/���=��ּ�׼g��r9<����Oj��Nf����K�(%B<���;!�ͼ-}r<Ɍ[=?`,���v�p��<����I\=�K���,=�T;K=A��I=����4P=j|��<3�ٸ���Q=e�k�I�Q=d]����f�pr�����^=����p"�?��<�
���J��{y=&�f<���r�ӼÛ�<L=+�=���i(�<��m�k�w=���:�f=Cl&=8bC=hD=�Ù;��!@����=�Z;=���<Uj���%�=�9=Y |�[��\�����xd��+������T�%B]�oAm<ng3=\���7U�;MP��Jt<bX�<nP�;|�<��#=��g��:!�ʈI�Hf�H=~(9��!��k�=�Zy=4fI����<"�<���w��:#��G~N�dD�<���O��F=p�ɒF;_��<ש��A <@J��)g�<�p=��g�C8=�:�<|��:4'�<J�����<=�;����7U�'j�<��8��
=��ʼS���y���7<��;L\����<�kO�#�.=��һg���G�����&��a~���g��Q���f=��<�9%�����a����;2����b��R<=��9=����$�09gR(��H��r)�3�=L�R=�z <ґ/;�AF=�jn=$�N��'�":���6�H;=�n]��ι����<J�G=�ۅ<(O4=^��<aQ3=w��:�8Ƽ�0d:��B�b~@=oi=�{}���<`��ۘ��Z�(;}J$��8Z=�R�;�PZ���E����<5Ƅ<r�=��<ɂ6<��s=P)s=��<|�N�^P'=T�=�2[��7=�i�<)X�|ȥ�1%�$J �_�O�B�����c=��m=�:N�i<��5<����v�+=�fu=�Q=Ѷ(<a�p�n�ȼ8et=�N(��z'=T�=Ų�;��K��<�������/����}<<�Y�<�w��L�*�}�i���f=�eY��'��:�<��=��N;~ݻ~^%<������<�g���̺u�S�� ���ڼ�v)�[����)<AM��Eŧ�'����)=�咼E�;��0�笧��	źq:=rԣ<��(<��<�p��:=��=f6]�L[R=��<�:̼�e��X��F=�OX=�=U�d�BR�RY<��f=�N�'�`;��S=�%�;W��:y8���R�<.#�y���'��h;e�2�C=/���A���Y＆sz<��	=�|���?@;@�@�=��0=��l=���l�=gZ5=�@�<kPK����<�E׼I�+���I�s��<�A�<A2���N<��<��=��#;�ڪ�jh=0j�<�*=>G��
�<W�$����<���;�F�<0��=�^1��'=T�J��=C�<�a%�ȎԻ�#�<�<�d]=9�ݠ,���=ޒ���L���V^:��,�cY;dg=��L=ܤo=�G<Yx_��8=[��9=��J=o�=b�c��>���.<�,t<�.�.L���f?=&㥼�����D������_=�ހ=h߼.�O=w�"�ݘ�<��/=knV=H�Q�Sf7==�ջi�*�7}=����<7�;��a=�k�[����ۼ��"�啻�Jv��>�	N=��<`��<���<��6��`=�E=�\�<��G=�%b���t�;�9@�1A~��>��+�V񫻻�9�,�9��l�j��`��=r�"D*<�ڵ<)C�9����B|���R=�ȼّ=�$H��O���=:w<�e�<�O=.���<��9�{;�I=�H=e�=�{�<�n�<U_$=����*�"�{<�p=${I=:�<�>�<d-ɼ8uӼN@�;~}��ͻ�!��	�<�.��v=U�^��zs=//��ԔO<ف��(I�<n2����j��;"��=�u<��<��3=��F=7/=k<�^=��9��<����L�$=����|/����>n �����\0�
��<���<�ؚ��$==�Ի�	W�߻��n�м�悽�)��)=7�9=�;�^,X�'����p�|��;s쪼,�Ѽ������:>`��P�:��+��=Gq�:�軅I{<\�}��D�<��="'=��!�R<�~��'=��<�!���<��Z�'�<����<��	�a��+���}�B�<�=���< BZ=��&������!���&��Q=����Ӽ�=�Ƹ������PZ�I��<���<�W)=O	n��tܼ��j=�w��X���E��Os�<7.3�!��<�a�;S{%��_V=`��'���z��3����<��+=��=ó9<؜k<m�޼���<�3�;�L=,[�<��
�g�3��n=��d<��/=�YW<A���|�o�<3V<2=�d�������g*�;�;�B� =s=����"���)=]`6����Lߐ��N�<�5,�Y�?=�j�<���<+;�V���<���<:ሼ���<��_���&<�=�:]=N,0���5=tC"���˼7Nm����]07=s��=��"��FF=rȼ
Ɠ���/;+�D=P1=�J%�i�Ӽ֮�������mL���<|T׻vi��e� ����<�b�<�`�<�ޚ=�⼅R�<���������Z)@;�����;�`i;Pc:<y�<���<zգ�������<\��:@�6�< �=��=���@����<R��<���?��]=ȯҼ�&*;����W���Z����<<I�<X�|�����:<3qX;�J ����x�6�Z�ּ_�&�=~P=EF=�.@=�u���<�Õ��q����<�G=B!<�\�+��Ŵa<�q��;CR�[W4��et=Npm<�߻6S���f��#�<�}��Ap0=F/�a�T=v����<@C��_N=nƼ��8<"$<������=h�&=lF�#w�hݏ���;��\�
��id�
7%���R=�ؔ��V	�n���&v�%�/=C]���<M<A�T=�a��]9�3uS��-f=RS���}=JM��� �<d2�:��¼�x� �-��<U�����~��+�<=^���]�=�t���`b;�~�<e�;}<�s�֨G=[v�<h�/�^�'=g��;$���c�Ѽ�J���=4��<�3���qU=�\���:�<����<�Y���c=��.������F�L�B���o=�T�a���U9=�'�;��2�R����7��|^�^�^=��~���v��J�<'p=޳�<�/i���v=7�-��ۢ;�*�(�5uF=��<�E�<~_Q�|�m{������A��Ӽ��	��J�<��̼�iԼ�+�;�N��;�<|��<ً�����2����b�!;UL�����8:=�/9s��F���&���O��<X�5�
;�
� ���:�d�=�d<*��m9=��	=�.%=@B�<_�;���<c�v=CG,�kn�;�>��u;<�ɼ?���S��e��;���<N:X����w�E<��ٻ`Ru��tX��Գ����<��&=�tO�2��l;O��+o<a�A����<�'�<������+9?�7=��I<�o�����߻�����_I�Q*P=|�'�G�=:��
�<E�U�3��N=b2=8�<��<՚<�a�Év=`H����<%�O���������K=070=�=k���8��<�3����<� ���f=�<��=P�d��~���B��ټZPb�e�#=� ���
E�� �_Z1=��<k+��ސ<��u<F~=���<��==*���;q����89�<�;�W��������<�T����S6|�����=��D�2D=9p��7=x�<R =��C=b��=�[}=��i=��(��Vr=�1�<�\���1��>B=HΎ=f�<����<�U��˲�=�Y��Da�Sxc�
s=��6;B�ӼX�b=���<��;=�W��w!=�As�W�\�W��<�X=X�=�T-�O�<���<w9�<r
H<�lؼ���
�O=�l�<��X='?E�W�Ǽ_��g�<\W*==� �<� �Y��<�M�<�5�<LH� /����p�N:&<d�ͻ8���8}�\d�Ȩ��}�tA=��:�;<jӼ�G1=�#X��8�<ĉ��̲+=|	L�{=�U!=��"=��<3��<&I�<%�<�D�;*�<]�o<���<�6s��u���<�;v��VY�'�;=�����lf�e/x����<���<yD�<5��<g<=��㼝=���;��;�	G=�4����<���<]�N<"ŀ�����K��QV<9�~��â<�0L=WH%�9�E=A��<`'H=L����=5=\)
=�i�<Rƕ�e��<�8%={�M���g�3�;q�o�W1�<^I���"=+X��Hx5�YY�9�<��P=�}����B=����m9=R� ��m����<�$=w����#J��z��"1<�ly�\͆;��=k�v�_����Q�<��M=�J <�o�<\+˼&Ј��G��S�<"��<�&��CC�<�R�N�<o��<�h�<5���`��<��V�S��<7l��d{�2mg�Y7�O�:�`t�8(F��8��d<9%"=�E�����<��<=T��:|59�8�.�=P�<W6="��;p��<��J��(�;n���e&=6@|<_�bۅ��5< ����:bjZ���Y��:<� ����޼��3�db�<N�J=��;�F=+��<�&
='�==F�;_��)<V=�r,�x��<�J*��H��W�<�Y{�CK�<m��b�nB뼚�=2��O_c��B+��`
=W�o=D�ڻ�/;=:�&�����Z�U�&��
=�9H�[@>��튼ϻ�I}E�����.V�cu��Q7���.=��<U
�����O����̼�!A�&������7=�G=�^�<t�<�{k��v���l<�����D����S���)
6�)Y3��]<�g<&gL�|���͝��	$���=>�p;�񁼰;D=�� =6�༃��blh=�2T<`K=rK=�%)�~G��S�[�O7.=;�P=��+=h�W����Ev�)7%<m��<WF�U��0�+=yZ�蝦�|�"<:��;f�$��wZ=�-=��;��<ި@=lo�<�L<�`�aY"<P@G=k�<~M�|���SG5����;ޟU��'�OG&�j~	����mP��J)<�͡<`Yd=�%<���
֚:�sz=[����!<H�J=�S>�ʌ�;���E;U�ּ�W�;�`5��N=��<��P��ȁ���<�7�� S<]Fp:!=�I��)��lټii��m=O �Qs�;��< r$�u��F�C=(��8���<=eJ��2x��盼)=ӼN
�<���PE�<{���ϒ��j)==RU<��v���c=GN�;d�C=�U=B/ =R�1<������ӻ���<����OL="�<�j�<dtL�SU�s���i�$<l�y�n;y<F샼�:c47�F��=��=��=�%4�6sR=g�P����w_����1���ڼ�������;V���O��:��OL��<z�~��Z�;m
��F=m����;SE1=dj=��;|��B��R�+u��(������<�!/�tɹ�x�^�y��;�4�0f9=�P3=?U��K{�q>�:谽;���A��&�U=����"{<��g�:�3�=���=��<����b<��(=��Y=�ϼ�L�<��l=�"=�F�g"R=SƼ�,<k0!���������x=b|=�3�<ݕ =��<�>�<�+4�_�&�['T=6z:���6<j�<�>�<|ed��q@��?��U�(=Z�<C��<�.�<�Sg=�6+=�_=b@4��zk=�78��1=�j<yV�{���W�$�,Xj��j9�ҽ<�8�=%1<���<p��9Г��r��`!��0�;BK��z'=��C!�''n<�K׼�x-=�E0��?������=�Z1�f=�;J}�<0G�<�$M��û���y�G�<��V�.0u��޵;.P���V/��ݻ28(�-�0�"b�]�=�4=��=������<��u;AD��(|$<O�t=�b<B��<�}$<;�<�0h<-�;P�=\�,�i����Be��}�<B�U=C���GX�\��<&V�#����U�=u���l5�$K���2;�n<'<�<��g����<o��<F͘;"�޼��B=@nW=�?=��==�'=8�{���A=KG5<�V�<��;=�ǻ"�F��9�v�)��`j���A=�伴#�<���;>ye�����\G�|0�<7s�=�����o=-M��[i<qa)�,�U��=¿�{�:�V����� =>�I=�;:3�9=�����=e秼e���<z'���6M;>��+v�05���<�0ռ�����<�w�<�V`=�Q{��I�<jn~����(��=>r`<=��μ�|==�%}D=���<;�d�k�D�޵i�;׽;��;��<@�`�99�8Y�>�J<g7�^���/���U��N(=�'�;�j�<�X%=B.=�#=�6=.Nl<�1V�T�=�s�b=T%)<�\�$����Y=�N�za+��q�9�����<��=�;�<�GL��B?<��ݻ��2=!�0=��~���1=F��|�����=�{�;�hC=�7s=���HE���K,�2L�<�Os��gz<WX8��C=���kE˼�V<)�;��i=??g�c-;f4G�7��<��;GG�_��<BKf�2�O=�-=u��$�'�)�b��E<�s�=v\=�=M��.������_�6������1=�p�d�n�:���R=����f׺8����߰<vJ�]�A���h=m���t��-<]t�=C=�<�*��u=ʋ���f�ь����<d�
�`�[=�<�Pu�<��}��;?��=�;*̉�=��<�&=���:l�h=�%�<�=v��<�s�<�~��wp�=D,<��b=Pؒ���=�yD8@�
<L�<�����W���<�e���S���J%`:�z�;/�c=*ځ<,n�<d��{=������==�E5��z��;�w<���<���< ��<��.=-�F=�}?=�Zi=@x��<��P=&L�-pw���<�9=*� <��/=6<=��R���("=�6;r3={�]<I4=�m=�<�/�;�s]��(���)�r2=O�=fL�;Xv���:�<�$=^="�;�T�<�d�XQ9=7 [=ێ=�q�ᄐ<�:�<#��;P
=��<��@�42a<�O=TJu�@Y(=�=h�<G�3=��9=IӼbE���)��$��ݟ<羂��7=mJ=� ���xg�.g�<:=9!=�W=/P(<�G=����o�;��10�<����z ���-=�P��AI=h ��ׄ;�d=&V=�p�<�"9=�4�YU�<�<�:==
)T=]�^�2��e]�q `<"�I=Ee=�%�;���<��;���z<�蜼�L*���=<��(�����Z=��H�2�'�-H�a�H��b0���ؼ� �wW���AC���P=�����<�l�;}�=�U=�	��,.�
r��)]���d:�p=hf=����G�L=�Nd�_��<\	==cM����*��T=��)���
�L=2�ּ���<�":�Ts<_���(�;�#���kɼ븶��?�<b*<�P����<�ͅ�ƺ8:�S���dA<�<��<=)�L� A=Dn[���=�*$ȼX"���$�C�i��D���.=�i<H;���==3�=���*J�<�=�x=�|��=!b1<����<]�=��Z=���<ˣ=�I4�ż�GIռ		���$<�l���%�;P�N���@��<=��c��!�<6=�!���A<�n$���b��;=�V¼
k�;��=�(�<��<�,���<����*,8�C�=��dǻ�t�O�<�>=W���ڿ�B�-��f��!�<�s�;�Gμ�(��V[~=�gN=�==VC�B�:�n��[�g�u�-�Y١��輴}=�=Q|��ݼ2K�@�>������jf;;$�XK�y��Oh=�z�<}Y�<��P=,��Ν\���v\<�����=�G�����<�o<�>0<|Ԍ����R~�<"D$�ݻۼ���<���1=8�?���a;�.�<�)@�@�(=h�ԼV�q<��=�au�� �<`�������Q>=� �<� =eּD�$���?�)Q�:?�<݇�<W#P<2���h����X�=�<�򷹕>��/����ŏ�li<��~-�<�)c�V��:f�G��W���ړ���3�h�;��8[=;q�����<�>���3=�U��b(�y��~�<%D�<P	���4�cKX�ژ�Ka�<�F=lq����;V|��6!=!�,��7+=H
��}@� 3�z|>��s�<5Y&=E.^��Ӻ=k�<�'<["=�l]=f>�i>�;��n<{���G�<�-e=w� 	�b�o;��=���,�<�EM��0��B:=ka��{�<�4�	|�eo!���Q�$�ۻ�ޗ;�ީ��n=N�Q�c)=�fP��H�<*�F�������<��0=FH�<ŝ=Ze;�5�<��;��V��6R���=U�`�<��T���<	�/�f�1� �n�Ռ�<�1E���K=��Q;cូKg=��_��eg�jp�I���YC��@w�<�뽼�k��	��b[���M=��M=�,r�x!1=��=����i8= L=픽����A=�|g;~+��F<��P��+L?��14=��<O=<����c=^gv<069�5FŻ�b���0=ۋ�&9d=j�B��V<|�Z����=�r=���=�=�G�<�*�g�9�69=f���}�q<B�U��=��(���d<��R�G�V=�z���ȼ+�<V =��D<~�=ˬ#�ؑs=<�2�ҧ�<+i�=��<x �M�һ]���q<=6������=�3F��U~��Sp<�@����<�rO�e��;)ZA=�\\=��R�t�w�G�;;Yȼ��:��DO����5J����;-�#��5�����PI��$=�[����&ڻ�f�S=]F<v���~{���
�.�
�=qȵ<t��;ã�O��;:jM�D#=�A=k���d=��:�����"��ZZ��� ��P<WJ�<ް�g�F���v��J�����U�S��<��Ƽ��>=���<��X=�b<f=޶N�2b=d�<��F=��8��$=���[<nM��k�+�q�<D�~=Cc<���<��O���:t�/=��t<X:#=X��:���
:��aE=�yT��� ;��z<.=�����.�>��<ym��*=�2q=�,�u!t�|=Z:�=ڙ=�lV��!R��-=��]=T1=)��<�t���<%����.:�M�<���}�����𼬜A<��B�Ӽ�F9<%&X��V:=N���f=�ӹE}8��}ӻ�J=�h�<�57�0K����x���<wLn<����K!�̗O������4���>���_�@���.�Q~��,�=�޶=[D�دq�h�G;q����O�-n�(��<|J=:�ϼv�7=T���7�6%���<Y��)�=r3�*~�ܬ��hA=��=��w�T�U=Fzȼ'�_=7�}����<�-=W�<ݺ��OY�y8�<��=V"� =F�<P�C�Z�H=�,���</�D��幼�v=��<C����<p���Y���Z�<E���ށ��T��?����d��= ��Z��d%Q<9ɶ��V&=�t���=��$���5=�I��Õ=-S���m���5X<��C=��-��� �/�9�������E�箼���<�j=��=f�Ɵ�1c�Pn�;R�<�r���'K=��=h�?����9GE��r����R=�<"������<�����=���[Ȳ�x/�sd1��bC=�"���C^=�^;=�P2=	0�<�d�����<ew�(+=� H��#��(��<�,�v�r @�u�=7_����<F��<���=4�z�s`�<��*��=:=2흼ǡ`�8�=
�ue�;],X�Ne*:��2=!�b<�%�<���<[�"=G���b%=�s!�
#<�+Y=���%�=���<��ɼ�=������o���m={ �<��<J�H��i=B<�[0=�W���&�^�=}�%=�I��5�<�;s3X��ׅ</�P���<�/�����c=vGO=C�f;��$=0Qb<|6<�㖼�@��ީ����A�ȁ =�g<qlλ!Z�y�I��'-:�:��P�߭,��`f=�
=WD�<��2&���=�.M����<o)=� ���d��<��˼���=�m�����џ<��������@�<��A=��)�J:����(�j<mV�<��O�mXv�q��<J8�;���<v!H�W��w��<��!=['�z;c�<TS*=��
<�`�z悼�{,��޼�-�p�.�CWJ=���;��8�h���-�C�;�G;@�!<ZO�=#	=Gx=׎H�9���J�;���<�]B�V�<�"���<���<	��=��C=El���I�k :��9<=�����&^��zO=����#�n<2JQ=M7d=l��-y��j%a��H=��<J
]��\�<ď2=		=�%v�6�ISB=�Ma��<��=�&<H�<+Ճ��%1=�}T<�u=j�,=��,C�]�|���=��O��$=]B�;�i=�������"�;�3>�ScS��ް:�,��ȓ��8�i�@=ۑS<�<~�~��Ã<�x<ϳ)��A�((=�k;��;�<1a��A=v<;һ<"�����Q�ȼ���<+�i��_�<G%(=3?�t����5~��Ŝ<��A��:��{�P=�m;�
:^<���<��F=�	]�0�(<p��<66=�ӊ<w)�Fㄼc=��׋��A$=$��< /���A�{�J�޾�����H�S=>��;Ai�k?�<��f��S6�;;aȼ6-`�F�^=I(
��N�=�Nr��<"X��T�<N����k�<J��	�f;�Ԛ��k�=~�R�k�x=Y�H=��ے!=nc*<ڃ�<��'��bb�� e<�t=4v��i�<�^"�u�e=�����O����R<�ı<��*��W�:=؁=����<J=�=(�h=�:m<Te=\�����<��M=߸_�}x���x��\<jw��
�;��L:��>=��8���E��<�9[<(9�<	�=����3-�;�;;j�=
d���ʳ<�k=¯����=	�b����<+k;�xC<	i�;EA'=�[�<	SY=��=��=�,�ňQ=Q~z�@i���<,�;%!�<R�<��v�g�Q<�<��3=�ʼ��=����<�����pA���=5_�:\�<�����:���=�:=j&¼m�=}����$V�#�=�6=���<3+�<a�_�̓U��=q;ߓ6����t�==(���ɼ9����R=la��%^��������/���!=cB�;R_/�k�=����B�<s�b<�o<B-E=~@�����J:���<��<T���(=��=2�=�o��d�=��S:�O3=�A=jV�<rw�坌����p�N���<֫�:��Ӽ�+��)�Ȼ�P�/��<�|���L;���;��<�ٻ|qg���<�#�B�c�t��>F<8��;I�,=Wt��e<�g<!�S=�.;�Pʺ
^�i+�=|�ټ���<�bR���f���=��]<�μ⑅��@=�=J���`[�<�[=�39=�}�3D[=���D��jr=�T7<�:;�X���<��N=?�h��m=>�;�ﴼ�}	��U�Wn<����"�<3��;��y<N�Q������Hd=�a=�F�́��6ǧ��R�����a<���<�!��Ԫ9�M� =C{$=�o�<Fj@�n΄;��='$�R=<�피x�<��s��Ҷ::�)=q��%��=�ξ<ƀt�܍�D�b<�K_=C��;p�A;>6����=��=�����	���T=A�=إF=�#��./=�j��?��8k�ּ�U��u/<'w�<��*��/�<��G=�(�<��i�è;=x	4�cT�<����G=Z�m�9r=�#��gt�%}=���a�<��Z�W2���9?<�u�<��=�90=`��;�k���g�VA�<�C�KJI���<�$��9.:!����<�NF=$�<]Fռ��]<��<���<ܕ纕��;���<zG���������+��x�;��ܼ�n<�M�=w{W=��=�?�o�7������1=��U�z�\�g[<�;#=�%g��L\�Y16=A� �@M=��G<�F��Fj�ui�=7�&<��)=r��;]�����<�������k����Dc<���������y�X�=���C:q��6��cu��-�=��1<�E2=�6\�F�ɼΨɼ�p����;��R=b��<�F�S=N1X=��r���~�>:�$ϼ�=`ݗ<�Nl=.*=�¼t���9ż�y5��V�(V�s</G�rz�>��<�ɼ�=5Rz<:_w��$@=�,L=W9^� �x����n�<~����Ns=�+�e�;H�Իv��<R���rɼv߫��Y\�^�?=�x��I��ZP=~�g�e_h�����<A��U	6��A�<NH
�rk,��=F5H;�	/=6}�<�8�<u��xnU�JZ�^���j<��?���<���U���+b��v:�5=\���|����Z����P=�D�<�fL�".K���;�E=Hg]<�����<�<���<�F0��+���Y<dq#=��<(ݵ��B��RT��=$L=��¼-Q_=�U�<r�<�����٭;(�s��A��f]�=�1�<!��&�l=qE�|�;<�i=~|�����R�̉��
Sܼ��D��3�<�l�<��<�%;��$=��N=�S(=�D����< �O=�X��<�=��l<"6ּ��.����`=���<�
=2�q�s����Cy<���]�f�.[=]<�<�����u��?k���<��&����<�\�92O=�+V=Ľb�F!;P#=��]Q =e$=��-;��ыy��[~�%c=�1Ѽ7E���(p��%:���H�2ܰ<{+T����<�����s�1��b=Xw�<oCH��'=��r��\�<�F)=�]'=�_k<�����|l�[X�=�,�<���<Q�Y����:�&ռ��ܼ��;��<���:'v�;{H���������5�<eE��D=�G=P����=`*��׉��������#�=�B�=�L=�: =urV=�*0= �=夤��_�<h�z=U��;�5�<*��9so8�Gd�<�߼T�=�3=,��<��;=�P=/H<�v=���:�/��$?���s����9*p��n�;f�@�nQ���7?�;��<}f�;zX�UR����*:�U3��5��3�<��?�0./=�4=u�ɼ�t?<�t6��`���=*=�us=/=�q�R��<�9ʼ w=AS�;s��+�����軹�*=�Q*;�S��}<{W���^=C�c=�g�c=/���1=�W�����=Lj=��<��=�0<��=A������OR�[[=���>���)U��=���<2hV�f���{���fa��
]�E����i�<6��[5=��1����==��<<�I����;ﳭ:��<s㜻�IR=n'�<�n��7�r��<������I=�=ü��b=`�;���<L�=��켸R=�p=�X��8��<�����<A��<�z:=]�X;��|���-=�4y=[=���y۲<�$<�"=��;�[G�Z7H�������vNk�,��T=���C={,���=.���w�=�/=�/w�k�R���\���E<��G��A?���$���⺖a$� �m�L�&����*0=x�x��a&=zeM��d�<�/h��;=�0.=rmf=Pє�����/ϼ�-��u�<��<��G�#��8���0=D�＋�Z�!�;;�S=�&���z�<�K��4����=m�q<bΜ��=��>�,2�<�gU=_1�;�'=���<�1���1�!��=Sb����a�ҁƼe�<2�<��u���<��R��2&�x�m=�5�\�+��q>=�E��Š<���<n�1<\�k��ػ��λ����<�ț<��H�O����n���+����<��=�����q�ú<��d=PH��v�ݑ��~8�B)�<��5���:���<�Y�TH����t�<�.<i��<� ߼��3=T�R=�i=��5�Ɛ!�1�����r<i�Z��L<�)����c<�q7=&��<�b���'�;o��w��2�ǔf<�<b=�)���	)=��;<KF������s��B!ڼ�Iy�E�ͺ�.=��r;?�/��[m:����;W�;#��g�g<��j=�`�5�;g��<�'g=��BhO<-s���<R�=�Xϼ�P������u����?=	��΢�(���u�<��N�3ଽ��'<AvH<�}��a	=���<�%��(���a�1C��$�A��XU��Yȼ�(��-s���Z�J�*=�@H���|��t�<��Y�C�<�=��3=4�k=���_�<��<	2�<���<9�8��=3L=Q;4�v=y�	=h9	=X51=!O/�la;�w���<��M<��</t�.��=����� =_����-e�z\!<&+=���վh=L�@=��{���8=y��;��=��>�<R�ʼG�.=�j=O$='=F���Ն=*_S<�Y:��B�Sy}<9==+2�<MC�<3j���=�iK��` ���=�;�/�;:Aʼ|��iE=/ܯ�9���$=p̼.�XBy=���<���:�F�<_R�<B'�<�#��4�ί�<�?�������  =��<M����4����F�X�2=A�3;����U�'��9=�a=ַz=`�B���]=Я��n�<��<_v�:˰==w=�$�<�7U�AQu<*�,=F��ҝ��a
;p=>=b>�����<���<��<�I��B5=/�_=p�������=+�j=��C;P�?<��ɻ��Z<fY<�%=r�0����<}o=J��	@��(=�x:��»��<%� ��U=b�ּ<�K=4�<0���ك�=[Cr=�n�h���'�<n����;�/;�BP=� O=��@=48l=i�;���x����<��м�JM='=m�.�K�=�Բ=���<��K=y�k���L<8P|<�ki�;�l<B_����;���R�D��o��0=�.=*l�<mT<{��	���,����Y=Uco����;��w�E�N�+:��.�����˜缴��<�D=��)��]�<#�=�<+�O��9(=�ǎ����i��n�
��%����]<h~�<�!���=��Ǽ�����:���;`@��ni�m9,��a��z:=p�?<;����!�<b��<���<t�;~ +��䒽ޥ�<�ҁ=s<U��<��P<�=~���K�<�0�������$�<�M�<5�<��[��o)��Y\<����]�(=-�<��J��l<�!;E��<�����a�L=ЕL=�N=�6�<q��;�� ��{X���Z��q�=0	��T��;h��<�=���<�~<,��6�X=�=��=��#���=\���FX�<���<�4�����<_s6�s\<��_�Ni�;>J<�؉;��\=D�4����<��!=kRټ-5�}��<�U�X=�P>��F�YƋ<e�$=�C�#�&�z�_� �-���;~h�<D�.��T���*=|�ļ�����U8=��+<gbS��<�#;�d�)E=W_����=����;����"�=�==���a�:1�˼�(̼��8�Uo��3��<팉����;﯑;۩n=�{0<s��^Q�UB���M=k��B����3���W=��L���A=3�I�Ì;r����p`���ڼ��s=
-�<7Lؼ��=�{��g�Q��z\=C�T�.e伤�=5=��;����1<���^�1�c�8��*D=&�C�Q�ڼ`�ȼc�<#�߻(ȅ�3V�<��"=�����A<6��{�N��B-=�AL��7M=�}�x���ID�
=�ܷ<2<���L�W~*=�L�<�b�~�=�ul��G�G�����U=�=��,=?p<��ǆ)=�|�=�=�����#=f����<B�((� ѕ<jDٻAMb�:���Ҍu=�h0= b1;��<�*�F�<C�H�
g�<�h =�ϼ<4���M������	<�{6<���; QT��-Z=��;���'=�4=�_���H!�:�^���=��C�<n]�$�m���n;6�&<����أ�=	��<ne_=�&�8K#='���d�;2�U�����*ʫ;�=. :;� _� �OD��n�<�ٷ�< Lm����<H.[<�DA=�I�=��^<)�ռsE=����VEF=�v�<�N=A��%�=�q!<��h���8��v���9��bT=�2X���Z<���<^๼'?�<��<�m!�>b=���;���[�^�&�{<�L���dX�q���= ��Fc<%s��MZ9���<�~���u=��=�5ʼ3`2�r/=�8=�0��.���4���$�G�Z=.D2=R5��$��d=���-C;4�1<�9}<	q<7�H���<��>�<^v<�ۉ=w�?���
��o=��伤�
���=6�ҼUD��lh;OvW=7P�<7Z`�.Hp��D#���7�R�9��<@f�<��!=���<*�*�F�,=��c���w��SV�_^`��kU<�,�;_?d�.D������ϼ� =��i������]'���<=���<Kcr�q��<=hn�<��<�Q[�-bG�a��U� ��֪;x ����O=��e�H���(k�!��g�<��=>Ih;M�=�,V<C��Jx=;�;��!= o=��:��/_�3#W�tG,�N��<ř6=�r�<�P�@� =�h	<
\��j��c=.EM<�Vb��X���U���fF=^v�}޼z�<�k<��;�;�v�K�$��L�H�&�G�T�)�<5����F:�:�;��,=
7��*<�qj<��<և=�\��h,�%gw��|�����v]=7�{���<�%�(�<�B.9m��Y�����:u]��gA����<%X��r�<�6��/�:�#�J��мKp:�Ѥ<螼D@!<�%<EU��C9M<gX��mQ=�<~tc=��{=?�5���e��5 <��J�>��;�`Ҽ�l_=6����h���w��Q��HD)��=�vl=t�P=ۡ(=fA0<�A�=�h*�UK�:�l���t�S~<=�W0��Q��Y�����<���hղ��I<�c��H;=Y"=�K���=�</�H�=`�h��$��|6��b���/=��I����F���=���i,	�i�+��Z�<>:<�E	<SU���)=�Vn=xe�6�;�3m��Gv=�y���>;
�/=�V'�4�j;�0���8=p�.<�2\�F�}�#�_;�Z<���)~�<'��<7�\:.��<1Y!�v�6��x�;��3<"s�[�=��3��<t��ƑQ=,�=Nd�<S'=
[t;�+2��O==�J�=b"���¼Ni�<��<�Q��T-~���D��d��u�;g�w�v�D<Yv~�T�9���:�c<��	��g�9�[���޻u^{�_%��y�Q=:�����s����V<����5�Y<o=��O=k�S=��C���J=6�O�G&=vN���N=u�(=J����k=_&=F`�V�.=j�=�"��:��y2;�7Q���ɼ���<d��9"������<�8"�.B����4�;$S=@�=���G{V���{��oP=# �4�x����5��<�N�=V6/=��=�g�p�%�=�/��#<��H����S=�J�<�����2O�=�;>E�n�5��V�Iu�?�=��<�"�;�zU=v�[<�/�;3�<��M�`��*�R�����4=Qd<H�}<��O=�Z��v��?v'=�y�<����6=4W��=��Rj��&�=c
=y>;5��;.�f=���<>�+=au��r=�R=���:I���yQ=Z�B=�I`=��;Կa��i/=`s�Z&T=�d����l��<�)`y;)Ǽ�\4<0���޼C������<�o��1��ٷ�90�<�N=AV���5�# =�*�8&��g�_=�/=�;��Xz<�9���=��n�x	;��U<�q3���5���û� �Ml8�L;�X�<<$�Լ�P�<����v<�i��_ ���#���=4!<|�<XLB��&e��zջ6	��b_�W�s�w�E=Y4M<lʼ�@���:�������<Qͼݰ�<-9N=~4���H=��
u�<m���d-���O=�#=��_�@�C���мRVs��-����d��ԝ�Q�<:����,b<ى�<��N=��7�;|���I�<��$�"=(�(#H=�w���>�T�[=K2=;3���C=�󾼣�;p=p p�لR�px<�:z��@;;a���5/�<V�i=�L	=���E<���;9 <Fq=Je=n]�xZ��OJw��j�/$3�%<����T=�g�H�<� $��(i=��<�_�<�B7���5;���Rؖ<*�=x2F=}��:�Bf��9]<2a'=_����5�G��<F�׼�;�
�6;�=��]=I��<�<rx'�D�XCy�o:=僩�l�=��I=;�)�:L���=>3��s�����u��*�-�E�/=�IA��i'=m�<���<�WI=�ļ��;ŋ2=�G<)����=f4缋Ɖ:L�<�<*<7�W����<XO���<��"�N�F=N����q�����@=�����	=��$��g=DG�<H}:�3��;Y�G��-F�݆p��d�<,�\=)@���o;=�%�1�<���`<K,ȼ��=�t��̟<��%=�6��ݭx=C
7=��9=�8[�lNA=��M�DӸ<����"=n}���	�<���Yb�A8=�=ɾ��-���$<�+�zz�̟�<Q:=9w=唲<�<�<��า��;.{�p�=xo=�*�����<,�輈���=�}j;!?@�sI'=c�Y=I�=�f.=��׼��ߗ�L�A<S�=�g��(d=����=��}=+=Y�f��:<h�#�����6Ɗ��%=���d���ȼ��`=�y-��YR�hAq��4⼄ ��	�!=�s��P<��{!=��#�]��u =�(�<-=eA%<�Ru=��8q�����<�}K=�m�<~y1=��t=��E�4�<
|L:��{=� /=G�<y�h�2u=PF���xo���9=�nl�q$`�>�&�E����;;�0�w%7<4�*�X��J���Š;�)/=��N:���vF<_��V2[��A<1G���j<_d��++�0�M��v=^���� ;@g=����
\��@=)༗ż�Z�l��y�I�?�m=��K<�*l�q�=�<f��<�K�CiT=|d�� =	��3��<^�*��@��A�S���R= �˻���;���
�B=]]=��<�=D�;������y������1�3�=��ƼW�-�"h<B��<J�#�e = +=?�˹;�1�;b� �H�<�p4��;u��<}�B�j�o��h?��?*=�l�D;=eq <�I���,=8׋<w~Լ�&�4��<�O1�@6D�� P�zǾ�j^�f�m�*MP��&	=0Da=ƣQ=��o�qɼ��;��@�I�?=���(�j;�!ĺ-���%=A�l=Րһ�jE=
�|��"=1�+���*�r����ݻ�V[�b�:��,�z=�hܼ��1���<=��S��?=�K�Y�< ,����F=�Y<
�<e>�:R94��=�]v>�2E�<) ۼ�)\��Kr=��`<�=�2�Ζ<"N�<?��<�M�9�u�#Uv�Ȳ=�8�1��"i �%R=����Z$<��;N���@�*=�d9��_ػ9/ =��C=���<`�\=X�<�;����g���Bּպ-=m�<<Z=�����ݛ�i��4=��s=Ro�* =�9)<��<�T�j��<�������Ls<k���C�;1�=�_�b+<DW+<J��ƀ���+ݼ#D����<TT��w.�4�мEe��a�<��_�Y=��S=�Ql���=�E!�R���@b=�A<t�/=f@:~�k=�}�<�d�<T��2P=����C#!=lu�;����݂=�{k�c^u����<��7=j2�c�=�3A=�=*��&#=(��T�,=�溷�
���<�c<YIE<���< D]�>�)=h�,=�/���M�Z�0=��'`K�8&=��<i�i�4�}<�>���	=�NF=���.-8=Z�U������O=zλ<&�w��R?=:o<(�2<�p�����R�<�b�<��B��-=.1�<���;i�=Kq�J�J�(z�;�׼@�=��N�B��<�O�VK+�ҝT��]�;��|��;�=�:�c�k�Xw�<�
2�1���L�B���T�|�ջd1��1d9��z[=�E�o��>�9FJ��s'=�)����}</=�d(�	w��I2�*H�<�b}�]wӼ0�p=�h=,��+���<�=/1=~�=�eϻ���dK <H�K�ȿ��h�%��LQ���<K��l���<#	=�DʼG�4<�K�.�����1 =�`�;��$�ۄp�C�S=6��ts;="|��b;�R=�`=�Z�<�2Ǽ�,ļ����8-��n���cU�dT��"o
��b�<T��8�<�m�<ϑ)���'��=��[=�o9=���c���IK=a���d	=r�Y�.�=]��<�M��ce<�YػC$�<��;�J�u�Q=Ѿ<Н�r%U=ro=���;�#�;�t!���i=�i!����<�Z�+��%�D=�;c�<�iq;2Ӳ�|�:=.�ʼl�o=����<�<�c=�N=�"���˘V=�$��nE=0s[=�j=�=~�X�}p:>���|U=U)=RgX=D���m��;�;�;>�<@�<�!;�c��N�`<�����<��I;�3=�w�;��6��5˼�u+=ĭ���5����;�?;j�>���%=�=5=���<�=;<���&G=i���-v�<֭�<t�Z�$}D�f���%��Fr���<%U���Ul<u�L�̓�<����{˼��<��A=ƽg<����:�b=������K�~EG�@�<�e1�3w[��S�� N���)�4Ǽ�׼&��&ʴ�y*R=�� ��k��N<�<O��<s>�<*��)�t݁�W�����ۼ5���|?�Aq�<W� =~�1=��d=D�"=�	<��J����o��<=Z(�L�7=��<�I�;�EZ:�s=��b������i)=c�^�4S����7<c�3�H�~<:�G=�s/=�46����;�w�\9<<������nr<�4B<�����f�<�83��`�<< �:���;�I�P�$=��I��M6<�<=G<$��j9��A��J=��i�ʲ����_=e���砃�`�6�y4�<��4�7W�;�:�w��ڧ<Nm㼜�ּ��'����>1�؄�PMX=S�C��Y�;1�<�O��g������t=�;��Vb7��t?:��]<-�,=�Z#=I����=�9(�s�h<=K='(���&%�7�<U:��v�;��<9&_a��u=k�8�M�/=@��<����?�<О`<��<�K�i)�'�o�jU�8��I�Zkd��b�<x(���/=�~C��/=�hg=��K�&<2;��e=�=앥�Y�d��#e<JTF=^Ƽc�g=�ἥ{�6(�<����<$�g�<��G:ƨW=��.�R�<~���i�U��0���
��W�<bR$=���
x
<���j,'=2E�<O�<�&�<ͼ��ci¼bl�<�I%�+�O�����]|���T�-�I=ݻ��՗)���a<m�k���X=�)}��j���mR=օN=f�����<zػ<�5�U՜��;��f�<���dʦ���B=��o=�2����G=�@A���n<� ��ܼC�C���<{�h�н߼��9=����]��<�(8=_�;�=���<�뀽���;�=��p=�/�<�A�<�o�28=9A��,λC=|�J=�%=�9&=j�4�Ǔ��8�<9޲<�#='�$=�����I=�c��k���66���伅Պ<<t ��0<l�R=!��էT�BA;����<�l���j�S�;=%:�%D��l:��o=����I���<=�b!��v��o�=���ۼ������t�SG=�y�<*䭼G������<F(�<,-��ٗ�.�h���-�'�v���;��>�<�%�<=�@��"1�B1��<�<?� ��;'�ͼ���=.��R2���p��=,�<wԁ=��,=oV���h=n1�<�hٻŎ/=[ :X�];���<�(T<����#	c��AO<�^=;��hg��~D<�Y
=��R<�ڻ6P���8u���=��M����<rϤ<���Z\6�x�f=��:=D�=��P��I)�8t�����ϼHN����<-��((��0��[�L=��!=%��<=�=B=�8��f$4�u-<-Ƀ��q\=�XM��:�<��3���?Z=W=�qT��;�;���������d�w��<�W(;|=�������<d�E=+=Rw=#����_��Rn�T���GJ<q�=
�;���</0|��]�&44�H��<@�l={<�M(�^ž����<���:Cl <�yy<��ҧ=�/=~���5����=��$=� }��9=�3��;�D�6��<�f_:O�����)�o�e���2=T�6���=���<8�*=�Ē<؄�!+��I���v�Emg��<=�=J =�:�;Vc=� �4-=ˇ�����τ�<^Y/=�����%��wo=�2<k��<�b���"м�z�-�!=�n<�XW<t?n<�pl��J�8�D�9�^���U=����N����+<a@=���<Q�ϻ�<���;A쨻��c�Xt]��j=}R�o��=�r��x=OE��g%��]=T�6=����*6�h����<����� ��@�<��Q=����_=R���O�@=��L=�B�`{{;K�$���O�e(?�����x��D�P=�T=N ��ż��u��VL�Eӗ�;Z������H=�U�~��`E�?��+����<�1��j�QX˻w�<M�2=��p�>l5�%��<(�9�,7<�]m<� n<�/C=R=���XG<\V(=� ��{����s�:ҋe�к�ح��X��
'���Y��{=��Q�Ş<"�����<�T�;�	[���6��Ԋ�p�*=6��tU<�� ;�9=z�s��G=d~����') �(�<���Iۅ<�P<Ó������]=]kJ:�\=�>�̜;�A=ƕ]���H���;h�B<2�k�>�:=�	-;�gt=�
3=s��<��f��N̼\���Ǝ;��	=��=<�|Z=��8��$<81�<K���Hܼ���<�M=�&��#c=�z� ��W�=#ݼ�R�d����4�X	���<��=��Y�<�/��9�I�<S�9�̗A;2�żł��K�&=��ӻ:�}=�� ���MB��h��<��/�}�=8I(���<|��<*����x�<9�"=���;��8=1�'�fn= �=bA-=O�[�T�=GG��S���d�VJB:ň=�����u&�&�_=�	�<��g��Z�I� =6�=q�9�^y7��r�<ټ�4=�l<5%=��=�} ��f$=�ꀽ)wg�m�=� .=��;�S>S=��e=��=8Q=9��<h�<�$��_�{���7K<9ڀ��=p=~c�[�μ��x�U=��hk=���Cn7;Hݴ�3λ�0�� ��/N�s��<��m�����r#����;��_<ԅ˼��5<�e<E���C�<��:�n}�h���.ѻ�x�N�`��f���=^.c=�/��Md=�t[=���G� ��	=.�����Lh�฼�v�#~=�𼶎n=Ls�<����'M��w5;�&���͸}���j��>PO�T�<I&
;�B�_􆼸�F��t������`+��Z�<S�����i4�b�ļjkX�-��<���;�4ż1U�=�й��#=X9�2=�qX��$=(�^=F	W=��c�r�;Q�˼)S"=nyH�e�U��:=<�v=���<Sn�<+�#=�̅<��t=�.�:y��n��:�i�#�`=��Z�˛R�4���'D=vI:��¼�ld=9@�<x?=� ̼n=>X�<�"��O=T��<">���?=�9��NIj;S�_�xŗ��| = �Q=�mb�'�=L�C= 4�<�M�A�.=+k�<���<]�<ZZ�t�D�o��<*T(=��c��y3�v �;�
���T=�D��Ѽ�V�\<ۼ����d� <��c=����+/=����}=P�<�=+����H�N=�s=4`��	��<ȃ&�ͦ���w=�=h�F�2�żH�J=a�u=�.=
�	���<�X��A4��B��<�:���O�;R8���=�ч��2=Zj <�� ��;�;��P=����8�1����H=�h9��9=}@���ۼ�)�<�𦼐�<zY���K�`�/=4I<L�=��ƻo3�H��̚�<�y߼-b;$�=�A�<��k=ޠ�;Ʋ;�+K�<��f=���<q]�����\-�<��H��v��h�;�=��M=Ff�p�$�*چ�Y��<�V=�Գ����;�r=]?�����?����<Id8���o=~M�3� =O3O<�R�<�>U<��=��-=I	 ���H=g�T�Zq �G�8���=�w�g-��@����<�C>��==:	=��$����T�v�r��;Qy=�n�<�����><���#Ȉ�
=X<1�*O7< ��s\6�/��<w�;���<����ޭ<�J4�1|a����<�-��>'��{R�;��S�6��!\��q�u�]��/��g�u����kHg�V��<z6���>���r=Jb1��o�;N<Tg=�[,<�	㻻�����H�!�n��|#� �W=#.��& ��2�.M(<�.?=�=Ur�<s��<�2";\\.��nu=���<��<=.���=���'�<�1=��]=GN�<W��ۄ����M��%=���ª�;�uA�xP=���=ztc=�.a=���Wa�<SD}<S�M="��:=&V=R <�BP=��7�&V<���<�W(;^r�<�
 ��Z���1�:~i=Ym�<��*��;Ѽl�<S
�<�*9=�.���:L��<�1�P�<�ݪ�X=H�4��X�8_�<_3f�q�=	ƻL4=����;f�SJлk�2�������C�S��<�ᐼ��ᅘ<�L=�,��2�d�q�5��)d�aAy�⊽����;�>�<���_�pB�<O>�<V�,������"0<�$g�;�O�[`��4�e���<d�Z�)�1=E��O=Co�5	�r&ѻ��߻��Q<�T���,ȼ%@e�x�E�Z�ټ�a���;��=`ɘ�oj�=�d�<-��;�wB=�;�ۼ�w=��μ���<��ļ�|=���'��C�������B���=�ȉ<�PO=��<��K���/��i_�B��<Ν<����+ڬ���ڻ#�5=F�O�mnD��%=E2���V�;���;D��<,�=9I�=s�5<$r�>q4��d��:^���㼨਼�퓽^e��d�<�[����<�ui��L=]�<ܪW�\[��Y�� v;�H�'����<EdU;��=ɜ><�fJ=+�9=g\���q�PxP�{s[:����[=��<����������l	=�;�଼�R�f����B<������<G���t�;��<Ň:񖸻ʍ<:��<t�<�A#=ļM=�;<����ֲ<+�%��!N<+�u�H#<"�%=�V��W�k��<�\�����3E�K�P�_*<��%=/(!������5=��I<�;����_<�+?=���=����;�s��_� ���ڼZ�#=�Ѽ{�ƻ!��2X���d�#<�L<�����0����=uic�/�
=>��s�;=$K�8 �����Ș<�<ƼU+�<9��부<�I���U�� �#��.�~=s:2;��N=cI��K����<�R=3�2'<i�<g��<]���bH��[=�hC��,=w�Y���<��*��j��G0�i�4;\�<�ʼ��C�cp���=���C��^(<Ҟ�;��\��fd=u��<=Lۼ��T��cS=R���ۋ�@�>�ͦ�<1�ȼs��<�B=X�l=��i='%���w<0�@=��<�/[=�=����o���2�s�4(�;�;<���	�j<�6;�uQ�qOU=�����:��Aɻ��<�:=ak��d�=J�=��?=��Q=8@;�?$���s����<nQ�h���W�a=��ڼ�n<=+�˅��W ��k��Y��7[���;=�JC<׶=we�<0�(<�pP<+"<|pt=B?=��Q;��������ք�s��=�1�<�!��8��88��,=����5�<��*<tQ!<O����<J��<70J=e�:�3�5��Ƽ��<�^I��L�=2����y����<�N�CC�;�m��y��َ<�~��d!J=���<��<i =�+j��,�Aˉ���C��᝼CE<M&��R��\����9W=��e=%���84<�UC����ڼE���T���ς<�c=tQo=���%o:l���5=�*��<�7���˼M;\=WD��⾻H�T=@�B�I�����9�����["<;J_��D<2�E��2b=0&�`��ťR=�s+� �<=���<���<N�<��=g����{�e5�<��� ��nLe���=���<0�9�����I���ڏ;��=ڌ��m�`�l&=L(;3�S=8������i�=��z����=��=��<A�f�����ț��g��踉�7��}J=��<ie3=�^��	 =ܱ���Y�<t=�L����1<��g���<N��;�R����a��=w^�<V�;>
=���<H��<�=a=�ܼ�HB��l��吽-X<=T~:)�<=��<�6�U&�;@�6��,��Xi?�b�����<1=�3R�C�(��tT=B���v���k@<b���k�0���e��S�;T���?��/��<D��:��g���7<�� W�<��0=��{��/�=�{�<�/�y�ż�@,=N`==<����4�A��%��oA����9����<y�Յ�y�<��0<ԎX��v%=���<0����^�<-�;�v6�+s���h�ci��֧<�`#<�4d<e<qO����D�w�=e��)�=0�=�V���L�<�0�� =5@�<��'=�e��v���(�8��1=m��<�}r;l����=�=��b���
��ϵ�w<�<_y#;sI��e�u��<<%�˼2����Ҭ<iUh:����==PX�%ԼF�9�c�h� ���o�8���6���c;xl�;��	���=������!�+;�*U�[7=6����q�<��w*=(,�<�B=��=��H<�,ؼ�K��k*=���[�z���q�Ą��j�<s�r��2��� ׼[�=�*<�)�$�=i�O<ǐ=�^� ����n�:�}c=�NP<��u��x+='���� ;aoq<�����Ւ<]��;�0����T�%�P�<�X����M=���<]���FL�<؈A�#[;q�_=\3]����;�ɼ��<����<ƥ���<F��< ��"�O���#=8������B����<���<E%�5�	P=�����FP���<jY+=�z=�D/=��@=ݝ������׷���ݼ�D��z�<�mX�,���< 8=�]9@����B=]�A<��@��id�-�z���=�Ҁ<@�b�\��2=&pڼ��2=Z[��ن=_;=NP5�χ
�)#=�4M=ǂ=���l�T�=ͭ;ЅԼ = a=hbɼY�+��f�=x�@��-�<9mp��¼;_x<� �<������;�07�d>��	ǯ<�������<��j=5�~=���<9"+<�-��(1�7�"��r����_����C�ʻC`-���p�^�a�/��<eH<�5�Ą���e��CH����ɼ� �<��C��<�m�����k���R�Ǭ���l=��=Ϥ�:�) =7�����G������E��^�W^=������A����o���k�I��Y(=�k=�<�+l���F��m=��ּ�^��t������hX�$���Oё�CA�=�쁽��<e��U0J=jJ;�x0X���3��=B�=h( ���*=�!-=m���"�O=��c;i�N=�u=u�=g�i<C�<G��<P�Z+��#15<ׂ��Wf=1M5=N�;K��T��/6���%;�(�k��g؍<��X��-=�+_���\<��z=��/�iJ<�_D�*����;�<��ȼK�e�tP)�ѧ|���ʹ��i=%�<4?=��<뫈�m/<�N�;��=���<k<E�����;��G�#jмfO�B�<��������<QY��?	��0�n�=�[�~.'��I@��{=��=��)�K�=�
6=W+�;d�<��4<�0
��I���)=:x�'��<m
W=D��7	
=,Ug=}�}=�%����<Z�S����=�oż&u	����3��;d+�<FV��*Ἑ6(���]��:u=�7#�y�7=����[#=��e�(��$\�C>t<{&�<[�P<�z�m�=��E��3:P=�BH��:=�L=D�"<d�M����d�<1qA��$5<e2�Gۺ�0��re��"<�d�92,=�\�֕Z=c�E=ؽ=%�oN�<� �����=�i�����WǑ=�l�
�=�wѩ����<�g��R�(<�BU�1\=���<�s��r�<�g�E)=�+t=���;��g�]��]=��*=������,��q �$�&<����4�m;��+����:���#�l=$~��x��
2��
<�ԻA����^=�,���`�k=��ɻ�{<Q^�hp'=�F��B�:P�5=�<z�=u���i	;x-<=F��N�\�U0�<��B=.L��uz��M4=�5�<�3=���;��֟N=o�,<$�ɼT�6=���G��<�W�]�����1<�Q�;��=c�6=��#�'μ(3=޸�����;C���ua��� � =Y��<~6޼)�B�!=p�R=��;������f=��}�pv<}�'��1���:<OZ=k�b��]*��b<Or��4�A�z�=�Aj��F=DB=�q�;���<�������ʰ�E�;�:6=�����<`�<�Q���3=4ʤ�b'�<��⼔��;Y��<[-�<�EK<1_=V�	<��w�}=%��;ER:�_6=�6�#���5��I�<gЖ��:�_l�l���H:	<)`�� W�w�$���M=��"�_�M��7l�C�<�i=��F59=5;&=��X=/�b�~Ͻ:�X�<�'X=�-�<�V��Ҷz�t��=�*=�C=�A�<U�<\,� ��2z.=g:<!��hf6=�i�����<�#��w@��J�U����i"�<��B=��!<K��<A�@xK=�Ov�_�+=���<<�&�Js%��=!o�;U<�<�?�<M(��+=T_=�����<�F�T,�<Hļ5�X�B�=�ٞ<�<�?��#�v=t�,<T'=$:2�6�I=_�ɺ�(g=y"2��J=�q=.ㄽ^7S=��<��9<�ω<C��o�ƻ�Kv=�ƻ�oP;�!�<��<R�X=Gt�6�R=٧^���"<��/;��=�i=~��ՠ߼������]���*<��Q=Ȑ=0��<f�9�MZ�<q/U=>��<�a����:q�ϻ���<��4��=,���Yv<M趺�R����;%��<a[:={g=8�i�yP��o�O=۷W<�DY=@��;���:�g<�}�Q⳻"�";nٻǎe=���<��=�P�<�B����'��z���>;=��|:���<�=��Z���+=�l�;�=@�<��/=�V�<l%�<������E:kM��1X��IM��=�� =���%��D��|=p" <��,=�5���3�\�����G=���<��<&g�<@PU=��=:Q �VO<���<}�Ҽ��$<�ř<�X�;D� =.�4��p6��ϟ9E%=Ý3=� ���)�<( �<��?�Mݼs�#<�0�j-Լ�Ū:-�;�AM����<��=�i�<O �<Zo(�b2=-�R=)��A@=o=�����}=��u�+y�/�~=�Ł:�ae=a�<�s;����\tQ�)�d��+��)=ɏ'���X���<mJ� Z�<�$J<u<=Y�;�;�x( �L������<PI�r�'=��=-W5���C�[}=�L=�����b=p��1&����<�M��ķϼ{Z�ܑ�<�5ֻ�9�K�<�
,=	�5=y�]�5��<�M��==�u��5�+=�Qc��;�x�<y7�<Ql�<%!�z=��<��F�j8=�_V��׼�d=��;7P};Sug=�c_�����O'=$/C=�5h=5�뻿��v�F=�b1�캝�Ǜ�����<9Ҋ�Y�<W�r,�#��<��D���<F�Ἲ�޼,׫�	M�9C��<����Ӝ�=ɶ2<����w��@�;��=Z���<�](����&����Gc��;,;�����;�p�<�����$�F4B��r뼰�G=
�<�=*=�ZA��
&�^�E��fG<N|�S�=��5�0�U=ޘ��)�pY=�Px���$�e
Z=�	=c*��0��Z_�s=e=�d�ɧ8=�R<b�=���?=�h�pC�菱���]��Z=ş�� ��;�<�켂��	�K<!]�G![<#��<�h6��I�w�<�8�#[�(e=�������<��^=��)��r���
=��K=I�3=Od;�/�9=��<��m=3~|=�z4=����qN=�Q=#�"=kR�Z*=gg�����r����Ԁ��^2�<�]�;�(�,_/=���;�T]��n�-߁��Ą��b+=k�@B=��=B�h�
Q�=ڱ&���Ἓ�=�U�]<������~?�/�]��@v=�=F��tD�=�c��Ϛ���;��\;b��,�����;���-�<�3���;�7 ��N���K=
z_=Q��<�ޣ<�2c��
u��c���Ŗ�  b�ʛ�<݅[9c_Ҽ@�Z��R�<��<B�;h�<a~� 1x��M�Ft�<��n<e>��-А<�J���:�����@T�wQ��5����l=����+=��W�XH�W�%��ۻ�R��D�<@W��"/�C�ڼ|x�π<�/;�"�OI=���%�=l�T=�EW=��n<��:�k�Y��z�`��IE�)o˼E>j���b=�j�j;h{4=�ӡ<	=�,������=��P=
2='M�<�<=��
<n�%X ���=S;W=����Y=B⢼s1\<�HĻ\�(=���[�@�fN��R��<j"����'=|�y<��	<f�-��o<<�r���{���
=�˼l�H<��7�*Q��2���<����}���\'=����7=5���Z%=x�h<<�\�q��-O=0|�������(��@=�Q<:�!=�%Ӽ�u�<��;n�<��ӓ�-�缠_j�G�=�1=2 l��TB=� 0��yJ<r��3M��w��!�<vui=Ԟf��jf�	K����;����'k<x�;6�2=~�';�K.=��
�|�@��<��N=��K=���(=�{P<K�=`'�M���P��N:=�O ��c���-_�@�%��� �����p=��:�����8=�]����;�[�:�:5=��J=֦�<���<G�=(�)�����I�2=h�Y=���wp=�#=��V<���=O1<���<8��u�i�ٝ ���:��H������m=ޢn�j���Q���<k�ü#1j��=Ab��c�\Nt�ڏ���)=\c=��ݼ:J^=�8�dzk�Jo=4LT�I5�2�<6�=����<�`=�/�jnB=��P="D%=YY�ɩ@=����<	�^��k7��M��ͺ{:��A=�R�����h=C���D=�}X=o�:=�';y���������e������u<I�Q���o��~P=�����~��P�]2���_n����;�k�F�����=ʅ<,� �o5�S�<���*1�%������e绅��:e1�:�:=n�\�E��<�=�Q����T��<K���1��O��W�Ĭ�fM<��<:�"E���<{f<�X�����<>k��n���7�<q�����v���V�p��[ǣ<�KY�2��<hP=�Xl�3t<<,A�<��Pk�<\B-=#˙�w!B���5=���y�#=��J;�^j=Lx=�,d�`�a�="=���<S�G��ka<�l���੼���<M�&�Q^O= �=nRP=lZ�<��ٻ8,K<�2�G7=�)=�6`�<�[^�B�i��p�
�;��9K���OƼtL�<��<ԟe=p���Q=�t<Ú�;��=� ���a�ѨO��Ӊ:$:ټrj:� \�z��5 8�v�<�#�<�zļd{f<��~=���OĎ<$����N<:��<�Z^=;�w��C��8�W<a��,e=O�v���<b
��x��«<��<w>=MQ<4�9���<�2ؼ�M�18=�)�<��F=��h�����Ψ=<��8PL�f�j�f�-<_�<�?rB=�g=�B7���6:N�Kk�<<�F����SК<�wﻘP':pA�<��<l]��p>=,-?�pޙ�
!�;���=�Re�FrK=�c�;�f=��v��[=�Lϼ�6��S()=���������)�<	X༣$!�c~���i��h[�;�<����<�=.�l=W���5�����^=vW=�䎼C2;��<7���k=P�Y���\nN=<nJ�?�����i��񒼆��z�=u��ݷ�<ŧ��>�h=�������V� ��!��Ys���u��;J�%��<e�;v-E�x`ۻ��滈�N;�=dj=����=������}=r���X��x=x����m���6�>4W�7�B<:�<�j�;���I6=�K���;�.5=��V=�_�<���q��<
L�<?�v���#��}-=�jĻ��b��;�U��x�<G�b��_J<I�N<@<�C�\^ ��?���?�T��;_-��Ķ�<�vX���d���<�lC=��B��M�<��ѻ�[�i�ȼ�$:�'��<P�=~
;�7=-e</P�<���;D��<�=pK�1�6=�L�<Fl��Q=*C�ױ��ÿ	�N�-=�ë��6꼇��<��R���<��,���<�??=z��6_�<�;�<0�_�D��5���K�*�H�<@rڼe.i<�bG<v*ݼ:aj�D�r;J�s=Ѱ���2<毑<���<��=KbԼB�=Ù��<�A��,!�%$;odl�U�D;=��<����d7��$�
�<���<o��+��r�9hJ=yμ�&=s��<O�=��=�6=s�-=���<����_<��N���<~�v=���<H��<��I=�{=X��ؓ;����w�? ��Q�)��=��#��<m�<�x��v�;VHd����6��<��=��L<�ET<'���v=�U�5�w��I*�P:꼝g��^C�<������!�]�2���<*�����<��<"�<<z�S=6��;wg���B=��H=t�<R	�<�܋=|����>��5�-�H�F�����0=��5<.�i<��O=\���3q=��/<�x�<_��<�<�?�q�R:G�e=,I=^U�;��&�ü��˼�"�RH��2�H=HӼ��<����lK:��]<������<�.���&=�	��M=�����H���;vm�n�9<!�<;��P����a��
�<��ܼP:=+�<�[�w�<�A�<L��:�=<�̻X͗�[�=ĢF=(=�M���x�9�9/)0=9#�<�0T�U�D=�=����t�<����c4=@�3<��`=�=���;S��<\ql�� ���:=pK=�ޜ<��ܻ(B��~t=���<Gu=@� ���H=2�N=Y=��%���I�=�e��px�?�<�s+���=���:��R�\=���T�=��pB=���;;Ӽ�d������K=�tx;/ޙ<�,��u|=0�|<�_��'=,�N<�( �~�4����<�Bs��͒�7'=�%���k=��=�2����F�r�=�V��:=0�\=��g=,G�Ĝ<Y��z��>�*�f�(�06��b�p��<��o=J7�<M�.='��%뼫U<='��� 	�wr�)xd�J@=Q�f<�iR���Ҽ���:�\��.Z/��QҼ�:=X]���R��<	鋼��<���:ռ�t�:�
=�Us�2*=�,�sx�<q���-=��5�Nن;��<N�i<�Xڼ5�;�~�xb�<�+�G��C�/�A\>=Iw�<O�W=iV��9<�1)=����$Ĩ�H��B��<��=�=�+3��?Y=s7><�ɡ<�=���<p|�:�]�VM>=z`E=�Z�<�4���X=Β�<��<-x�;p�.��F;Sr�;n�L��'a��ټ�Z=�%�v�<�_y=1�Q�bc���_����fL=�?�:��[�m`#����]ީ�5��<����?��-�;"�r=xI��R=K�P<\ñ�K+��#꼸x|;mh^����<��<�ĜZ�8�=T���|��ɛ�;��=�q<�����=:��M�%=�߼�W�;�<�<O�#=2�8��={%�<�|�<a��<�z�n�<-�J=+��<`07=w��<��H	<��%=3�?��ǋ�o�����H=K��<��<kc�V;=�M=	�L��;%>��Ү;�#;�u���c����'XG=ק�c�5����<�mS�&�N=�s(=� ��<n�<�?8=����|<,lk=�=�A(=��S=zK:N=u®<k�n<�A¼�o����6�����4=�P�+�+�����h�;��=!;=��=C+��Wm�V�y�/���W0�ҹּuIռ10<��=�{<��T�����<����ƽ<t���,�ܻΖ=��w�漏�P=�+��[��n:<AR=�&����'��$ ={����<_6 =�+�<�Vu=�m�<��:��)'�i��C�)���"���Z=?z߼a-��f��<I��R��<;<����}�A:���������YZ=�7O<���;Î-<L�=|S=�t�p,
�"������޾�з@� ߪ;�<=�-�Aɧ�5�=W�X<5%B�)jm���ܼc��<D���, T=m&=�a��}�<If��Nd<��<$tg��z��<8-���V;O������j�<���<�l=�,��%�<$�T�_�B�}\�<�[=}�a=��(<So�;4
c=rM!��쿼�{;����<��<����gf�Z=�M�<9u�<��ݻ"�&�U=�3=���<f,˼5�L=F��<�9M=J�?�$h2=��4���m��-�=o��<�J����k�9=�f+=�h7�	g=#]ʺ��#���=H�q���	=��O=P�<;u3=��_=QbQ���o<C�<�<?���$Z�5�=9)=�Z�<��"=�y�<U搼=6I�}U�;������A�	r��&��,��<�T�<�4�����h)��j�^�Ai;�	X�T1=n�^=/9����<'E?���i�i�$9�<Y8=�QY<������.(~�;r�r&9=�2�۠g=[�/����<��9<r���%c,�,z�y?`���Ǽ.�7�-=��R=��?=����@w-=w75�A5���<N�B�@���Gf=P�4������R=*�u�1U.=i��<����)��[�(w�B�e=�}�<쀣<4*=@�ĺPЩ;���<Tճ<�y��1�����X»�O=�?=9�8�r��=��7=̼ބ<�q= �[�[���<U�<�G����*=֤����1=��4����=�+=VV�}z�:������P�P����<�|�R<�8:;���<�C���<�ʦ<M�=�<��<w�U=C*='�S�eP�h�Q<2���^0�;K�����]�<M�I=�L��dD���hd��#�<^�<q�ۼY$n=Le-=�Ơ���ϼ��<[����pV=��A�_4���2<��)��^
<]�ڼ�E��ʜ�Y �`�7��.<�1�<�d�<�k��Z8p<Ϸi=��=_�<mdo���0�Z�8=y"=�7H<�%x<�zr=��	����d=�8�;�J=_�t�'L����<�^=��i<�)?<�0s=�A��W�D�뼇fk=Ll�;��/���+��߃;dd��5�ռ�V=�?)=V謁���|:�9´���x=�r�<�^U�>:_=�;�;�v@=&.��M��Oa�<��q��Ɍ<�zo=��C���R�'^%���;ri��\���<ᙹ;�켶rt�8º��s��1�<":��#=�v�<7*�5����<��)=6�=���y�=���<��O=�,���O��Go��1�<���bFR=��R�[�$���ϼ��L�E�?�"ȼ���	��4a����<��T�<;=�ܖ=wֻ��=%7.=�	�;���<r!�<wƼ�I�TZ��-�h=>�G=�^=Lл���<C��'���`=��i�=R8=�-G<���=��j<嶡��PC��6�L�<�����v���<=G���}�*=A�Ǽ�g��2��]�<�L�<|��=���E��P�0]I��F=��=��K��Ӎi�5�=�/)���<�e:=}F�<jbM���<wn�<;�����h�<�I=�ݩ<�&/�+�<s:D��J`��;�:@=�	a����<?M=rP;�v�<Ÿ�3Ⱥ_���c�;����b��+!(=��=�(;/6<	l�;h����G;�^z��V�Ev=<�.�B�P#0<�ɼ�\���WI�i8Z;�h=��w�y{e�}�-��<I�D�d�<>(����*:u<�ၼ�I��z�Ѽ�'�<�"?��J<�W�3ga���f=�g�<���Qc�<#i�<[	�<E�Q;㙧���<L�Y��}��} ��):�=�A�X;'1���Q�Y=����%�2�u���
=�UC=�T�a!=�CV�Da��S+=`�m=j��<p!1<Of�\�=,�"=h�|�*ů<�������xs=5޻�o�<-�<�Z�<-��<�=<]���,=�&q<�D@��L<+�f�(�s�xVF<l���D S�8����<�E�6+�<���2�<�<�<Xk.�jkμo}z��L=r.��>�<�K��� ]�I�^=��B<?}J=LaM=�=޼f��<�%¼~��<���<k�=!	h���.�G
���>,��V�{EQ=KZ=6�μP;�?��0W�{�==�ؼ$����$���<Xc=�=sla��2�/�2=�0=�Ԩ�N=�ʼ�M��m:�;�g�:d�<a:�=�Rn���d=�n=�u#����<�Zg��E�<z ;�J=�f�<��;�T�iz=.0<�>oC=����_��s7^���9�&��<��<��=�+�<:D�6�<���<<��;pԺ���Du�;!�:��R��z�;���<}-=�h��A.��}�1Z<1}=�&i��h\=���N�=D��;\\=���<��;�XI<�eI=��E=:;4<��S-��WN�c0=WP��;<o�.;<�R(�<��t<q��^�7=&;C,5��y9�
	�<�"ټ�=�rJ����<�e<�0=�j���ӫ�a�<�K�=إ�<gr�ihX=�"ɺu�v=��,lM=���:�u�<��>=���ǌT=��C�q��<�g�^F;ո<�]�qC���L='��>��;A�-��x<��=��d�f�m���w;�U����ѻe#+<os��#~��p��	�a�j�=�ζ<~	�q�N=��]�Ř'=d2h�U���O4����a�ܼJ��<}�$���W=�/L�%�n< ��#N=�A:���<I�A���!=Z�d<�;<�7м��_=!�x�
�<Cq?=F/<�b?�F����;;3����=�G=xМ���6���=�|&="lL��^��$��:��<hբ<���;�x;d��<������<0xc�-�=��6?Z=E
��@���=4=��<D�=�[6��=���<��g�X}��R�=#�=H'�C͸��W:=Jn�-$X���|<�����c�\��m�^=�<�Z�<&��0�E�X�ۼ��`<Ni =�s��z&=w@�x�<�f�R=q���Ͱ<�Ie<�.6;ʣ�����<
WX;�0���8=��<�7���<��߼�E"=�U�@�=
<o�꼺v�<qa=�8��n����;B�8�89 ��7s�=Ƅ��j=�����j=o�����w��LI=�+�<�k�<C�;H/�;�ϻ�n$=���<��;�
S=�=y=,����(?�b�i=���<��<�b<|�<K��;��$<Ǘ�L�|<UY=2�6=wTD=�으8�s�r�:=
�=+��<3�1�m	�:���ؿ�95f�z�l��G�la�<�p�<�'����=0ˆ=0ui��,O�pR��(Q8�wC=������e�;B�P�7�@=�K=8Qe� �=U��<��x�١�;�^���=L�.=m2��S<�t��<�CI=ޞ�<3B�=�C=����y�<�.'=?�_=Փ�|�:��w��=�Pd�}ƍ<��<��ʼx�7=E�(�2�<Z�>�Ģ���`μY����i=��q��=�����o��R=y�a�݂�����M=2��p�F=����;F;�^h�7��� ="�;=k�#��V�;��-�i�N<��=�=�B�;�;�>`�gZ�<�v��ς���7=ͼ;��s����^��C=P%<M��:`��������I$��u+F=|�~=�N̼�<DD7=3�&=��5=��j=M���B�,�s�=��=��X=��;�<���ǝ$�4�����<Ϙ=�\4�V���6%�� ;����g);�#���N��#�<����*�;�7F<���VL��`�*O�<� �= c˼;�;=��;��<b���AP�=�=(�:��F<[8^��4=v#w�N�V=��ȼ>]�<�9�n4=(�4�w��<|�=�G2=��=|LM=�2F=�6޻��'�"�^��=C�G�6�Y=�m�Y�S�aT���<��@=�V0=�6�<tyN�V[�<��Y��Ξ��\Q�&�F<.=��ȼR�<�/�������<�Լ܈<��bL�X�Q�����<�L�<�o =�{=8׻cf2=@u��q�>=�{V=%�;=�f��ܴ���y=t7��|���6���·�eG`�fq9�]e=oqX=��l�-�r��eͼT���q=�8f<+_������	=h�j=q�=��k;x.=��l=�������=7ԅ�ZCI�窼9D���u6<ЙE��>&=	N�\>�<���;`N�.��<*OA����g|��l=^�;����;��q��Y=�y/=g&f��b6���9��{z�~��r=M���.$=��;�YC�xK�8���}�<�w����-��ϼ�:,�ʸ]=�������(&=�\��;�;���&��<�<Ł*;�x"<*�|��<l�1=����b�}=�8�筻���<m�=�$2=d2=P��� t�:�%=��I���=z()=2�j=f�;<�vۼ���<O��<��;�e=41=�!�:څ���:&�Q�jrb��gM�'=�?d��L�]�����"��}�<�`=��=� =��=���<�V=�<;��� =aП<[��<����9��=U����B<&)�<�-=��ʼ�^�$$����*�P�,�T����,=�Ҽ`��7�=R�_<�-��u�<�_=�m�J/2=!G����I��`�<�j���g<�C����<��켊Һ��~���ؼ�E=�2j=u�;<	�G��m;�\�=`;0�}4�-��;Q�2��P�������SV=R���`4�BTK��(=k��<��
��<�=�h9�~My�*�[=�/=�_3=��;ֈ��'��q^���=؉ =����SZE=�L�:���"�}��M�
V�<�5O<X�<8{]��[�7�<k���K=��z=�_<�4��k�^<�$����;|CQ�����8��a-=?�=(=��=n�/��"����=���<�-�[�5�L��\L�<���R�=���=�b;/�9�%L<Sgj���.�"�<�+�+�8�^+��b��<ZwC�n���k�=I�м}���5�ͻ�SP�a2�� _��l�<}=QQ+��X)=gD�=m���/��1�=LX�<<�ժ<�Ǚ���K=��^�Z%,=�A�(�����~~�(����8=Y쉼u�ҼY =d��<z�<��<K%���<G�<��n�s0=��M=�,�<@�)����;�O_�	ۻM
4�.7���끽	�����M<�,���N�Tx�����<t=D���c<c������=�[�R3|<6�L��=�_5<{ ߼�3F�RJ}�뤺��MD�J?���ˏ���)=�y�</�̼�պ.H"����;ME�'-����<�:=F���Y����<#�M�}��9�h�=�`�C�^\0<�R������~&�g ����+�>=�FH=p|�;��0�3X=�YT���0��=g=]�%;�ZP�����K
=�r�<����v�~nu�9xS<W�p��si��0���ͻl��<V^ =���<8˽���@�f$J�|�D=jD=,=�=ky�h!�<�8=��i<��t=�)k�RA:=���<���;�I���,�C�Y=�:ȓ�k��b���	�ؼI: �(|X� 0<u�i�SWF</��]d�!�g�)�8=O
=�r�;��$=j���h�F*�=����C	��ϼ���<�(#�%,�<Z�+=�4�x��$�<�@=B�c<+弘�<�Q0���&�Z�3����<��:����'EɼNV�~Z7�F��<Ecż0N=-� =���<4�L==�¼i����.=�U=�؇���<�n*�O�~hv<�?P��R<qS<9�7���c��C����y� 
=w�^=~;i<��s���n=l琼��<��v9y�����S���-=��3�LǼ�}P�OۼOļ8��q=*G=��1��:�9h�s��I�&�)ﻼ\��G=�@�<L�=P&��/[=0�=ܯC<O���ZT=R�<��p=2��-Z�<`��w]=�^Q����;���;��༫2T�jr~<�߻�W�<���`Q=ydS<K�~���O=�)��P	�;?��;�<ûϴE=��ջu�~�YqI:>�S�6�g=I�=*��:���<��<�80<d4	��@��y���l���;xG=-^�<��C=���HOE==:�ճ(=�.�<��<fx�<^�I<֨^�͓!=���<}"�=d�4=�N6���=��;��������O=b��<>�Z;����������n0�͈2=S#ݼ2�����9��"O>=��+=)!<X�p��Y�0�6�).Z�Y��<�q<i�-��I<��=Z�J�hPk���Լ�).=S�<����R��!	�!֪��J==��:�kQ�Ĩ��砼#��N,=.�W�P�j��=+�=��@����<�*=�~j�HO��,�5u2=�]1�:ö��������T:�=o���9=�0��Փ<����BA��?=�&���=)�<�&=���<B!%=M&6=@�0�3F=���<'-d�z_$=��=���<"=g�����8=I=X&=L���1�<��j=.` �5=��O=~��>��<t����6�<�o;e�O���&=�B=ڟ��Wn���!�M7%=p�v��)=�=�6�<wn����<+ͯ�A=+�#=��D�=O=UY�<��W�+��Qb;�(`=�7��������:��zG=��I��c<w=�
m�58�<.��<7�X=���<�ʜ<�+=Ac&=�Iw�������:�����<#L�<6��<G��<�N���M�Ҽl� � �=҅���-=�<QsI�1 =�k��FE=b.V�w�u;Wt��7����%=��s=ݗr<���<�w
={�=b��SM�����<0�T<<�;=:�<�F���VK<��^<�sk�t<SIy<kI?=�@�<�IмYBJ�1%��5̼��&=	=��:�W��<-�e<�[�����9�<z:<�}�<�ɼ�����?��eNg�r<� P���=��S���.�7�=���<-D���^ּtB=�J��mh��
��3�<4�<	 c;53#<�(1�>A=y��9���<r�cI=��M��Բ;$9t�k�/<���:7Jv9ޙ)�3+�)���6cq<V��k�=��8�Iq�O[?=:,=��;Q�w=db����<��T=�� ���#=B�k=��������C�j-2�'>޼�{Y<��=^�|�L��<�I�<����)M���<Fς=x�j<�n=EJ���=����� ?<o�B=���؏=�9<N;!<��<DÌ��#���oH=�$V=����=[2�)�
�����(���k��؍�R��:��=��¼ᨿ�-vX<���<I��<��༂&����T<uF5=ٜ�<�N�<O��<;c��3-��ߌ�M\���u<�ǲ<�d=�/���F<V0C=��1=��;��ϻ}Vz;�uݺA�b=|�f���<���=�2=}P#<P}�<.*M����<]u���M=)@<$/<��3�KI*=��<�<��ح�C᰼�b��P��_���aL�p̀=�4<'%�և#=�%=���.=J��<E�λcR�< �1�����u�ۼȁ��Ó��c��u�¼+6�<ؑ-�W�<}~�<3�0<�&%=��,��SԼ����o=�bļs1���X|<7���󼘰��_�<)U	���P<i�V=/�\�3#c�U�.��"=�>m=�[m=�����7�f��y��<j]K�&B1��{B=��]�#���n����<��_��o�<��(=dW=O�ƺ�\�%�<��=W N=6,B=�#=��=]�˼��%=����[�<�-=�[v=_����	�w�ܺ?�=��|=�cf�?J���A���;M��ꌻ3?��e��q^M<�D<	��<�S����g�5�ͼt`�<��A=~���ӟ���<�e=%y/�Ŋ^���so_�z��=�1��4b<�<v=�B=����ŗ��Js�I(Z;�<B��<�xJ�銏�uR�����dW�;�����1��Q��I��5\��c,=uW=�w��l��q��<9�K=H��<���;|0��
�<ҏ;��i=�	��U�=&G�<��-=�-�u0'�G���R=$=�ƼX"���� =af<=��Ѽ�_�ƍ�<��a=��>=A����<=ۈ<OCy�KH=v�(�����b=��P�҉��'�\=�/����I�H��:B.Ҽu�K=E ��V���@/����:������A=ߌ�:`5K�}�05=K����;B�0=�L<��<HdU�ߗ�<���p4����r=�!�<Y�l=}���K<W5�<5b=7==�{Z���<:ۅ;���<ͱ|��EI=�5����̼n�=�U���}=��W<��<��|<��_;���<ϸ��'��:�s<R=J$�<�)�;h�<}�����<�~�<��X����;�����C���/=� =򏰼��U;���nP=�� =?�<w}U=�H=��<ܑX�Y$�<��c��4 ��թ�s�.�nހ���$=sA�[[;��k?=��;���������9�%=~ʊ�v�<ܸV���<��<ռ�<��ݼyP�����Rj���:N4J=.��L�M=]vټY-=�e�mn3����<۪����=Q�<�ݶ���<�ل��%=�
�<�RM=�.����=:�<D�;,s�B-=lU3����<���<�����ӉP<�U:��>1<�u����:�,�;�$�XE<E�:<\;=-��?�G=�:<X��=�t�=)d���˼��<&i�����<̡�<UT=Ug<�o�9!��0��<�T��<�t<��@�^,��O�=��<=��<T�T/�T	L="��;S<k�ܻIs��ۿ�@�^=Le^���V��Nƻ��<�M%���tr;=:-�<s�=���㼀�a=�>�<�r���B�C}y=���<��H=-(�;q�==^DP�{�἞�0:����0<��4=q���	���
m=VaL=��<=>LN�3��<S�=?X<��f=�^A��(�7V����=��2�>�<�7=�$�<�Q:�:ƻ� =M�j<��~=��f<U��<OAL=Yz�����/��<�O#=�/=[U�6M=���<��Ȳ<o���Ӎ�$��<��E��t�@�W��=~Bw��X��o3=�W-=����l+=�b���F&=X�ۼ=�A=ɬ�=��<B�:p�9��@=�5!��Ԡ���s=��"�����I�;��"=en��^=���J<<��N�#��<��<�C�����+�[C<}I�<�=��=>�������]���g�һG6���<�o��}٫<{t=�
f�2�<Iwo�j==�T��^]=q�f=��弽�0=aX�;>�z�~�<tC����;� !�Ȱ)=��g=��*=�ڼ`�Fh�<2��<VH�;���<~���v�<�'ɼLvx=m,�6�)��	���N�!�tN�� �<���B\�<���<��x=CѼh��<|�_�u�r�T�N-=��μc���'e&�9s?�̝(=[A��M<��r�к� qf;�z=���=�t��;���;�+���d����y=cb=Qݓ;F�ѡD=Z���q�<�3�=~��;zk�U�O=k-=~=�#=���<�hH=6K�N���=��.,���<�+z<F&=Bʖ:0���G㽼���y��<��c���K�lE|<�L�;<�I��N�Pc=Uo=IѼ-]�<���<j��<PU=#��<,+����U=�\�<���fh�8$\=�����C�՗A�[`�&e=)+=���;D �<�v<��]=��h_A���W<e�m=����kt�}�S=E��;��>��"=;�式t<��'}"=ի�;�r
���O��;��؂�3�)=�r"=C���y�=g	?=�r�<q	C��[8=�X�����&L��}2Z=���&����iQ��n��@���nR�;���A#5<�
�=�-)�� �f��"���eA��v8=���<J�!=?�'=#�B:ł^<o�=o_��;4ͼ%�7�N.=�gC�2�N�����;�<�s�����֟�Dh�^� =��=�OV<���;!=�9<�kI=	 =7ü�� �G|T=��0�eI=ᔰ�f`O=s��<@QD<�g<l��<C=�V�;�<'��I�<�yL�_�=�
��[�� E=��]<�9;� g=�>=ZU=�gF��8T��<*�<�9��4���z�Bf���,��%<�:Y<��=~b=�&��t=H�O=��+/P�k�=���<S|���<U��<�3\=ne���~������H=�����^C�oFJ�P�$����Ί?=�=�����6]����1cl=Q���<w�=��!��ܩ<8D��0�;y�;G�<���y���|�<-oT��Y���ټ5+;��M8��=��"=\`�<�=3=ۙ7��L�<��U=z]�:EWS=�<�K;-�D:}f��z(�#��<�h���cM=��ּ��~=��D�CZ�<�����l� �=�=[,��m�=25ü94�;+���'	=�d�po�;-v=��<�'=��P<Cm5�b�Z=�#���%=5�T<χ��
���!�<{�I��=Y1������^/�=9�9c��z���/��D�=��<+��:�ی<��1���e:[m]��#=9!�������>=��<����VG���Q=���R�%�.�=T�M�ǉ#=�n�����<J�2���(�}��Ɗ=<��;��z������'���Z<.s'=��,��)=پ��G9�:I=*�q<�i����ȁ��Q<�u�<~�0��_��WX����:�5<�BE=��1=�5N�I ���T�<<�=��*=>�M�����,=���<��*=�4��n=;�I=*����s;�{E�(�N<���<u�?@�=_r��	^<%Q�
A�<�=	<���<�#.�"e=I�T<t.��/����Q��#��S�^����<:7��7�X<Z�C��MV=�=�͹�
�<�=�=��u�<�P���.���;��-	��ɼ��=�=�╽�+d<s�b=�ܺ��<��E:�;9��<~ f�%�c�٨@=�<�w=��=%�p���<W��i�<5L<�&�<+$�<�q��`ߥ�%N2<B��<�Ή���q�-�57=�%=g���Ё�14=��<p�\���<���<�pF��_j=�I��5�m= �<}mu<�jB�$��<8>-��"6=N�d��-�<�n=� =���;�=���<e�"=Pk�;L�9<����?������8bW=b�������&z>� �x�]RK����q.����Rpz=��V�݋�F�V=y�n=�#m��S<=�q��j����i=L�!=�1�u��<��N<�=
C<25X���<��<�[=�tp=�IB��@��[/=zOU���=g�0�@<l4���;�5=�(��&=�Pr����;�Q=�A=�@A=o���
`^�ݠ_<GL���==;:�B���=�-�n���[Eݺ#��<ڏ�<�0���<�i=�jn��[��%�<J��<���<]^�;)�<.�q=�E�;xT>�]�<z<�<!��7(�<����>=���<`��=�=�<��9��l��Z�=�$"=�u�<��V�N�<��[��|R=�}��v�<�^�<�h�<���<ƩO�^r缄hF���$���B=j����ͼ������;�#0=�=!=���<��;�K�Q�X��D��J!�H�J���3��ؙ��	*;Yn���[=4VA�@G�:_p���n�<C����M�Ǣ�8D8����<8�y��������щ<��$<�@�K�7�Ꝛ��:=��<<�m7��)W��1ؼ�O�<��;#�K�EI=_��h�`��(�Q��<��-=���W�L=��O<��=�<8�nL����Z�8_�E��5���<���+���b�<�Fl=�K���!��w	=IBݻ�����`��������[j`����Q�~<�&�<[:�:|%�0�����=���3���~���@=�p�bL<QH�<�-H=�<�ו<�J8��%=l�x=}�=x�;B�0=<cl<�{�<���M?K��s��-@=q��s��<M���^b =u���=��_a=��j=��;��h=��[='|�<ak6<)�T=�<��� =�D=�P��{m:��'K�O�z<��/=�J=�:Y���_<���<]���'{=� �<g�:1z��B����a<æ���=9FV=��I�('<���W��<K�:���'*�<!�I�Pu�Xkn��=�uM<R�b��ip<�G=�[���<ǳ�;)�;=t�¼~���'��A�)=�]�k���	3��u�=>��<�E�F��b�Ǽ��S<��\<{��<h=i���+�O����<m��<o�+���=<x1k�g�;�i(<�B=ΛN��_=$�&<�ϥ<Y(�o8�,>N=i��<-�O� �W=+b�<��<�k�+�\�%cF�9^-�j	<_ ==OhE��4���e;:Ot=���%�g�:E?�E�˼�������<���<�eB�M�k�ˍ1=��M�`;Y=�桼]�-�D=�3��df=�p��xH���y��n<%V=�Ez�7Y=�+7��X=��=/�_`ͼ��!�7�o��k	=�E�ow==B���\�=3I=�I2�T��</�2���
���P="ߺ�JE=��w<i)�=t֗<���<�l'���J��!:�W�<E�$����<����C<X�<�<E�~�<�<=�C�\�,=p���\<S=�N<�d\�5T=~�=r��<}��e.�Ń�<�G���h=��z=`���%�M�Sf"�v�;(���	D��4�=,.ټ�$3���C�����)�D<f��<�v׼��?���z�k��-��<(8<�k�:r�8�C.�<Öڼ�{:j��;B=c6#�r�q��W��w!�;�<�V(�ni;u�:	��N!�<���;����2˻W{�<�S_=�d;�B��϶;/|��i�i=z������B�<u��<rUk�2�H����ڼ�#üv���f�b<��*���<�2@<��������P�<�*ĺ���w�0���o<6݄��2���g�X~B<��g<ٻ�<�f=�7��C9��<����I*��71��`���¶<E=��<
ʻ�1���=k�=�W=�y��%=�h\���=�@�<?�U���F��i%=�=����J���1=��=�`��F�<`��:��=�=U�/���$�I�<�=s;��$8,=�%�<K�g=���<��� �K=Un�6O<���D�;�<a����<��i=�_�<�>=h{�<[Y3��-?:�S�m���Hs��Ĕ��6�<,�<�"�<S�g�H����F���� ;�$��sY==�B=/���q�<��=�=�V=���:��t�Le��n=�q ?�m�-���R=��<�w<pL"���X=a>w�W�f�[YA;�ؑ�^xE=�&�<�3'=�I<V/X��t�<lYN=�U<_׼�ɼ��E=����Ў���<�N�<�<w=�.=�g<�������<���<f�'�
�Ӽ
f=X�?=����c01<;K"<TJ�<��=��������$>=�'<2���+�=S.V<T�=�x�>��9@����d=!���V=[#-=^-}��/�P��<��=����<VE^=�J���s��(�<7n�<�6:*n��ݒ;�=�f=��-=�e�<uu�<5D=����Ҽ�b=��U0���Q�4�;�;�V������<[ׅ�/�<|^ټyּr�-=d�<��K����<W@;s�&�@�l)ļ�x|���߼FdK�O�߼�h��>�d=y|�<%<�N�X�L=\�@��L<�[=��L<��^��c���'*=!SO�P�;kq;߯\=��ͼ�P&��pJ=s�3=y�[��׵<=�R�/=}�S=�l=�%�\�r<�ol�"�d�\�"�.м-m��_�U=k��<�꛼�7<��Ȃ;��6=��H<s�w�*=w(����H���|��Ļ��#��QV=F5Ҽ�.�D\�<bp�<˯*<�Uϼ2��L���JR��C��߈<^��<��<�V=�񈽏!<�7�������;}��5m��R�$��=��)��<"�!�Գ<�5<�鿰��c.�.�'=��.=j��<I���=xv<!2�<��P���<�_����;��:Դ?��C<Oü��1c>=S��<L٭<4�=h�z��<v�5<��;�����u<��2�8I��+����O��<��<fo-=�[h=�L;���::!��_eY�!C'=���h�J;�zm<SL�Ә����d9��`��u�9�g�;�)��V=�%=���4��<��_=��˼�@X=�d]��`��aϠ;��2<6?=�x����ϻhM�����;Cɵ�P*=v(��=���
<�8n�ζC=�~=�$�>F_=`����V宻�y��ln�@��9-� \=P=n�>=7#=�m��H��ы=�z���=Wh�<��=R��jn=��g���� °�t=U�1�K=�z��L
=@�<��w��JZ<A}�<�}==��켮u��譼 ���+9�C�,<2�<�<�)�^�޻2�4=M$��0�<��5=H$a��v�����<n�A=��n���=�2�8$-���J�G*T�<�>=��ռ�� ���F�U�E�<�����=J �<��:��=Վ�;��"=c�\�=��\=��8=�'�[��kɼv�zǼH=n/�80=�Ba<r�=���<�,�;�F�U<� ��} <�^�<�R!���\=�L+�D� <�]i�ھ<��ܼLC༬rG;������?=E^���:�0�<��<�/�<0��=`|=�v<m/�ZJ=u��<�3D��?!�V;ȫ���M=%��<&s=��5�D���ʻ7%�<↼@�]=��;�$,=�m=�;^�a�5=b�(�A�=�2�а�<
<,�-�������<��,��@�<q,��K��Ȼ1�b��<���<=-�=����/0=�9�;3���Y�<X�<2r�� ߼��&����	�;S�<3��<[�,��%�;������`������3<�$m'�uoN�=����=-���l�:��(<`F�;��8G�U�м+VM=�Q<��<O¼n;'��s=Ɵc=/R�`�<�AG���%"1���[=]�<�}�	�y�7�<��ۼ�ǧ<{M¼[�J;�b���b�vyݼֵ��|S=�
;�[��)=�4�<�ɼ8��e�&=�;�+J=�S���w��
<<�5�Y�����<L�=�@<#Qx;Q�5�����<[����×<kV'�B�,��o4�l� =���<��<={����O=Qj�9_N=��i=�
=H t<�2=6l����<Q�}=� =�L��=;�}-�r-�< �l�-�=�=���;�ӂ<0/�<0s�^b��,��d=�`м��I�i����<X��˒ ���(���m=��ü/O-:}�3�^�.=ߘ:�Қ��FT�XNa��u��e�<�gG�U�����<Q�6�m(o������58=�U�W�;/�;j3a�|��vz�<��
=8b=+�=��:�o���5k��IԼ�x���h�`�=1=M�"=�ϼ�6=��*<&S|�K+S��׻����3＆�D9����oL��I�\�B=Wi�=+'e����T'� ��<[�!�W�j<x���R`����?�G8���ټ���*��dUL���l<�Z���+׻R�W=c�@�'�'=��<�?S�z;�l|&;�]G��˟�>v�<�5�<�PL�|Y=��H�?l;�m���<&*ݺ��N;CY�<�V+��T0<�:=��J�(=�4=-�P�_��<�,��A�v�aW����<񪐼V�J��x���u�[�ܼ �+���<g���yv@=�T�jŻ����|�ؼ#ȓ���W<���<�2=�<�$�<�;��3=�J���9�v�Q=��9��F��է�׻���T�m�=�6�<�eJ=��<�ż)��<Rȼ[D����<��<��;��M�y�$:)�c�*4B�<.j<�ol�[�jP&=�O=��9�,�<��<�������R��;nR�9�<[!=�.1��>:�^��:E����y�;��������_=I#,=�q2��y���NF�M9q=/���f=A�;�fq=�l=�s�;.s=x���==׏�Ԧ
���Ҽ;�����<9Bżvx?=@ X<%Jt=f�H<�ec�P^�֬���T�̅X=z�ڼR��<�W�<tB�<�`��$/=Aφ<%8�n�#=(Ӆ�M�;��|= ^���y-��#?��ׂ<^=4��< ���DT�<y��<����Uq�
����<�3�� �4=Q=�;�ܼR�7��("�����Eʉ��F�Y>.�6����oQ=�-Y�A� =/�㻺�p��� =yP���y<2G�;�'=iH=���\=�Y�<�1T��ּ��7�</��<>Ο��=�;�É��J:��=kn�2�w��L9�t ���r�;$=^��<���<��>�*��<��3��K�F>��Ѿ�a�W=����&W���%��:|��:��@H=�@=�/ <�܆<õI����'��,"=�Ma=�5=���o�qL>���<[�+=��=�z��L�%����<ţl���=֞h<��=W5=wB�<2WM=)"h��⻦�9�����W	�;��=���<�>u=���<��_��N=Wh
�+��<��ʓE�0��v�����b��pG=2�c=)=�O=��^�\=�V�^�{f=��$=
+�C��;����^*=�H�<Ϗ	����D{����yFs<�Ja��[=����/=��=�B=�5ϻp�<p���z����<$?<�7c��\o��0�=�Og��_<���<r�b���{=��?=d���m�<�O�:��X9'��$<�g�Ͽ���{���b���]9=�=���=:8�4v|=h�1=������;�{���������K<=����q<�=�=]��<YV��|�<��<���<F�!��UI����<�U*<����J����<4=��J��d�f�o=9&;�#�鳁��G=I�0�������<��<j[<KM��06��>==��S�Vh5��[`�5F�<��ܻ�f���A�+n%<�^ ��|!��V�< <a�y�p�>=Ǳ�<�zl<�͏=jV$=�D�<4�ڻͦ<�a^;��h=��ռ�UH�2=�YO=F^;��\�tC=dUd=�4�;pֽ<H�
�(z�<^�C=�gR=��+��Z@=
c��Ɍ=�$a=�N=4Ɵ<[W5��S�<|��</o��v��O��FF=zM-�dTҼ�m����;��=�>C=�Ƥ<��
=~����<�7����;jl	���R=k8s��̼!�A=�t=�6��<��M�|� H1<<����n=/���j=��<�<LX�;t���4=�1=��}�?t�<T����/�5<��<���<���<_�:	��=GY\���=��Z��=M�8���\���;f��ݽ���y=�����ȼ��.=g{� E��{1==%�
-=���m�<�e3����<a�?�:ג�L��<�}=�@���c:&��<'Y(���\�B#
=�`�<����u�;tUG�i+���>��4_�������8	=��r��0[=z���>�<h;<�)=�D=lА�u��;��I=D�����:���<��~��ݸ� =Q�g�w������6<�򳼉5 ;f��<��k���6=�����F�(F�~�*�;���(����:��a<hWK=�`<������N�`=@��<8�=�$O=T�=��.YE�(L�;����
/=L��eRh=v�#<י��@Q��K��^��<=�f�:Р/=�k���K=��7�j�ܼ��=ƴ �Ub�<��=z�7�4�?=��3=P�D���=a����0=��5�
~�<l+�q�y������#��+!<9_=��5=�U�W�=��4��>��x��1Z�<�K=}����T����D��Qs=Cp\�;dD����a��S8�
���<���N=D��<�]"���< �<�=x�,=R�8=4���XDü2퍺y�鼇��2���[�.�k4���5�A_B=��8<��;!�X=aW��qͼ��ļJ�$�6k�q�U��^�<�>;���!�m�J�V��mȐ<�#=[VK=�WK�" �<VR=\���?�=��a���T<y������MV#<R'F�t'q<l���2�7<�
=��_;�G��=�,=�t��Yo���!���'=p1P�|Bd������'�S=R�Nt'��xM:�V�:߁��9�Y<_�J=SlF�A�o�;@̤9Xt�[�;�.n<ȸ�<#�u=����6w@�/��aD�<:0˼�&=����d�;n$=I��K�N=�#	���������c�=d?d�u��YM�<�bK��Lw��������<���<z@<ǿ����e=ґ��M=�w�<*"����q��W�ԕ7��5#:�>�<`�7�~�5=��E�0J=4�<��%=��\���=������:�C��g�л֔��\�8:pZ==��<D��<@���!�Z{'=���<��;��h=bT�<?�T���;9�x<Z�䜥<Ƽy�=�5=!�@;)n�< )��{��7=������=rM�<�&�<�h ��I=�^K�i~�<��<@|껍�G=��ě�Hm|��,�8��;�	e=F�6=�q��g,�a���nSe=ݻ;Z{�ŘV��y&�rV=�&׼��U���R��4=��5=���<1�<d���ըu��j�R���T���:DH	=j�<���<�7h<?�;t	<�{���4=�v��A=�<FG=��3=8�<�%W<H���� u<��G���@=	�S<"��:����!��J�wG��ǂ.=�(�<�	U<o��<���<�\>��"�����*��� �W�<�"��t]<em�;��{�4��<�[����λ�fż*W=�07��^=�'��.<r|';Yi2���O�Eg=e�;-�a���D�z�<��$=�'��ֻڬ�=Q_����,r��lr`<���!
<?�9�-@��SH=i�@<�ѹ<��9�/�=��=2��<Ǉ=�8�;�L=�bc�$�#=j�<=g�<����o-�쮎<�� <$����)=���<S���c#=f��f��<�-��*e=sI�<�u<�].���� ����O��s3R��-J������U=�������zܡ;ڬ#=��x�|}��T�=/�*=�%=�N=�c���{����=��fơ�D�D=[� =�d�<��R�S듼�)=ԇ�<p�=���+<��=Ǉ2=4`<��G�HK*=��t���l��~��pR=�.�of�<�ɋ��4=)�$=�=��,=0��]���<1=�bؼ�F�<I���=�I3=JI�<���<;(��U*��T��:g�b=��k=Lw@=�<N=��<���:[:����&��[%T�Q|�<w�m����<S4<�ɥ�4A=�17�oje<��^=��Ż�R���t;�%=N���E�}�,=x!;ᾅ<��<�ڳ����<�K;���<ұA=��<o�<$"d��F��U?���P4��̅���X���?=�]�<�n�<;G�<�{=W,):�� ��):��T�	�=��;=��;Bo ��A�<�[=�?:�@�<�9�����<��+�>V̻_k#=�f<��<U���/�ػ3�8�V�й�<�h=�벼�E)�c*=N����=
���t=�=$��;_�=+���`�;���<V����w{��O�0Ek��B���>=�49="x����c=j�Y=�eN=�Ӽ��ۼ���<W�Z;��Y�[h;��*�qr�ߑ��[nh=]6�Z�O����;�rY��C�<���%W�)k<i����;In��y���-6���T=�d��
=��ϼY���ڔN<Gࡺ��; ����7����(�)��O��b�?��	[=���;=x¼7�<@��X����<�f��҆	����;!*��xK�TA���]�VZ���X�,�=����<�����y=Ȁ�<�9==@=ٲ�=�m�<M�:Lm��t9=X�:�f�zW�<�;S"�5ҼO'q<����;T=~D<>G��sU<��m=w^��1?;���	=��ռ��p;K�f�IsټZ�<�m�<��u<q��;�[�?�b�T� �&�G=��ؼ�>-="�U��������9��� ���-D�,����Z<�`�¦���Qb��L<A���y������y���E�<��4����_fB=���<�L~���{=Y�T���Y��k�<��Ѽ3u=�z2=�x"�r $=T�i���]<��?=�7������弲�&=׵<_��<3���S�%<`���4N���\�5��<=Td�<��@��!���`���`<m�K=U
.��b�,�+��ʹ��=��ȼC����ˉ=�d����<v-=�f�<�7;��:��VF���=�D8��	�CuA=H��<M�Y=gm��lD�z�S���_=0Lp=п���[<p��<.Q����-J��<[Ｌ�,�B�<�-�<�::�lW�O�2=R��}(n��g=�5໛��<
�B=����Z�<�;=?wl<�Ԇ<�g�;��8;��R�	����<; >��=�.�=�@������}�
��<,�޻��ɼKeO=�:T��0Y�p��<4cO<a�	=�,=�.�:��<�S=(�����~=��Y;��<W;<B=tܳ<xx�<<�#��<��$=bp�;�:���Z��@���Ll�83<�0�3e<��*<61��ө<�j<q2!=˂�;am��
��L�~��B=�����CS�DA��p֢�Y�	�˯��2<�&.=��@�猡<|u�<҈<��<��ϼ����&=�v�WK=F�A^=E��<`jD=P4=��<��<�=�)�=��<=�q��{Ǽ�9���6�r��<��2=ֹ
�v�1=�q@�ȍ=���:�Qܼ%�s=T�꼊�~� S=3I=|��$i=�����<p#m<`9��U;���9��R'�:!��<��q=�v<OP�B�=�cj:��C=�\=�E[�� Y=^��<�P���; �3=+Y����I�|¼jݻ�컝ٍ���M<(BH��a�<	
�!���;�u$��/1���=�a�<ea=E<I�z8C=A�P<x�-=EA�����<�6�;\@ۼ=�<�����������`��������<צ����k=n�	<hU�gdM=X�A<�u=���<�g�;�~s<�'z;��o=<�;Ue���=����ہ���E>=�A*=��=�=:��Zx}�D�<�����<I	=���<�W;=E�"<T?�?�T�-ƚ:�wa=�u���=(S�*~{�ڃ�<���<�A"��>�<��S�Ћ��dLr<� E<�����*a=��<G����<{;�;f5F=�z=�1:8�Z�iP�<%�=�u,=I��]>�<q�<�`*�	��`�=���;�b�;���;�5G�f�;\�;�'�E���pz��e�H��<�^^=^א;o�&=��=���������؝�t����h�:���ǩY�Uj=L���*)���!��v,=� = �<ч ���ϖ8��z<��=J_���%=�/��;�Ep�����@�G�;�#B�*�Z=���q��ԥ<d2l���'�ټ3�U�=V�'=�-�����L=.�B:pe����X<��T���A=ۅ^;ZV޼5�m=JsּYD<8���s�=���<�=/p���玽4}=�vi�g�<=���<�������Y�)<�=D=��x=4��<����;W��@��-=�L��F<�e5=Jo==z~�,ͣ��g=<���\==�$<|,�<�ȋ�7��<��U�5	2���=�]5���1�<���b�P��R��{L�2Sh<3	��E=GЭ<L��=�)�<���<��T=?�P=��=����]�qr�<�6�;ĉr�W$�F�=��� ���>���%��2<E ��:��T�<t�I�_��<꾉��!J��s<��<�q<r��;d�='E�<x�*��ה����M#x=����X��<�Sa�n�|=�(���B^=��v���D��'�;��	��[B=@t='g�����̻���;�S=�@=�	<��2�SZ�}�7=X���``!��lc<��<��>�.��m@=<�=r-�<�Ch�q�=�n��Ǌ�<3$p�(�4�j�)=e���L:��(&H=�B3����;���򦿼u�J<!g(�eD�<^iJ=��Q�օ=H4=���9r��<���x���h=���];8@�<�d=:o �R[�;��<F #=;��<Z�꼏h���=#��<��h<�V�<� =<��<F�c��6ؼ^t_�22<��F=��5�u�o=�(�;�Jk�,*^��H=|u��<	�2=��D��� =x�=Z+���!=s��Lg��ǟR�9��5	(=Dd =Z�@���</E=��޼��9=%�.=A(���?==�5:;��<^�����(=8�#=���;K!<$@�nL=Y%���=�F<��ʼ�����;&=��޻�Da���*�X��� �lM =.��<e:=�.)��9r<���<}T\=b9�<s�2=��1=�S*����<�L<}5�<}Bs;�����:������4=�w�|:��>o���弨�V�Z>f=w�b���A��e��G��d<1_���d�{�9� �����={�(=r3���3<E�4��;�mK�@z�8R�y�L������I�ټV�4=!X!���k<C�	=�Ӽ���<0	%���9=~iu=�.��}-=�r�|X�;Q��<�!=]d�b��Y=�s�<�Mr�5|�G�Y;�!6����}=!�=Y��<���=��p�k&=_hF=�1��Y�N�ޔ]<��,=��� `�P�6=��?=�==��w���#=�H��?=-�T��GS=��\��x���i�|�Z��L�߀B���'�I���CD�?Bb�Yp�RfK=8����}=eX=	����m5<�P����s�8���y�[M�=�:=��J�<<�:=a|!=;�A=~�컰�F���4<qn��˫��^z=t�.=A��<A���L=��=�+�;r�N�����t�W��<[JA�$�ڼ"�;�t<�lR=��S�r���E�[�+�Z=�z���Lp�b+�������5�[7~=c<�J=6�*=hF|=�vH<#�T�b��L<��?�\Q<l+�l�h=K���J$�ce�:�E~:�x����<�[��q=X�Ƽ|�<�0=	����'=����i;���5=bf���d=�5�ed<1�'�S�5����w��y�=��<�HI=2��8���/X;�S���Sk��魼H�߻7T�\&�^R���b7����<��y��=��e��-�<���L�h<󑆻j�AG��OQH�_~*=�J���c=Kp���T�P�=������	<=�>=6㊻�(=f۫<	�<h,�9��;����}��_�< δ<-��Pyp�44p�	��<H� �.�7���ݼ���=v㳼�pR=�)����r��F�L��;����D6<A�@D,�qHX=�L=.<��	��a5�T�<�9�C��<)ܝ<��0��\2���_<M���(b��K�<e�D�|s�<!�ɼ�G���^�l��;L�o��>�+L9<Dڄ<�0=~꠼�=؄��T⼐��@PD=HNy=ֶ�<��<�eb=3c=�vL�,Po;�	|��$=��Z�|q<�VH=2�=m�=<�<&�7=�5.=�ʼ����'��0$,:!Ԉ=  u���<Q!=�1�<N�;<=rv<��߼P�"<��2<ӕ�D^=�W
�qh�G�<@R<��<�ʌ�\�3T�<~)�<�5��;<�ǎ<п&=�{=�>�=�xռ+v-=p^�<ߖh��t'�������<�4=���3��<w� =�)J��j=�ꊼT��b~D���L=D�Z<�oM��m��jɣ��	=K�@�>�D�5r̼����xʼ�U=N��j-B�I�O=w@<� �S��<:!�<�g=��>=�T=�����u9�{S=��<�Ɇ�j4h��N��U(л��:&C�1b��r��a�-�p�u=)9�<����TL��M,=��.=?]�-%&=�5ȼ��L��Zf����:lL�����%�c��<�T��n=@��|(�LpY=�q޺��R���&��@?��+=�L=S7J���;��PJ�g@�<�VI�f9��"=�.�<x�=%@U=�(=�돽��-�Иټ�6���<9)`=�ZV=Tk=��W�2ts���<M�l=�����&%=�<�wj"�<:?�-���;#.D�4�,���G�(4=��J=R�_��T����;�h2;�h�<�B� 挼�\=�&׼�.s��O����,���ļ j=+L��N�=@��=AB�e2=�){���=�6L��B����;Ι���!�<)&=���Ư;��;��<pE=�t\��+�<�� ��M:=���-�M�U꽼,�l���@���|^s��K<D,��V�<~�:= ��<G�M�F��<��5��_�<���<n��D\X��I<�>�7�sj�=��\;z�&�E����dZ���N={�߼��(<8��=�J=#�<�<^�=�pJ�����'�$����;��Ϲ<0aY���U=�"���@=*])=T����r�<�̄:�쪹�#=���m<��ڼg��<a�<l("�e�#�o��<aՕ� �=n^�;3w[�StN<����+�!F�<�e^����<vL���=� ;=q+�<�H$�RN���=�f<2ÿ<&p�� =nU�cs��m�<�Lm�����M
�n^�������b�7Lb��I"��"=�и���<D�9=<� �Qv=J��m/<��
=���9�P�<� �֞
��[�3E=��`=Xr�=�!<��� <"QK<Q�޺w��<�_�;�#�-�E�%xC=si`;��\<�Qܼ�u�='�;��8�]��<�=��4=��'=Òe<�p=YI=]��Hې;��(=P&W���=�L<脎<^w�<d��"�$�>���"h�>�ļ�f;=�5O<M"�=׊+���W�ͤ���<*�=� I�k�A�G��<Qf����iny��uT=�=<�#�����Y���Eg��V���e�;��;7�9=:Cu�d�=G*���<RU���SE��%?��D��5J$�S�I�󀃼�<�"*=�=�<"S�N�����	��\��l�+=�?���@�<��<u�ƻ�0�����(�}ud=�=�Ծ��0T=��
�.M1;������2F=Z=;�)E=X���!a�9MQ=p����h��Ƽ<(�<~�Ӽ��t��چ�5<L=5�C='�<�����.3="��<0�9n7��P켓a@�h[��4򼺑�<�\4<6�=KŦ<f�]=��=B��Q�!=�֥<�==��=j4�<��O��	:=��<��	=F������<�ғ<���C���9�<�A���C=�<b�&=�4F=(�;=����Cp�<#����}�>��</"�:Kd=�=����~=�'� �w�S5���Wb����;�kq��M�5<�H����v���C<g`G=?�1=�X�<�Ғ����<���rA��I=,e�8�c��C4=g����{��Fv�<��;c*=���=#�~<`>�<�e���<���R="0A=*�<g�n=�*�<PpY=o�v<��DżcK4=E&�<�b�{��<4��;%L��>�<��Ļzt�<
*Ｗ��`����<dJ���<xvȼ��4=²�<D�J=*�:��<��=D�<O2=���<�<5F���<#T�Af�Dz��T$�o� =�:�;�5=%Y�<.�ۼ�b�<��:=2=|��1��*=u�b<�>�Q�yR�<Q��<q�������H;F�
���Z���=�\��19`=�T<��<�f��27��3�9�R=�=�p�-���.�=i0J�_;�e�`�_�d<dF=5 �Cu��=�n�Xݭ<�1�{U���=���;�Züf�\=WS�<�`n���S=�K<������<�k�<��,��-B=%=9�,<�R=E�
���b����������=�ĉ�ΰu<�=y4���;�)K���,=X�g�C?1=���<?*=��<m�<C	=H��<u�=g5<"�'�����q�E=s��<勝;�K=p�C=�"=ki=�w6=`�n=�����<pED���C<t�߼��<Ly\<I� �����T<ج�;���<�<Ay(�f$�Nxb<0��<&�=%ļ!XT�b�<�=	ơ<������}p���R��g	����=C�o��q�H�<�@�">Z�Yb�<g���?B�
3,���c=	!���3=H�b�W�m�����$c<�ꊼ�h߹��'��Z=mC��[<����Eb�:h���C=� ��o�<�ù���	�S醹����)����j��<.#r<@s�<�ST�btd��=�1�|\�1B�p��!��jzż���<���;�a�<��<D�`���=v'�<1>Ƽ;�;ĳ�y�F�Ye%�u�2=����}z��U�<��/;�C=��R��O2�������ͺ���;>\��r�<W%�7�;�F�����s=x���F��;.S�1+=Ի�=�eq��l��`�<��X�S;���ּ��<�¦���A�c�&=�BW�J�U��m������n=�qG��&7��=��L<�xj=m�;C�̼Y��;�z�<��]���= �<h�&�(�����-=��������4eS��:����m�<�?m=�ty�ތ��C
��Ƙ;0u��6���+�X<��<$�=�?=$��g��Q��+=�/�;�7��=�<��I=b��<S���=w*F�{4���u���k�(�<=F��wB�<�BA=@�ۼ�U,�Q|�=����k�Yx<Λ���<�����y�;=>L���/=�K;��<�Sݼ���<�*���(ht��C!='��9�7���9(����ź!{��+=BsV<`��<=!`<�X�;�����<��R���8=Pw��.�]��<���<��:��l�9�|�;��<�?=A�j=�-�<�n����<At����j*n=���<2(j�t��;hpq��n��=�¼�By������=I:!%�[i!=h��C���0�Z=�G����=!�t�=��=�=����u�#=em��|�:�Q<��<33�Wa�:7)j�;dL=i*M�g�J��'=�}w:u7=�:3=#6�;�#�ݪ�!=w<�=��V;$�=��`�U��L�f=HUG={vz���l=Q�T<~�\�]�� ��8z
���R<�I��L�<��%=;���;�<1�<���o��<�g��(������l<��1=�L9=8�ʼ�'켃�h=�����H=Դ�<�Ww=�5�<_	߻��G�ޱ�i�(=
�3=����tF=��aڼ<'�f�����Y� �E����2�\��O=��	�b�Ȥ=��!�;ռ�^	�2g��x/���q��_==AZX��L9�[x"� X�6� ��1l<.
�<((�<�=�6<����Ln�ɕo��7<�T��� $< 0�S�3=��z<I&ϼ7�����F=S��;��=�SK=��<s��<�Jv<��ȹP���!`����<��<��ջ��{�qkڼQ�����<u�߼��;=�]�;�$v�n=l=���i�G�ļ��7=tqD=�م���(=��=Q�Ǽi�s��\���>�BJ=�aa��U�?e�«��{,���<�$=��u�A�������]=�mu<�`=�\ֹE�7�n|<]B�� ��&���<�?��Z7^=�8=|�G<XN;&`;�kx�;ط�<2�<��<f��?���H<�\(�d��<�Rl;yo(�]\<��<��J���T=���n�W�yL.���$=]7��j��<r�@�u=��p�����Y/��%�<�����!�UC�;�D�< d ��CN���t9r<P|�;p��<1=EF�Ϗż�T=H���D�<㮉����<Q��<j�����;��<5����_�<��h�<�}�qu��w�<C�<U����/�O����:~Ѻ��#�"�e��Ⱦ;��׼~y�\M��_Q=5+ü,�����P��y���=.�-=��c=���;b��;M��;�̼[[�<��;=~�<m?1��Ӽ�=��(���;��<H3=��>���b=�l��v�3�Y=��<*M��n8=���;�<|�̼U�J=Q5.�,j����#�m�D�	��Q%<�|�c ��y�Z;6�u<oZ��Fg����=�r�;�t<OP=�<��ۼٽ?=�Z=q�����<�t��Զ�<�=����$��s=C.=��l=!H< ��< JL�j�E�E]�<��=u3�=����ȇ=Yk<^=�|���G�;����jW=��G=��6=c�^=MC�<��;6=߻=F�j;n�+��J�~�������5��1�1 �r" �h�"��������<\�nw�[u~���ּ0򻙗�;n�o���U�����.; "�<�ʇ��a���:7�sH<i���pe5=3]F�5ھ<���%��ώϼc:���.��D=^� =�Ҽ ����Ƽ����'?�ղԻZv�;���<�x���><n�$=������I�~O,�GN=K����0�Tɟ�ss��S<�::�(L"=��H���h:_#Q����m����}���=��[<�A�z=�;�>Q��#��\m=g�������7�;�u/G=�<	=mXW=��ڻN�W���{�\JX�*Ȇ=f� ��"=�˷<��3=V	=\��͝R�7�����Ǽ���<-��!���<�=
��;�ye=�T;�3���F�J���BE[�͝^������%O��[�=���<c����<>��<m^3=�!)=�8�\R��
��<q�¼��.=�
���1='+=�ߨ<��Ѽ����V=��<鳼�1�b��<�0q�c�	=@�<�7`��q1=�9�Ó-=\Z=R���%+*=\�r�XS=jD��6=�l&����:�-L�<�<�g�y��<��߼�x�����<��u=ui"=3����<�g��EF�<m�<��[:uU=H��[C= Y�<l���V��jtf�ZN�<0�M=�n<�K=�N<�#���;U�<�R�����~���N=�_W���=�:d�f�2���e=E��|7>=�$�=*Ú�7� ���L:<�c�o�����V�?�<V��e�(<�� ����<DqM<"�E='X3���=����ւi:��l��w��QW���:<b"�<��������3=%g��Q@�<�3����<B�,<�oP=RrP��x=���<ԩG����;�#�<t�#=�`;n�K=�����l<����=��<^z��=�S�O�d=�R�� �3���D=��[�T������^���r;;֒��	D:��N=��ļ�D�<4�3����<�[��!\���$;�.<��E��I��\A��<�t�<۳˷Dq&��ZO=S@=뼋�x���:���軘[j=q�<�=gx���l��BY=0<�5����7�Ul��~=6�<��6=��6=�D��2<�M�<ɸ,<�w��8=��R��R<�=��#��� ��+�=+���=	l"�P�A�[]8=rW=�!8�TY߻�� �r�H�c�'��L�<u�ͼw�2=\�u=�r7�"�Z<��=)|�B]��28���=�8=��)�E����+��	%=���< Wu��1m=��<�+z�;ޒ;�6=��=.�>=(�=ֱ!< _0��D;=�G�����k�!��ޯ;l߸<�M��e<P�P=�𝼉Gz�4���+�:����Hf=����J6�ݐ�w�V� @`=�*<X�m=�S���D��(�n�κ�&��R�j]Z=��1=y�W��`�v�<NV5�_�<�=�3���s�<�k�<׶�̪E;�0<ysH=�)���ݩ�#E���t�.<Hw�<�}ܸ�f	=���)�a<�55=�k9�@=Ko���dd�/� �U�<G�����=߻)=��_�6�=��8<��s}]���C<1T5=�DѼ�UW��+�<�=,� =ʫ�<�&�"1�U��<�ڒ=0=;����	+=E�>��4S=uz��_;<y)I=�Ja=FF<`e5�|�<��<jP=cb�����.�<�Y^����=�A;�~a���3=��A=��Y;��<mo�<�9=�g�Ļ���<Mym=��;bT=ɇu�Vg����Z��S�<�9�<��;�ُ�"t���d�����%M�{4&=T���Q=kjY=��L:9�9�Y����Y��)><��8=�$;�,��V�<p���&o�}�\����9ɴ���b��5.=gq=&Q:=gq�9�����;{>=u`�`���<,E�<�	8�f�p=`Rm:��<���.j=��Լ!�m���]����2k|�V��w�<��<���<��!��{��q��g;=��'�Iɣ<^���Ĉ=��<]#����U�<LEA= �'<�{</+�=�g��Շ;/�r��.�KN���=�*��g�*��<��<|����(>=Q=]=$��f��F켵5�<^�<�LO<aԼ���;F�b=�l=��"�g��<��=`�l����=�_��N|��>n�x��M��U1=k��;�h
�=O]�����dR=�$=��X;�|ڼ'��<�S	��((����<|n=H�:=�(��=�Q;2��6��n=�1< �,=[B���?�6�h<@�$=�AμN�=ʋA�$(C=8�ͼ�=�QL=�i0;?����;r�`���<A�P��><��&=X��<y<3=^�=��%=�*���X=0T�/G��7=��E;��/�b#�Z�:<cƿ<6�;�}��iD;�������;}�J=ӗ0��M]=�� �s�Q�=6|<=���a�<ma=������_��<=�8�9�p<];?<�y='��<7�@=�$�.�g=n��� �x����L,=�����o;H��ԣ���<j�c��s˼�+4�J��<���<b]==we$��<.#��#�*�����>@�VS=�-����<�[�<B�<�[�#M=�%(<�&��{R�&��<��ϼ�<=@�ʻ_u����B=�O�;Y�+�E�Ѽӱ��e�6��,=��=5��|L>�>�q=�Z<�ZJ<�݆=�#*=�)F�ql�:#��/]���n-=����oL���:ޟv�*�=�e�<����m��<l�<��w�F �<�ּ��:�{��<fhL��K'<&�2�l�<���P�P	v�1�]�]�e��C�<'���uk<� �<m��I�6QD=��8�kH,���;w�O�s�;���<��ke.���~=���f�	��*%�ouu=��(<�L�<s��:`�g<���i��:��輵q=4�a�
��<�N�;@e)=��I=K]=0|,�.b��@j�<#M;���O�M=>ؼ�}=od�<DIR�*�R� Kd�o�<���;�C�f��`��<�J׼�S��t�qb�<d9�L�=VO��=p>���ތ<�/m=��n;��ռ1Q���<Prx� �0�=&Sw�EC�<��<�) �| �{���0�=%��<b�%�<U�D�g��<"ow<`Y@�/+W�^S=G�輓Jk��,B=�3I�D�A;z�A=�<�|(=�.=~�h�<��㺞�/=	ZT�KW����<��=U%�����KL�N���R;���<��F==������O=7�Z;��I<�W�;�,O=_�T�e�=�ja��Ҡ��v=
�;��xoػ!�=�ɀ�ǻ��T����=��,�:
�(=},"=�j<���<<�m���v���:�B̼;=��<%��o���K��$�<
�<0_=�8��<��޼S�0=�Wٺ6u�#S��CU}�&
�먇�F���e(�ཉ��
<i}=�)=�LT=�-���s=|+�b[=��<Ԋ=6�5�z�=��X�HV��&�<0�;�f�H���';���<��<Or�2}F����<���<���<�L=w�S;��;M��<�N;;�&=d'0���s=?��:<Ӄ��=�Ϣ�z�8=.=�ۼW����:�מ��03=*�<}n&��iQ={�l;Ӿ2���L�L$�F���<烣�*�E�#�N��O��� =����緼P(��x�00= A���&���=���<�<�w!�'	o=. ,=�=�[��$;@��qI���X<�w<��=n��<<�X=��A�f<#L�:|�=���=�w�<��<2'=P�]=b�<~y�:���k��G�  ����:�.�<=�J�6����9E=�ke=)n�<�;���=���<�3��mȧ<��s=ti����<��}=�G<K<�Z���q<� =6�$��M=G-Z�1�<�|D=-�<��\=��J�6�&=�%�<�=�i
���$;G*����<�~;=G�<�3Ά���=wZ8���=�S<��O�<6=�&��O�gf0��w�<z�W=¿r�W��I�W<̡<�=<������=1�=)s���^=i⦼���7G!�⫽��#7�GF;�!��AZ=��<O{y���<A�>=��V���G=��+=���;�8]<_|����"�ǽI���6�ܸ?=��3;e|��k�Ƽ	R���̼�WM�h�E=3��eG���u<�� ���`��Nȼ:�@��8=�<�;�U�=��<�B����S<��7=e�==�=xl'���P=�(������ֺ�^e�&�n=�y=OG�<��=S##<]=�ވ�e-'��b��m>�b�Ҽ�ߥ��_�'<�KO��e���?���	=��¼�
��w&�:xG�<�c6��{����4�����pѼ���3<�r=�a�b-�;�֊<�����<0�?�D���=�sY=r����m=��;	$;=���Z_=Ne_�ɟ����l=Ý�;�,T��v=�ļC:=�.=�0;��d�<={����<I'���뮼��S=w=�؆��HD=V	���i���޼b�"��\���}`��=&L�S䵻�ş��_�<���;P�n=�;:�P�j�
�G�iH�<1�˼+�=�k=�=><\�Z=�0h����<Z��<�"�<ԣ���==ċ���;��2��ݟ��]<;Ԑ=�C=2f��n���j=#T`<��Z=G�.������<I�0=O�=$-/=��=!��
�<C�?�H=k+=W��=�]F��Ǐ<pM6=��X�rI��F�J<�%+=���` �<fl�<��t��õ<} ���W�=%~��oM���X;���XP=3�p�h�<�"w���<������I��9=z41�F��<s.	=��q��:e��<.�H��q���>�=I��v%�<D�������^K]����<�/=MۺŬ=[
���h�y�����Fh���;�^=�=w��:UT=�I= z �t�\<r@�b_=�,N=������2��.�b�)�1=1��ǂ��&���0I꼤{�:�V$��ں���9`�U���-��Yh:�����r��Lz<n	�=t�=u���P�=�r�9�<(��~���\���b=�4T�3��@�@��鼧�=�HJ<}dܼx�=��h=&7���=<�;��#�;"�ӻ4d�<=;����<���;��\���[=+F:H�3=���;z�?��D�;�f��F���l:�v�J�Pм�F!=�<w@�,}f=�j=e6��>�R�;�i*=ڸ��R�`����<����k�.=�nV�J�<�]��h�˼�=\EY={�:<��R=�@��ٺ =H��<��<���< ��<����x����I�}$��j�g;�<�&�<�F�gRY��?� <�f�8"=S�B�]�U;�b��
��ͩ<��@=q��<��׻йZ=['=mb)<��(==b<HF��g3=O��<]3�<�:�<�`1=��<������;v[.���K=o�ܼ�꿼�2����߼�J=�z =[!=�BX=���e�5<���!i��q�<���<V��\�/�4��|U׻�fT��菼-1g��д<b�h��mV��=O�t=}��b�<�#��<޼H��<��<�.C=��^=�E��ڃQ�~yH��4�ECR=?�5= <�>��bp�;C�F�zhӼx�i<H�4�sp�<J��::�(�3���)���EF���8=y��<��N��ie�V=(=�S=��>��P=��w;�m���=If;�]-��vw=�gP��bH=��{#�<� �<�j�iO=2(���G=c�5=F�d���&<O��z6�;2<o�G�c�ļ�=�<T�+='�<8��bS=K�.�'JU��\��2=v��G\��*=%x=0��bl'=�/�<W'N;�����M�Nד<�J��W��M�K�s�v<ٯd���>=M�<o�$���2=	$�<^���7�<����ϙ;��<�|�;��;>IJ���~���<=���Bu��P�LvX����<�B=���sI<�rZ=
����-�LYX=+��<���v�v=�2=��;ue=%w�l�<�S׼e�E��#%=N˓<�d#����<̪J=K��=�<��9� }���OK�=d����<�Q������ܼ����w]#=?S�<��ͼ�ʹ��E���(��ׅ�<h�<�?W=4���b���;�<Q������;�\5�S=�ኻl`���nf��b,�s0U<�Z�<�E�;7�==�A��,�H=,�!�ka�<.�	�_�ȼ�#�'E��tK�<�k����"=�Mv<�FL�ϻF���e<|m4���}��-�jh=�_�,���p�^="�K�˯3����<��;/�o=�[��xac=���<���<;�5�0�J=���Z�<=0+D�tT6�7g�5;?<�"`=8ZڼJ���:��p2<��= ���JL��1�8�'��j��}�I�o=̀\���G��g8��� =�%�m�<����tf����;�<���:H`׼5*�l�<Eq0�˚p<b�=�IL=�B仕�&�Q-`��n=W=�Oh==�=wA�����܅���=���N=���<O$9<��:��Kx���Fh:=�u;��0�<���< ;>���P���V�*��:G�~����<s)!�*K<-e=�8P�S�N�A�[=dM�Z�D���?��3;=��$�ҿ�<}�<7�!<<芽�����=�h3=�HT=*��1<aPu;�l�C�/�%P��o�=��T�W?<�������<~�+=Л:�L<f=,ee���=9�[=��j�~�����=�yk={O=��6=��������D�[��<��D�U���L��O�@�}.s<Ȼ���9=�X�<�J�,켾�k=�@a���Ż�AX=�o[�Թ~Α;Wh=��8=de�<��,<�n7��*=������A=G��<%I�<.?#��[<F.�{s=�=�O���p=���<��N=V�<l�=���<7�K<���E%=O�-��T�<N�;��\��!JZ<�)߼"3�<s�n��[�=1�<�*V=�:��zA9� �=ri��0�=w�<��U�:��o>#�ߪ<*�:�һ�9��爆���b��<��<A�<0��;��T�<x7=%/A=�7޼�k�á <
F���iӼ�8=sԽ<�sx�A�<�==�C@=��m<�kɼp�9<�8=�}��Z��y=`K1<YTy� �H���C<-�Q=kJ=�w�:p���zB��'=�=2m+��;�d�<
�.�oS?�9,^�J|���J���<�]L�Ng�	�1�^� ��a<��2=��;���<*f;>==���h�v�K-���t���M�4K�з���μF�9c����� ������lN=ZV�[U#<i�L=�`==D�ּ>	!���;��L�h4���<(j��i��:��;`��<��-���N<�E�`�=�@\<'���YT�n�<b2;�}a=��ּqT&<���PU�;�x+<��m�h�<r�[�*~ռ;�g���d��	n�M�J:�*�9�,=��d��	�J);=L�/=�S(=>�	���:�������<V=3F˺�A�X?�<.<|K=,�<� U�;~m�;�t=�Я<��M���J=�}*=�e�;������׻B=��<���<��u<�]�rk=�w�O��J��x:�<{�껑I=�]=�{ =$%,��׈�K����<�y%�i�=�I;����T=��@�Uw+=Bώ��� ��y��)�:)t=V�a��3:=��H�%ҟ�F�4�!%=�[]� E�r���m�h<�p=JOu<�G�g5=��F��/j:�)=R�=g A���"�M(%=°�c�t<���<{o���b=��<t�==�*j=-�=�At=�D�<{G ���<r؀��苽��su=Q�4� ��<Ɗ��y� ���
;%��<dD:�o�я0=��;��=��e���5�p��#�c�DG�������5����i�Զ���=M�c�U=�<�;$Ӆ���	� z�<��%���+�<Y[����>�<B/�d�{�`��7���<?��;��=��<*�<�A*���<��75�L�ۼx�&�@n:�T��n����-<����� �f�a��]=gݼ<C�p�B�[��	=�u���̃���a=z'��Մ=Nt�<�P�m�=��:u¼��=0���Ȼ?N��n�v=
I2=�`�;�<P=��[=�|F=!VM��f=|�#=����ػ�{r�A�=�>=N�:���<ߛ���i�m�<�~�:z�3�_��9�<��<��G=:*=��-�;��<�ؼV$��摼���{d=�5�<��=��=�=�:���Sp:J[���K<=su��Z��X뼙�Q=Ɖb=mbļgl�=wv]�je����6�^�,��?Ƽm�0��n����M�l�c=���=-�<j�M��P���5R=�Z����:��L=9�<�a=�=u�;m��<����D������i!��0y�<�1��ݞJ<�m ��s.=�b��O=g`�Wo����v<�Wh<#��<K*���� ���=a�*��qD�sb�+d%��_��EZ$�G�1=P�=��<��0���ʼJ��2_� �мL�����6�~���û�b<\�Q��0S��	=q;�H=��<���.Q=���;y�$=b&ʼ/�=9SE���6�S�&���<����Q����x;N��i4?�k�=~Nw<�3=�?&=z�]��-=�	�����Z=��3�G䳼;W�<�"=�<	I���.V=�$�<�A=���Z=[��=��=~�	=�e�� _�t3=�',���O�P�=�6�=G��m���򺙲��vd}==��G�<�̕<�"��fg��<I=�!0�=e�����<�@<�����(=s�u��$��$�0�.��;\�8�Y{��)8/�|QC=�cb=��<#��<iXż���y?�<��Y� �u=N]���&A<��P��~ʻ�E��p����ey����)O�<�J�e�8��y��!!=�yS��VX��� <,�}=�TC=�g�^�-=����ѿ�<�](��ej����5�w<m���y�= ;μJ��<�r�I�F� dD=q��S�����Dv�H=�!�=Qs���5*��������/��(I�@t��PΜ<F�E��;�<oqn=|�<�L����;.ͅ=�(�=Uk�Pt	<���<��t�@�¼&�%=�w���0�d8�<���v���C9�~�	<OP�Z�=,{����{�:uz��z=U�1<�ޚ<��f=2�=OR3�]� ���<��=9Y&=���!�=H=��&=���<-�;O�+Xq�����I6�Xx�<��=�F�<!���;�o�<j�'�U�F��Y�<�~%=�c�7v.=�:/�D�of{��L�:�.k=�-{=��9��<ǘ��
S=L�i�ۂ<kb(=�<�<�:��Ѽ�(e=GR6=��.��DJ�sv;@F�<���=���<�р<�z�V�4�q=�W=�n����ʼ:6ع	�Q<F]�V���/�;y�<2`�;/^ȼ��K�k��:��(� �0�o>��=4� ��"�<zn˻�ͺ;�8=�v�T|<��=�XV��ǉ�j������͝{<3�X��9�����x\�&4�=��<��w�ｽ���3�qʫ�t�;oҊ���\�M����=�a$<}3F=��B�;}=Z*<�xW�G1�2U���?�;���t2=���<�Yq<��żXt8=�V==Wj.=�+#�~�#=��R�.#��-%=R��<�E=�]��k]G=�F�<���<���<�E���= �<��f=�w��A��<��<�裼wL?�YL>=gN���3<mL���=�َ��==�5�<^��9���8o�W=٧��Ak�>m|=Ä�<e��<p�;��^��c\=��;P	=��2=ާ�m�<s�a��>���L3��#�<�9= �< ]�<
&�9�?��-<�6J�*a߻%o�<Y�<�{�<Μ�;vI�+� �f}s=*S�;o��<M�û�oC�=�<�b�ofм���:��+�����m��<1��VYW<cw�<r�<�4��"/Q=�U���j��e�<Kޟ<�<4�(��<p��<+%�<<u9<8�S�R�M�ܽO=�w-<A�꼥���C]C�حA=l|(�U�>=�(�W
=c�_>9�(u�j��=B�=�~�<�	��\�l=�?
����s�<#t�<0���(�4��j%�VV!=��D=B�<�d(=}+P�5�<8ټ�'d=�*��$<�p��1�6�|v�<j椼�(��=o���:=D�I�YՑ���;�����9���S<�-��4(�ƶ��)o�<�$|<��s<�]�:w�X=kS�<���l#Y�D�s���<iBҼ�=�C�<y�G=֪�5�O� �0�Z!�J�F=��C�̼�<A
�<���;Gt�=�V�<L���n=��e=������<�b����~������;ܴ��M�<eS��|q=�+����<��</�w����#���
�L2�<j�B=��&�.w�9�<���9���1�e�+xg��}=�����ć�U{�`�8�?0�<)qj=T�w=A#�Y�N9�_�;=y��2�b��<�;��D����<�8:p�<�(�<lS9=�.'=��j]<��-�_)H��'<���<�]��]��[V=h;�hؼg�(=��:={	���N�<�����6��~=L�ܼ�oD=?g�<��;�s��/��H���1�<��3=4-_�hgZ=��w�+��mKV��'m;7c=ej<Hd�����<,�<=���a>3��<yY=1b��1=�(2��p�v�ټH=���\�<�]����<��p��}��C����b;Y��;A�H��������K˼❂=���=��ʼ�t�<S`���h�o�_���4=b�<u�Q��.ż'e��@��L�!�;=���<�����������0�`f�<v���� �Ɍ;(�o�K��<6�Z��Q���<�5:��r=�缴�=��F|��=[\:���&����؅;���z�ۼ�)��L&_=�P��?=@c1=�a�<q����;��<i([��$?=���;�g=+=�7H���=�����H�4��I��$=�5<�Ι<7l'=��^���</�z;q�9�Nk=����N��<�����G�Bt<=`⊼��N�h#=H�=<��:?���r*=�����)=X'`<�*=L28��Pn<wg=g���B=#��<�[��Q=:讼�6<,���h�=A�M<r-�8�2=��ûrjK=x�=h�G~Q���=���;o�(<�Hֻ��7D����߼jU�;��<��K=���<2W�<����I@�<�0F�8�bW���z=�k�<��Қ+��R=�Ӫ�y�(=˱�\���_2=�(��:=�o��1�<�eZ��k,<�T��<�v�;<2
d�����;�<$��A,=��<�[�I<�͟�	�<��c=�[c�m�����V�5V=��ƻ�2=���䍼T�A=�	�!�=��<���<����;^=f)=�\E�)���L��:���<�Y���҂�|Ǽ����#P*�hє�u�ü�;�<:�=GCq=��M���:
��֮;�H�����Zs;��<ePW=?O=��q�6�2�o�#���3=���;~I��r����%X�[=<V;�~=d�)=�˭<Ӈz����<̧1��~�< '=G+<�QN�'q���8��>\=��!=����<t=��N=��)����5ۼv�i;��<=��Ӽ�O#=�4�<��;�`���
�=QU=|z(���:��D=��<R%==Bd�<��U��
=,�&���=�"=g����Ҽ"�˻nN=qzY���<f�7;~se=�c0<;���,=��u���F�~�=}��� g��y
������x���o#=��Ż��5;���<;0R<x@�<�=td<= �����h�<$��:����18�<�Լ���<x��<-��:K�n<�B�� �W���^�g�+n�7���'=D�Ѽld<�X�<�ߺ�����)<�sB�ZG.�@���("�+=�kl=���2���
�V=�C����H<ģ�<�� ��xݼ`���Œ+=���<n��<����i�,�Q��;o�:��(<�-=�=;<�z.=��$�����˜<��<�S*�wx2=1<�<�e��ѼD���d��4=�s��i�<�`�˔�; �B=U�L<�7����
�b�<"�/=�(<�=0��6�<��G= +ļsP=���N��;T়��::�<4��]ۼ��=�68=�g=g>����B��$1�ٙM�K�<�Y�烌�C4�}gI���=tZ=��?=9�+i��
'���	=��g<dh��a@=�����x�e�F�Y7�Z("=#I=���:��<tb��y~�<��<_�=	��<�N¼��=\a�;T�+��ż&�=���+=Ԉ&��E=��(��<���w=�	,�	+s�]��<L���gF���N�!���q�/:\ɻ%�=�8��� f=��Q��_H=l2v��8�� �����&tz��u=@k�<��)�Yv/��&K��Kp���[���8��;{���<�l�<��5=@ϑ<U��;)QK��ү;� W=?�=�v���@c�Jz=Lw7=�S���g���K=� �Z����Y���ռ�������:��<cb=xR��8p=t3@;��=���:��0�|�-�|�y���<?�
��c�X�a����<�5Q;��Q��<�wH����Ҍ#<H�ֺ�ĸ�Pc�� K�L6=�4U�CɼC���z�N=�ػg�<�4�<*:���m�/���9I=�0j=��=��3�����<t�c=Cǒ;�n"=�X���!=��r=���=/߼���˼�
<��Z�/�.=�~�;*o�8�eu<!C=���Rݼ�8e��*���漼�:�<�����^����;���W��g�<9�n<�B=t�s<���ɠ�fm��#���<���<�D=<x[�;��>��<�<97=Y&��E=��;��<� żs򛼧�=!�мw�2=D�>���o;��M;��=� ��U�¢�9�I[<�=����;����@��q��_� �z+=u�/��A��5_<A�S<�8=~�v=N�<���9�f=N�ټ!��UzP�ɼ�@���%=�F���8Q��t=��	=?`뻓S{��2�<-�X<���<��<��3��d�<,��<�!�<ZI%=���;l%�/>���w�Lt�<�\���V=��%��I�c\=d��;]*�<%���1==J��s�����<��A���b�!Mk�ۮ����4=�P?��`8����<ף��Vw��	|�n��ե.=\�q�x3-���=��o=D�=��C=б�<y#=���nt	�ѷ=�2���r
�G2C�<�-��v���·�~�)����;���8_P�;UӖ;�gӼ��
�f�C=�<����<����r<T�1=��ϼ��<��]<���}�);�V;+�.<�/%=�c�<�C�<��������<�!�<���<��C�X=(�`=\ �=Y�<���<\� =m	=5[	��P$����<��W�(�=��=�X=v�d�X=�eɻ`��j���@F=��m����en�>�4=&�	�t;��)�;H* ����;�}n��с<�g߼_�$=�9�p`ʻ)5=2�<|��<�]��ΉS=�9 �XG=;HX����;�浻�b=�h-�9�`������<!���=7&=��P=SG>�H�=rHk=22c=n��<�=�F���dV���Jz^�r�<��5I������@�<0���P@5��nh�֞<EH���Ӏ��:��"�=�{�d�`=G�;�����<ףT=��=W ���׼��%�J�n<�}�<��-�U�{��=�9�=gLL��(����<��<G7���W��=� =S��{��ό(=�)�<�X���<f2�~7��o_<tj�<��,;���Es�<�<M�9�����ݼo
,=�f%=��ۻmX�l꙼n� �_R���ּ"�G=��<z�/�<�)�kr+=P�=�ɉ���1;L=��<	�%�=��;�>ż��R=򦘼c��q� �ީ�<i���=��h�6
�;$J��[�͓F=����j��g&�f�ؼ�I�b�e�KV<��/C=�xW<�?��1Q��� =lj<J�<_�˼�%�<W��<	6�<�J�;��ۺr��:L4.=�~;��޼A�&=O/=�2K=�x��"=�n�{ԡ<I��<�W�<��z�d���h����R���t�a����W<��Q=��:>}����<�MM����<g �����}˸<�3��u!97J��z?���ͼ������\���RM�lv��O��<��Ӽw8*�k<��O�s�H��0꼯��e��<�-<�Δ�<��=�;�<��<��<�R)=@,=�p=j��;*=�O�4�A=e�`=�`=?�T;t�!��C:�Ik�f ��4�k��©��8P=� <=a�+��o��dz�rvC�a	>��D�����0(�<�� ��N< 3���O5�$+=#z�<�V�;�<v����q=7]��w�;�][�!��� ��s�=��':��C����X��+T0=ll9���e���a!=��O��#$�^�=�/=*f�E�Ӽ]���Q���	��L�������5���䚞�8<���=V��<�A��]��X�v��zC<�n�;mY�<�<<�2=�7�.����;�Ep=�u�<S�r=R�1�T�O=�=}y$=L�;O��<l�=,�=.D9={a��|��R��X�<�˶���A=�*�H�<�m�;�S�N��/�[�-̬��R�<%�<�x�l�4=eK)��T���n,�&��ysM=�Y�<y��=��<�s�<��4�!͂���Bk�<��<뭇<�}�;���;�\��/i����7��<�=��A��=J���Z<��|����<�^C=��}<D?�<�`��ӛ?��;ռ�7��['�<J_X���<w1���p;��Y=�]^�:#=RcM<���;�Z=T�;��];;�<�Y<ɔc;� �<x=�;�9�Z�W=���<Y�̼21�D�<��-=j�n<�� �Q1�<��a=�� ��S=�=��F2�R�IW�;>�<~k�<��O<WRV<uHƼS��(=x�?��G<[_ �TI�<���xR�<%h<��ϼՇ��>~��5�<}�r����;ѿ8<�+=+ =�=�|K=�꼾Mn=}N��3p�<}�2��/��-q��;=1�:���=\G��mab��"������T=�i�.xF���b��x��
� �)=�ϴ;D<�g����1=�x�:��</�<ŧ绋���f1���.;j@y=�Y������D<�l��<�ҩ<�����A̻rGܼQ�=�l�<���<Y�'=�	�_�=��9L=>=
%0=��N�z���AS��Q&=�=�G�<,�D��`r�Wa�<~�<qx�+���r�(����è�<�oG���=T�J��Y�;e����/=h���Q�޼��伟����*0=~x����;�W�E<c�D�Z��;��:-vR=���;6/�?9�;=�*=�W���'�8�	�x���gD<ڻf<�L<~?�<� 6�^
�76����I�uM�<�ǂ;e�<���<�>W�n���K%<�}��.rX=��;��g=�<g�d�=�;�/T��!E�y�T=kռ�"<�H5;�,<��M���V���9=E2�<iM2=���Xۼ[�:=��<���W	���=}c�$l��%�@Q��,1���1=q �&jg=?
���;�ϼ���<�=%��`��=7�?��¤<S�-=���ť <��D���k�F|�<�T����<[�$�kV��׺�<8B�U�,��)%���=-^�<��M;N$=�J1�Ć�SG����<*.�Ɇ.�{�=�ܼIH=�T��'ڊ<���<p�=sDn=}<`৺q�5<���<�Mr�(l����P�+����@&��sW=�M=�.=���DI��;�E=���<��2�J�ʿ\=�yD=� "�������w�=	�1= ��<�^<b�6=�Q=(ļ��;I�<�t1��9<C~��9t�&�"=�= ��o�<���L�=t�м�c���<�03�Ƞ�;8�;rS)<�ļ<����ˁ�����_;��P�=��<4I�1�p�4�a<�~Y=�<��X<r�q;]�8<�_<�3�9�ݼ6r��:μ�f���v<cg =��C(����P�̼��;�C}==����mT=�<�1W=��<�g'=y~d��Yg����5�T=��;����M^O=��]��+D=`y����<�q'=�o�.n�<a$��^	�<��;a (<[1��N��<Ax	=��̻%�^=_=+0<��޹>4n���E<ՒV=|m�<�<;�eF�xG	��o�<`�)<�<:�ʺr�4�D=>�$=�����<��(='�)�筲�5o�xB<LBO=�I=6�Ǽ�Rڼ��)�mEA=-/=�D
�Dܸ��f;�X=Y9��3�#�1��5<�N红�<�&;�$�:@n���J=l�O����<��<��=����B#=��C=��A��O1=pM<VVn=�5,=��ٺ��=!s?����;�y`=백<��d���<�xq��&=\T�U�<x*�<�*M=�w�<�z��"��;�4�Qy��*=[�=��d<��#����=�r��t�L=V�9��8=/�<8=�¾;0<��<�(�3,Q=�_x=h�H<��Z=R��;��jh=C%��򎵼��z<�h-=]:<�N"���GB=�j�n���
�-=n� =1�
��>�(���=%��6���^8=�7�e�ɼ��o�� �<��=\L��r�<�����i ����*���Z;�t/�)B�<����i-<׾��<9P�钹�'O?�v9I�lf<e�,����LX�Ճp=p��<Eh=踟<T�=��;���DBw<�wH��$?=�oq;{�<j*z��M;&�	��ؼ�/=��<�n|���u���q<��<ژ>��Sżk���iU�<Җ	=��c��7%=}g3=5#n���,=
�?p|��ǟ��͉;u�=&�K���x<rj<�AL���z�<[[���N=���c7"=�\��9 �<��P=g_.=v�YZR��q���%��RG�8�^<p��<�U�=�^S��i�<�k�7�G�hCi=�R���UI�5��?!e�)>n�8�)=���<S=_��<um<0��:t
x=��b�y�<���<�ٿ�S�L��o=+ =@�<n��<N�<�O���=Tl�<��4=X�׼v�'�UN�ӱ=&Z �k�l<�.0=B����;��U��(a=��;�/l����<O⼵<Y=����k���b=��w�ȃ�;~�B=B���)[�<���<��l=� ��r��<l���h���=/���=4�`��0�&iq���=*�.=񧢼��</�mT��..��#3�v���m<^K:Dr1���T=�F���<�};|�z�o����-<��W�Z�pk�xh*�8 L<�1�=L�<�}���A�;.�׼��D=��o<wYo���z=b[!���.;|�<E��;+� ����c�/=xM�<��Y;�y��)=qE=����򫻪x,=G=�x,=(
�;�0����<���� :<Y;�<�% ��`G��@=/�ϻ��_���-=�������LH=��j=�<^�Ѽ	�����d=Rڤ��=�����w*� R���L��\9�s�	=
_�;�9T=ۡ�<�*=�g=k�t��%]�����%�R��b[=�/�<�}|�N�x<�y��#���|4���<�=ON�gm�	0��(V�\t8=��׼�+��W��
�<���<�ϼB��<�<R�=㱅�Q�<K�h��z�c���{&<��Ӽ����l1=���=�����~��v��Fm5��`�;�%6��"���M�F0�;s9=8c<���A8ӻ �n;%5=�bw��V=� ��7�I�W=`!L�L�=�r=��<~LM��Ǔ������=�ݻN}=�^D<Lȧ<7�蹁��<6c=SY=bJ�~w<ٱ<��:=:�O<�Y��)���;=��2=���<�SW={�C<%�>���8<�A)=�.J�f|���=�i��+<*�T<��=�=�f��Ɖ��݅=������N[�1^=��;o6�<r3s<�x�<����m����ʼ<9�d��="�����G 7=5�=LH�<��'=��E=�a%�0~}=�T�<��5��.����j=��V�'�?=�	4=��>>�:)�;����#ż�M=I�=O¥��1�"ͫ�����;d����)2���]=1�l�"D3<�G9�Օ*=6�<�֦�Z���x=y����4�������O�L����=�Z/=��G��"=�x�<Y�:��	�8�<�W��:�6�F=�ڼI<�d<��޻d =G�ݺ�%C��;�;�v2<>�I=��=�^�Nfe���+<�(v=��N�:��=h�O<�~=��N=X���Qmg=���]3)=���=j���6�����<67��q��k�d�%�R�=?(�-���T�0=;[�t�L=�m=�a��&�<��g��t_=��T�Q�=�2�;�໓_	=��:�`��"�<���<�������ʺ�o5�3�=��<��;�S=%�a�� U����<��B<�^���b���=�:3��7=���<H�f=3\�՝2=��G=ؔ��E�;#:^=�"=�Ȁ��
��R�<;,m�Z�� �O<C��<��x=Ьy�_f]�Y3��,�^�3S��C���0�<?�o==�A�g��;��(=X{L�1���7p=p ��U�N��?/�r�
�{�=�>�<�A5={pҼ)O���A�Ν߼S�ʼ��@=J���+�J=a��+���<=�A�]y\�1z-��#���?�<���cq��|�Y�h�=��ۼ������>=��� �a����a��y��Y.���缞���F#=�}�<�H�<��<	�<%�b�d�e=?`�=�O�*mJ�Y0=��-=orͼ����#��;)2~���*=��$=~~���D¼t�3��N�!�����;�E�<3]S=p��27b� �M=�rv=��<+ӧ<�JH�29=Yd�=�tR����<�=xE�<��U�#)=�Id=h�j���A=���gbD=�۟<��}=>U=�ؼWsd�B>��KǺ<��<	�=��O�i�V�W��t�;��;������Lz<f��l�\��,A��6��~uI�iJi<�����i=T^>�0��������)=]�̻�(�=aC=�c=�־:�
s�Ǣ�Ǟ��eW�<����� ����:�Ң9Whi��1=�ω��x��v�<u�'�C=[r���Ҽ<d����>�;a.��b�������D�}<8/a<=���.�<��� n;x�ϼ�3��sv��m8�T
i�$�R�>J+<I@�:Z�_�1;�� �[����/�<g���d8���E�U?==��n��@ݻ��}k��7$=&�}<}��<<�D=B[9��@�;���{|b�'l=Z���7WU<d����[=��=��(<]mg<�) =G>=����$��E�/G��/h�<9*=�^�;�y��=�=V�>	��Z�<.h=�j������<�$,=A����l����ƻ�}�<r�>׀=�ݍ<��;�Ȼ��<e�*��?μ��=�мm�=�H=>�=ޣY<��'���W�i�����6�qU=�%F�}PW=��N=�1�<��^=ի=�����ြ��)=�M^<>��'=�((�|�i�*
=Œ�O�ϼ��{=�o�<�Y��C�2=�V<��S�G=f<m�#<?�<"*=�0���<�H����<�o^���ӼZd��6�N=mNP����<�Q�<������\=c�<����6�<"��<��8���r��8�<{�@=��*�<���^�<��~�� �<��K����屮 @��so��_����;u��;h��p�������c���<���j(=��;l�@�g=T���Bf�.�c�zG<�����0<:E ��{�;lY=�IC��]<=�W��H=V��9�3��8g=�߼'*=�-��9W�+*��=?�����<1�=��R�� ]��E�<�ml�%�G��[�<|$)=�XC���4����<k��<�7L=E=����5H=4�D=�|<}�]��	E��P��	<3G�<���<���<`(C<CR�<}���e�R�<<�� ����U	�=�5�gK'=�=�9���g����_���o<�'e�&C<+xм�o�<7���#�+���%�n;���f���J�ƣ<\�/�k�����<F�ƺ_l���ǻ+ϲ<��=\z��g=���<)j�;�݋�;�$�V���g��c�V<J�<0E1�3�� ^<��<�1=�-ٻ�>�<�X}���2�����Ym����m�N=�ż��F=�/���H3=8]<=��f�u=��<�xռz	�k�';���,���H�<��=���=|P��t��<�&\=�x{=��;B �=��e�p=���<�ae���<�cc=J=�(�<�m�;M��<�Y=��=��=�5ݼo2N�3��<�oY���l�J�����2<a_c�
P�;hMU���V�)��<\F=�l���S�=����c>�"h
=J,���l=qF=�&��s=�:;=�J��-H<=��ۼi9=;Z�<�
���^<ϊ�=J=�ô<�Y�;��,�us��8�<��=IU]�qc.����;��޼X.H�]��<3��~"!��B�<�U.�]��<]���}
<=)��	b�n��<��y<�&���e<�-[<��F=S�U=�ؖ<��;�y?=�fr��A6=�:y<R��A�&�i�B����<K	���O����,��[E�U��T�<W�S;.V^���f����;�£�W��<�%�v�<��H��s�-> �0F�,�ػ�E=��ü8�g�<��<�
)=�����d&=�l��e�=��2=%,��鼻�uH�X�E�X�*=j�\<Z��-=(����냿�L��yh�<}��;���ҟf�0�<��=<�	�<7c=4��<�V����/&6=�#�<��9�}�4p=[����]Z=�{Q�˚	�OՓ<��	�9C=��?<܈9=.�<lT�<d֓<c54=�`м���:���<Kϯ<!�=Xl;=�N��EQѼ���! �X"�<�晻���ڴn��=�����ټa�:y����<�~��7�.��<S8V=T�9=T�'�_o�����p�=��,=m��<�o7�
L0<�BZ�J�ɼ4`�<v��;��*<nd)=ڟ\=��<2ɟ�k�R=LoE�%�.=s=�c���鼾>�<��=ZB<�V�J�8=0�C����cN<��\�t@�����1�� ��~��J �i�r=�/#<�b��sp�<5v��4=/�!�)��R+�LW�򸆼�U8=ol1�fa��������ۼ ��<���;�@���Ӽ�f�<L��;���Tq���B�� [<e6<@*�3y/=y4;��"�� �<�o6���7�YC=�jJ=@n��a!��V�B=Hβ<�a�U��-��;I�w���P<�z���d��8�1��:P�U��wƼ�؀=�J=(a5�L��;��=�=o���L_;���(=��:n�r���������/��h�<�I��A��<_j8oՊ�=�Մ��X��A\=gL��&Y<B(<�� =-�k�R��<��=U��<�xҼx6�<���;d+���'l:�>�=Q�G�
���68�Z�.=xg=)�_�ҩ�<%�"=��f�2CW;\Yļ8��F�X9ػ�9n=柤�u��=�1�q����g���<�g���V���=3�O�H;ك\;��= iK<���;DyѼ[_�՛;�DH��^���c�OT9��Q�����:��Y$��-�=��n}@;od�;��U����<5���.Q]</0V=2#$�b��<4@����Ἵ�	=�`�<I�=C���B�;լX��[<�vι��¼�	лQ֣<�Ұ<;��ʨ�$�=�'=ՙ&=�**<�������;dI�<����T��Ĺ��o��(��	�`��<.�X$a��߃���=�Y4�V�w�X��<u#�<�g�M\���h���|��<5W6�&W}��.=5�=6"���xU=R=��,0.��<=��
<�i�c�X����<hh=m��E��U�f0=�����=��=��R=��;����s:l=��'�0(��w�����<:�#�2�<��P<q��t
��U��)���K:G8= |���%�{@�K@T=D�r:�4�:V�<�?��[����7��:�����!&�y.�;��<�$R����;�"���!���N�n���j��<�Z<=��"=�E��Mv=�	a���Z�:���p��;��V=)��<��<ӛ������G��n/�<��t�9j:=-�=a ��k0i<�� �y=��e��r;n_B=��<-�
=�!�6�7=nq���	<PO�<#:"E1�L��<��?`_��/L=�5�;C���+=�=���[O���y�����r+��8�����<E���{oD==���"�<8|_=/��'�3=��H<K(=2��J�e=lF3���<�ͺ��(�<�%�b#G�h��G#y���M=Ə���ɸ:��IZ�TQ�j>=�\=p݄�kb|<�l:{��<�M滑'/=��=�9=��L�g�=�#����<b6��]=+�S�~����m�7��Sk�;��=��=��=�D�<>_���=�寮F[���=���t=���<Sħ��q�;�c,��B=��8���=�C�<�@ =�?R="�=*�<�40=�Ƽbk:\��<jP<���5=;Bs��6=t9�<&=�=[���M=I8黚J�;��8=�ֻQ`�p�7<7e ���M���+�ae���&J=��v�t�<����,�;�"8�^�<{K7=�W���?=.
���zf=��;=�z1=���<L���=��&E��#�d�=�M=�Et��Ƽ(S7=�4=�@ �u�'=�9M�W��<���<;�S����?�=<� =��<�=OE��<��<�|$�I�e�'E��Ԛ=(}�<&m�=�M�<Z�A=�*<��<Fx=�nm��Ei=Ӵ=�̺��ᢽ�Y=�@<"����\<�'�2$'���ڻ�=P������<��a��-e=iX<lk��a�;X��^t����<�ӫ<��a����;_w�z�;�<d?`���^=�~;	_��(<j�,�7xD��c=�&=h�A�J�Y���ֿa=k�<=�!O=<�����D<"^h�3�=�<�W�<��(��(
=�'U<�!��''=�<V�P�=��H������	��;��<�*,�g'=3T�M�Q�%�$�R�1 l��������;U���)�J�,=gS�<�+W�[�!=ȴ�<���=��V=��6�Ｌ� �O��K̯<��<���<���;~ܼjb=��>=�}��xj=�T=xE5=*�q��Y�J��ļY����=��<j	��Ǽu�L��<T<�fd<�*�<������Sq�<�<,=_p�<��;�?��3 �bs<�0��)=sy=j4=RwS�u�u;�m�<�;|� ����<���<5A��;��G�ma�<o$�w�#=H��Z5S<O`=����3�8=����\�i�&ռ�n;�T�O���׻=�=���<pq=xKc��<�糧4N=���<n�8��ě��1��\��}��d��&��;lyü�Z���<�ό<^H�</)�(�A���<9�I=n==<�=\l4�{�<CA���:�=�=A�;�WR<Lv�<ǿ�=Hm=��o=�;W:�=Z���J=z�p=Z�<�N>=E�:�{Y���g��w�n�R<�#W�C�	<?8><��
=S!��=U	=����Ra;��:b!=��<���<�X�<�QV=_ ��G=� =q^��d=���;B����-==ڄO=�6�=*=�uP�����H���l�.�Ѽ���<h�T=����;�:��<H<=f�S=����n���k�����;`<b��00���
=�=Gc�)�m=�fq��<�aJ;���:j��<4U�<Cw=Z��CI=^�<_��/��[�W<1W���=�0�:���;�(�<��(��>=��!=$��<�?���F��H��<֞�5A���t=ԋ<�Y@��;����w��m�P=@I�=Ѡe=��=�+��9<%��2�<,tƼI�D=�a�GxK��;�e��<�����(=`X�=��<=|H���<��=FN�ޚ =�������+C���6����<bв<��Y=�� =���Lԋ�S���)w;e��<��V=��~=/=Z��v��<��O�Wf
�?�ǻ[~*<���ۗ=�s�<�b��P��W�;�N$�%N;��)=+n=��"��/ =�X��7n=v��l;U<��+�5��<�=�s�E;�!�=��/�.��H4�;�IR�8���輇�G=�Z���`㼒��ҼL=%0���<��ڼ��+�����<1L�_�{��O?=/?='6üԹ+���<��<<�=�<=��f��?���=���<A/J���4=)N�P�kX=��m���"��"м��1<o�=���*)a���F��{<:�$=�廚�=rh�X�
=��Z�ڥ<�c�d�P=ȏ�<s�?<Fl�=¥=��c=Jļ�!=�B�HS�;��-�񏵼�BJ<�;�\!=d�E=J0<�X��{�o;�S@=�q=���<7����2=�O����� ܸ����<o�H=\���^�f��;x�	�{�[��M@��ښ;��"=�=���-�<9���E��3��Pt�;�ǿ< P�;�f�<��<;�j<���12;���<k#���k=B[�;����,����<�p���=5=~�5<쓈<�Wo�5h%=Lw�H��O<�<�._=��c��V<��$=/>=�%����;��;7]����<�\=�K=>m<�N<��j���1����� (���[��Z(=6!�m9#=���;oB�f�<�`�;<d�&<�'���o=%縼�"n�A`%�罚���ݼ�X=�\J=:��HO��E�Ҽrj&=t�l=j<��8 �	F =N!7=S�A=؄�;gD=+�V�s�7��y_�f�B���@<V�=��;:=��DC3�%�3�8%Q=�3 <�L?<VkE�]>u=տ�<�<8�<'-�<^L/��a	=�Ad=�l�\�
=�υ<��<�F�<��ڼ��]=��<�=����~�0�<�<���<�s�ME=�dh=F[��C%=Sqv< ����� �D=ޢ�j�<J��<�5���r���}<�2���f����Q=�m�w6m��U�<�?�R����(�ڱ��=&=�gb=�q�<�
�<��H�G�2=�k=�]��^�<v��<�I=O�d�J��<�}}<�_l�|cE���y�>6�<�YI=�W��C�='��=b =^D���p�<{�[�C<��=���P=��	�2��;���<�,�p�2=�8#�L0=_�N=�#b<��s�>�޼Ҍ����< �S=?$h=��μ��<|u=��nt2=�1	�tCY=�Z*�k�1�.�f�w��k=�6=���S�<���.C�<<w_�ʡ7=Aϥ����<�x7=��7��YZ=�5<�ή;�@(<��(��7'�^����o=�j�:RI=p�W��n=�OG����,f�����G�	=7��d<i@��M-=F�<(�E�G�G9��m�Jb��] �c=��1�-�E�i\��뼐�*��zN�w�E=U8弢:����� ��<�T=V���&:��6U���Z�>H^=�'�����'R=�[��G3M=�<hx\= T)�����Nh�+�-=�X��S-����� ����M$��5N=��<��=��_;;d=�P��т���j=8-=.��<ײ^=W�E��;OR6<^O=2����;��=��;=�T7=\0s<I�<�"= t�<��=) �t��<(���X�05Q=R��3�#�f���<�<p=a�Y=�s������Ok��3���=�|�X��9G=�X�<�
=���g!=�ؓ<�Rg=��L��=�Yx�i�<:�s=c�� �v�C���ϼ��N�f�D<�����|�<N�<�Cx�c=Zw�N�=)��<�ά=�Vu���2����=91=!/5�~R��d�w�Y�b={�M����;�eo<	�KF]=��*<�7�P��hr;���<��j<QZ����[�ʾ$�� ����T��<y�F;��<�a�<�MK�汞�ț��.�4
����^��~y<�-�<��<�s=x7=_u�i��<�=��a=^n7����u�	<��=��<k�{
�<��O�YF�<kļ�ST=&=�<
*}��D���$=�S�<�9V=I�,�<�����
�<M�V=�ϟ<�&�h���cf�Y^�G����:y���<�F=1��;��z�	
�<�����.�e�:��)=�r���(���:<�'���#�o@v�d�h�[QG�K)�;�N�<�=�ݼ.�����K=�o�<�ɻ�p9K���$<I�<!�^=��'<ɞѼ�wX=0��A)�<s]Y�Q()=�m���W�<t�b<�u�����<�:X=J�E=o�=�:D=Ձ��h����\= B=���<̿@�I'H�c�=���<�Ӽ��)=}�f<#�-=L|�{�"=T��<���ٜ��f��4�B=����Fs=���<����*�g=� ��8<M
��R��<��J<O�9(6�9#��;�,<e����:����<�"=.2U��
K=O(<)j��ɼ�J0=�.�����(=,9�����$=|��8���w(���� �ӣ=)@�D	�<��u=�A;�?�d=��=.d=]����<q��<'��9�7���m�F�S=8,�<~�ü��7��Qv<*jr�p�Y<MzI=2\�<�˘��m%���ƻ��<��<Q�˻��g��Y:'�?��q���q=��$==��S��V�X�f�`=8�3=#�#���?=�[)�x!D���+�m��<g�N:g�}�c�(=��z=6ͨ<��<ٳ]�\���I�;��4=c����&;ٿ��:5�Н����v=�ʰ�Mި���<M�4=���<��ռ��	=�n*�e�@�$m<�tn�)�Q=��<��(\=�}�};<I�<.=c��<~��<K�I���<K�=G)�<*�4=�=~�|������m����;�;;�xA=��޺��=O��;T��;A�=�5���:��<�Q<Y��;�ȉ<Y�<�2=.�=��'��t;�g�<���>=����<� �<ҿ[�Hh���G<&��	ou���\�3=9< �9�u�	�Fy�<__���q���"��˱<->==��<P�<��^���lgW���;��\�U�����;z��<���;�+)=�vS<��<��D��,=��
���2=�
����/�S�=s��<���<�0�0_=��ͼ��<����;�w=U@<f����)=V��,Z+�ęW�����w:�rI�4�<^�<�+3;�c��p<0�s=�<��@���<O5c=��F����<?L��%M<3i޼(k��o</ּUn.=�<d=������:
i�;빫<&g�<k&ؼ��W�!ԣ�5����<���w=<jw�B9]:����GUX���=O����'R��TP�lI缪 	<?,<㓇�0���R�Ҽ�ݼM�'���]����%]_��F+=���E[;=�x���g4<͏2��]�	�=2'����1�˼��Ǧ&���V=�
�������W#��@�(�<���<+ޕ���2�}��:�<�Լ2�e���!=��$�e�˼���/�?�)$'=�q̺|�=�Q=s�l��pʼCuQ�3���(\��׼sY��==�/=��J<n=�y����<�&=���<�야�I�!]���&U=1��='�1=�f=��<��n����/�<9̰;�І<^�<� e�TF��S��Wy�<'�<b��<� <Z4<�P&<<�B��|G��-=1%��'�Gt,=.�A=�R=� <x_
�����Z����ek<���<��a� jI=�/p=Dq<����s=}~��=j<R�<��+��3�\8���D=P%=�y������E[�"�>�I��:�=��<VZ伹օ��=��Q=]~�<�B)=�.�;kyI�{�>��3u=r����=��={R���W��M\�o_�:)@<BxN=�ea�_!L���-����;���;>9ѻ��<��;�O�]�A=��h�?j�ƿ�&�g=2h=�+V=�y��9~<O��;l��a���F�<��K=P�"=#uV��+�@eG��zԼX0ӼڗJ=�T#;
 9�s+��L����<'fl=�1<�I�;��j�ɼ>�<�5�<Җ=L8=�2z�2EM<�<���<�rn�U@=��RU�����;5���R��nz�d�d����I1�<�|�:�&�:n�m=�w<m��<��D<9 滟de=ŷ¼�$<v�
=�$=Rⶼ?}v=ZQ!=�4�<1+5=�YD=��m���<��4=H�F�`'��O�<YR;dvM���N��l;V�=S�o�=�M������=-�j�$����ڶ<��af�����׈�<�R��yMO=��]L�~f<�j�<�<X�Ys=�M�`o:_m:�6@=��L� L�ji�:F�O=�μۅA<�~�<�;�6���L�<�\�RHV��E�v=��:�W=2n1�G/F=�"=�� �=�_<��=�t����C����<x�û}��-J�;�{Ӽ�6�;����|ۻ�}�<u�Z=���;�L�"��<k��<`(�;~�ļ~�~��F4���=ތu=��j=B'W=L;3���t�
a�2B:=��`LW�?<r=Ƃ�<�����_�f��<�^:U�v=Y� =׋<��	=�T!�mJ�<������<��F<N-��SP��8<��k�'�z=���<�^�<˽m=~�̼H��_�c�7��;�;=�m���c��=��i�K�=~Jw:`��;Q^��v���+��.��o����=<��!�Z��<۸;<�7�q{=^ڒ���<
x�=���v	��?�]~�<��=e��4�;=+�	�#��Ab��
mg=���K_�(7�)~Y���h�S[�p�%<l��<Bq$���g<��$����o9j=_�'��	t=O' �X7Z<��޺��%��<qY=֎;ژ3=���F��:@�f=�3U�˛��B�ɥb�c��3=䨼r�<f�g��QO�ݧ9=;�)�q�<�Mc<���<��4����<���}0�����仼���2#S�j��<. <�ث;��;�!�<a��<�MF�������\�#<k��� N�T����< �<�5=ܨ�T*��"%ռ�`$=�);[��/]�<�J=�>B�g�C�I53�@�j<�{�<5v<�A��R ?</�<U^��U�;3)=�x�VB==7�"�b�u��Xd��Δ�A%���il��c;β=��6=� 漅�S=�/�<��,���ü�(O<_� <���<=2�:��GQ�;;=E=Ț�=5y0=�2�<e=�'���;���<?uZ<k�@��u�;�<n�<9�X=���Ԯۼg��<i޼5i=Bt���/J</L?�L�f=��1��7㻈gS�~W�;��Q=[�d=M�m=3<�<h����@=
����;aZX=G3�8���(��~{,�K�*��H+�h�'��10���=0.�<��<��@����<9H»�4=@���E�Q<c�2=���5�߼�y�;o�*��sH�;4Z={ka���H�'��E�bs��[=�<_<��x<��O�����Xx�����DR��S�FR=d,�^�r�g�޼n������V<p��<CX(<��>�M�L�|#B=!�=��0=�x=��%��.N=���<�T���C�<Օ����<�Q�=A�<�y��P��<��A=|^=v8�z�=��_�/�ݼ'L����C=k��6��5P�<19Q<it/�f2K=�#�m
\=�.<�`@�	�i�y3�<�� �Z8=��<B
 ;���;��=���+��=�yb�0~7<��8���H����w�m��B�B=S�=�ZW;��^���V=o��%�0��<�y=������<��d=E�
�d9Q�0M�`ؼG�b@Լ�[<$��;T��=���R蛻���-4�;Si��u�/��W���Ƽ��</w�<?$=�70����k��<ܪ����=�1�;L�t=�ӑ���99={�;r��TI{�n8����:�t� !��/=9�9�	�1����>;<�	=�7�=�b;��O��7�����J)��Pq=�Z(=B�����7)� =�Af�t~3���a=�%;=J�*=pC�<�4&�?�=��=����|>;�������ͼ�hѼ�K���	�=��\�K=�Am�y���"$�%�!<ǐV=�W
=�`T=��2�u��^3=��&��bf:Y�<Y �̭�<1U�;�/�;�)<3V��m�Լ�CY�0+1<l˼�)=[N�<�+��D;M�=�b;|O=���<y|-=c�M��� �7)=�b*��"��j��,��H=C"P=�@%=�i��ۤ���
�	
<�B�V>��P�����e�
<�x#�
~D=�%=��r�� F<����^C�}�y��?<D�g�ݻ0Se=�Y�<��<=$=1P{=ղ̼�y�t�"=kW<��=3Mb��w=��q�=��<HB��л[}\<,��x�;<��;�&� =A
���6�ʴ<}S�<)7�P�)j<��0=��v��¼>&V�ظm<>c�;k�Ȼk�><� �<˖��
�����<6J��`(<�JO��<I=��*�Y�<"��<,�$��k��U,��ɸ���������|1�{l�ʇ��M�<s��<2�m;�����[<�����0=��<�Q�j��<2���+�<�`D�� �;��)�jD��R�z<><�hl<R��`)�B�#���Ѻ��=�i��O=V}=Z=������;�&����<� ��	��:�G=�.=/1[���#����=%*����K��G�<�!�<�p4=C3�=�� =�;jm���)=�Aռ��7����^y�<MU�:��8=*'����2=t����z�=��<��*��ex<*5d�|�<�=�+���~<��߻b8��|�:bL�<���;�^t�\-��*�x���;;:���yj�u�=�0���a�]��<��� sj��j�<{<!6��=�����<�<����<�D���t�	�3=�4�BOf=����dmQ=��r�]�������4��n����k�?ȼ#.=��<�Ё=x�%�D�<�.w=�Ի�Y%;Ĩu�/G�;�h缊r�|��<���(G��%�cGU��F�#X:��9<p��<k�?=��k�B�Y�u�����9=�v7���W�{F ���#=}���s�����>��;�o���\]$<4:p<��3<��\<�B^=�k=�7 =�/=��z==���o��߆)��ms=t��<P�L:��y;7՝�C�C�uO'=�*��{���3���=*�<�x��g�D<�5<�����0=#{Q=d�ټEis=�V=����W�H�μ����<S�=��<�&>=����G�;O<m�d�R7[=[0a���6<q[a<=����'=��˻�xP� g��Mg���<Rt�;2I^����=�u�E\����63�����<Ė�<g�[�,��<�/=�4��;"=�c��Dq1<-��;<�3���<8��p�<�Y'�;�[=�pP<�.�;���;�u ����<|��<�����=��=g���>�1�V�i=��=z�<n�A���ؼ���<V�=�#K=�Ρ�ԭN<�i�bH�;rz�<���zԸ���b�e9H�T=�漓�k;�ɥ<�T����伳��\�<����z�h���'[�� <�u���7�꤬;�K9�Ɋ5<>�<�D�OqN�4p�]=籁��i~�Ι"�K���T켉kX��kL��%S���<9m=�b�=m�����"�X�W�����<@�n<=�_���<T\�<�Xj<�:=�#=��Ƽ��1�W�4��oһ��9�缯����V �:�����<@���d=\��zr=E�=���#��B=S�=�WN=4�T�����U=L�v=<5��q��<B=��(=T����t<����)��h�<�����������<�^U��[�ܛi��J�T���=s9ͼ[�<O�R=���~�<�@<[Z�����R<aM�%"κ�R�Q޼H��<z!��>�F5�=�#�<�����Լ��ۻ� ��߯�<DL={u�����u���J�<�DH=�p��􆼙x=����-�<�=Uq�:�P]��N>=�;.���;��E<YKg<��h[�<{A���� ��N=i� �=J��Ȼ���%T�wc#=��O=X,T����ù&=2,����+=ce<�N�)^�<A��<���;���v`�C����"=���=M}�Q�N׼��N=�޼F==qc�;+J���<�n=u#'�M�^=�-=Z�ռJ��;�/���;�����>ȻmB;���L��J�c���μ�eڼ$��<�^/=7,��,�=�H��L����M�;��$=ݓ#�����H�;�7�����:��};��s=�I=`��)���E�P:��j3C=�ZF�f�1��I=@�#��%����=_���p�<aEc=hj�kх<D����;M��(Y��Y�����E=�^�X�x<��=a-�U��<ݸ	�B+�<��)��՘���R���="~ܻ�>�<�=$<~[���<�B<�-:�=�!�������~�<=�v=���<�z�;0$����;�����=��=V���L6�<�Pr��Ƈ<���PdY=e%-=�� ���<��<W��I�n<t�4�e1 =^P»vz�:f��6*�i��<�+�=c6_<=2=�a�=� =S)�<vq;s�<�q�<=*�
Y2����:��0����X=0=YD��)���g3�<qA�>�»Q�29]�J=��p��.�:s1;^U=����)w��M�<��C=�x<��=E���n�<�8	=�*�qND�.�h=g���8�=^�߼�s�;�0,������H]=(�<맘�Ԅ�G+�D�C�}6��2j������y&<;�=�z�;��<Mq�¿�<V\�<lw���e��\�xr=�Yκ������;Cwջ�E���F=yJ<�<j�6�%z<�����<í�Qﵼǟ�԰�<ڂ=�����	��Ӷ>���0=I3=��x��E���a<�<A��V��Fμat�<i]=a����n �6z�<h=Ɍ�<��
�x=e�X<n�b����<{��%��� M	=-�P<m�<���-�\=�5:=;=�?=�P���R=�3 �w�=�<���<~]=��m�Z=h�:=[���C�ln<�V�}6y���;'�=?a=�TQ<�̳<��!���(=��1�U=����Ҏ��x�9�����Ҽ�t;�w �@�<j-<����zؘ�D:=��9=�)¼L�Լ�p==��R���D�Jc������� �D�U=s��<�M-;�gf��U�:�;=MW�_	�<y-�� ���|}����=<=8�<�',=L>��!�<�J�L�<@|8=�`P={���hݼS�j;U4ܼn��:��<�<=^�w<���#=��A=��I����'
c<St���i���d:���<w>c�?Vd�r;�M����L���<�˳<6ZS=�v�;�A=�J���V�y� =v�l��|�����k=\Yj��P�t�=�*�<:��Fu<�)=q��ĭ�<�E=Ř�<�u�v�i��+=ۄ�<��=C�<z�<O�ѼڛT��}=�>�ˉ���� :�O	��<@&R�#/s�F��=��=�1��v6$=��O=��i=���O�һl'o��`=��;��*�Lc�]�n��j伇)Q=Da�<�o��ژ�;�#��~Q=~��;�[Ȼ�[�=��b:�)���ʼj3=<�<�.G���I�ov=pP������<�:P�*pa����<��V��Qd���i��������S9��� =�<�y<<j�<�l=��<l\,=Dz��!���i={������<=ϼ.��:��N=��N��0)��S��_0<�=����f�-��kI:�N�=�+�<+�;
T(�W@=��;��$=0�6���K=1��<o�����@=20S�ʹ/�B =��Ђ=��<*������y��<u��<El�<����D=�E���<��&��l=!W=v�%�*:<�����i&���c=þ{�U�5��_����:���܉�;����ռa��@�鼙/>=kAP��7=�m�<,�<��4=��#���A��Lμ��<�<�t�����=�B�м�=��R�$�(=#�x<c={�b<������Y=q��<��
="܅�|���S��l��:X >;5�K=���<oe�<5�=�*0���r=GJ�\24<j��<}=���<�o�=D�0=3#	=ϻ=a�=�xż3-��8�<p�L=�f1��,�U��<����%T���1< J>��Eۼ��<_N�1ռ�u\<O-�<�l=[ �=��I�S�	�\������y3a:�2��`P��K��k=s��<J�2��#����Τ<]� =�]�<�K�;��<(�o��x!���c=�q��FQ�!$�<�$=*`n=H��[Z��5=`۪�!�2��b=��L=��T=�2�<e�,�*�&�|n��ke�=s1)��ֈ��9���B���P=u9A=H����ʹr�}��<�������t��<��<�Vq;�;��U"�<�7+�����u�<w�=�XX=����gj��#*�(
<�88=_���_�<yN)�^�n<zX�=�b~���.<��[�/@J<6f�<-M%�4�ۂ'���T=/���< �=��\=����T�=:�=;M�;�:}����<������9{�<9�<L�a�L��<�%=y�&���<���<��z���q<yy<=��<Q=��<O�&����v�ǥ.��t�)q=S8K�O=�Q`���'<�+�<C��oG�<�4�/T���T�H��<pD�;�_�H� =-Bj���{=�"޼��1=g�8;�-���gG=��@��U�<�;�=%Vl=��X���p<��=��B,����[�`��<�8==�>�<[��H��=��9�	��[oM<�;��l���ݻ\����q��=J�#��@= �=��;�R<�a;��9��1��o�<��S�/�<�}��Zg�n�L=� �����ъ�'g=��=��8=0�޼��<[&#���<|O���K�	c=�4*��[0�����;����a=�h=�Jo<m==�cG�@��<3��T���r���n�<��
��8��Y	��ͱ�}I5=�	n���,�y���T�;�Լ���;���<��T� �o<o)�<�QN�ɟB<^Lo��et�9=I�<
���R�S8p=��j=�0�;�E,=�����Í= �&=;�<{��<�U�;`Ǽx)$=6�<&�A;�s'=ܳ��K�HM<�K��Γ<:ۡ�)�<?ȅ<q�;}��97�N��<��;�k<���i��<�����a �0�U�#���{a�h#%=�ߏ�	=�C=$��o圼vtE��ht=�^3��a=^Pϼһ9���V=KM󻋡j=��a���!�B+����'=v�����ͼP�N=1V��V=�l#�o2�=qd�<qg]��_�;6��c��=�Id�g�l�#<�q䶻��&={t<�^�d�q�_=�'�<�}=i"|=�X��)�{�=�e=�7=-}�<貝��~C�& ����C��y�;��D=��;�-=>i=�'ټو�=�<���<������=��<��s<%��;��<�P6�������<��J��؀<bv�<������&�H=`&3=2%����0�1�%=�X= �0�+��<}��b�:[〽��w<��8=p (=��M�~��<s�;Q�����3U �2�=i}(<��¼�r<LRs� �k ��<�v/=�
��ʧ<��<�����]|=4!?��ic=)�"�aD���E:PW,��}\=�_ �%/�<
d=��<"�"=:�;�+��h��,=[y/=�����%=�ǋ�-^�� ;�]�Qo<�żӍH�wT7<�2���O<g�=�;�0��=�������~D==
���=�G�ӓ�</��=�q<�\�<%��̓�t�ݼrH�9Y���@r=�hi���
=q=d ռ�ݻĠd�x�~��Dg�$!�</57=��=��X���`<���n�d�]\�:S�:	N��.�%<͎����<�3)=��g=n��U��;'�N�	9=�)=D�߼�:�����z}<=�;e <��<Нn=*�=I|�"��� |<��P��=iq���N<)Z�<Qҷ��W=W?^�!)�ŀ{<���;�%�<P�<�Q�<TQh�G$�������<gb����<n�=��9=&�Ӽ���<;x��_=�k�*$���� <y�Q=x;�K�G=` (���+���2�2`�E�<��f����:"��'~�*=�T�<{<s4^=Z/=�ˤ��N�AI�: �<;�[=Li$��:K�'�M=�����<���;�G�K���B=��<�$,��+,��u�<��<)h���Ƽq��<�b�,�B;`�c���<oGV=/���h��#C=�J�<��	=(��<���<k�N=N O=�f�;9����=?:��2H�<��ü+����[���yI�9�S���R=����,�ע����T= �==�ە�
05��)����'�<%==�%=��,=���E����3=�ĉ<Ɵ.<ݡ�������<d��!=:DF���e<��2=,���&�����&l�R�u��<�E��WY��3�<0S<�d:U��<V�4<�)�7�<�K�X1���w<����=e��<i?��Wȼ Y��^��<����jԼ��<��O�X_�8.�(=¼�8 �z�\=�T�<,}i<��f=�s8=1-=�&=n�<E�H=��E="@=�9�R|=:�9{������n<��3=�GR=Ҧ���L�!�k���1��*=[q׹�Vl<VD=߄�<b��;�`�;,,=?�A�:�ż<�j��/=E I=R*I�k��<"�ɼ���<F�;Y�g=/�N/�<xp+=��)=�{��Zb1=�}��~�E<|6U���D�H=8�Os����;jl9�S]/<"m[�:���U,�J��^/=B	\���]�P�K=TyԻig=k�d����<�<2ca��0�4��������I=Ύ���rW�2��B�5�04@����.��<�!"=��<�=��ȼ��:<H�=�G=5~�<3�=�Њ=����M�;�I>=�J=�P��3�R= r�;7��<��X=�!J=qj��V�:�<8kw:�8��-=[��IE���cK:�ï��@�ͱ���0<W\�-_�<�W�_ra=
�	:������f=��m<�U]<*��<�=H=_EY=1A<[�*��3<n�B����;�i=j�\�ޓi���>�~�<��)�=� � qI=h�[=#f_�a?=�x<��)n��K�D�V���4������;˹ܼ�萼Ld�<�{���=�5'�=�c��|�=3��9*	.���
=�[[�-�=�LQ�(�$����q�;դi��$=�V/=H^ռk�=
@=��>=`�:�/:=�/<��7��y=�ּϊg��?=�5=�7�O卻�"C�7�Ƽy��:�	��x�<�U�|@�<�1=�[1�;�BW�#|=92�:c����8��J=x�q�A�,�?=��:=�_�Y^$=�{�<+�%�σ�<�� =�sR�\Ղ��Q�<�B������g�3<wp���ً��g��>);:��'=^���c	ڼ�p���I�Nm˼K}�<�2��G)��'=��/=7��Hn|�e���F"=�U=��-���<��=�銼����5�<��༊��;G�X�w��J'=���Br�3�/=�K���x3��o �	I��l�<���<+��<�?�#.5=�<�P����<�+<`�?=|�;Ne*=cU�X�iD�0%=i�>=ԥ+=e�� ���d=�2a���b=;4E=.j6��M���]=�q�;�<⹡<50���<�ͼZ?J������O�t�=Z�_������=�_D��B��[R)=�{b=w�Ǽm3����<��ڼz�N��I��P=���<)����U<_��<���i��<��:��XI�v*u=?�!=5M<��=���+|�Ҽ�<�^=��Ҽ;
L=UT�L7-���<$�p=:I�����:�io���T=8Qq�F������<����=O��1����==�4<���ר��~�<�ļ�G���=7�˻�^R�E_[<��F<4!d;>g�<e����c�<*Z+=���<<�< ��<��/=�؞��jZ���8=�<J\�\Ҫ�� ʼ��,=/�
='�ؼ'�<ݫ=p!O=/�=�zO=��s���B=��;)/1���$��8>�Էy�n5t�7��;\�<�| ���=��8�ɘ������b_�<ME�<��;�?e�ʳ빾���>��ʳC��_���0<(7����`��Z�<WϻXO��n�;���D��g:x�i���<e�W=k�ͼ���c��<$�W�ލ�[��;U׼J����z�Ѭ�<��#�ؿ�<}�S=HGp<'Z=�>��`���~S��f���5��߾�����.�w��<�2�=�����sj�9׭���u<Q���Wk��r.�=����1=�L=XB��BC�:z�<�����<�U�������$=E���w9<8�	���p�>Y�<���=)�3���<y��<W;_<T�����/�9ř<Ţ9="�n��2��0�=�<�_�<�R=B{���.|<�u����<�4=Z�9=ڷ��h4��2�;���.�H���>����<" <����HT=FRE�s�<�����^8�U���=�4����Ƽ}ϼK��`UȻk�K ��A�#��9�f�v�;=t�<�]�=�j�;ke��MK=�s��1�<�C����A=Y��x�<A���S�''��ё%�|��]<w�
=O��� 4*�}�;t1-=橠�� ���5<�:m=�:v=w�{��KȺ��^=Q"H=$�ȼܖ� �r=��=A2�::�����<�L.���=YG��ͼ���Eo��c=��d=��?�-���_^=g�:���'���<�e�<�<ql���=k2'��E&<o�
�G=��=���N�����ʼIL=Mڛ�"A��7<�=��b<Y��<w7 =L�(�E��;��<3缏���	=|�X���P<�U���U���7��N��S��==2��<RP	=t�~<.*��� ��W=�t�<w�G=�J�<ى�=���<�T=Uo��A�8=�:������2#���b��V=���pz�����<�8=�f��h�<�9<yǼ�G=�)f�6�R�ƛ.=,<ۼG���]M��]=�9��1Z�yͻ1X{�������O=0B=�O���J����P=U~ ��Z���<j��Q��Y�<d&ʼ��<���<��<[�Ѽ�l����<C	}�� =�<vm�=ּX�>�E�4��ȟ=n�<A�;������6=Q ��^=��=��H=8�R�m�!=ű�S��=(Ӽ���Ï<�M���;F=B ^<�#|��ɼ��k�h���KI=��ɻEh<c�}<ٯ�<�/=��#�R��<-�o�q�:��P=��s<���<k�=5�)��̚<��e��P=^=����t���h=��<��f�<b���׉<�zx=+r@=}N�:K҆<
*�<i�����<=H'u��|�<�!=<�g���"=|�޼��<�@=[|���o�����<ֹ��Ѝ<�E��� =���QѼݔ��6�:3K&:�o���>��>�<�햽�V=p�u=I		����;}٬<�*�<�i��Z:N��y�; 7\���=[��=DqW�@��<B=����qS׼}k;�Y��<������p��&=�T�����R=5KW���������=|X�<Gʂ=p�_������<�ʔ����D�<9Z=��[�p�J��~��ߙ*��I=���<̛�� �i=»h�u�g�`]C<�I�)�;�1=Fj�<B%7�߉L��n_=-�<u��	Jj��N����<8bz�<���J=��j�?ƻK
<^Z�<�˼z{w<ڱ0�|�[<��<�< =�;�f�����< 3N�qP�AE��J��<V\H<noS=$0@����<í+�1��<L�U=a�<5����O�M�=��<Vʇ�6�8���ռ���<9�[��7<)�,���?�I=�;�X�
��6j�<Y*��1x��s�b<D}�	�=w��M�L<�'��Z��aZ=6����>�<G�z<?E�&[?=L/=��=�O��@��n;=r<׼$Ea<�A�<֠��!�ȼ�>=����~�O=>7�EA�:�)���=���9S��<lAV���?<^��
=c�<f�<�=ꡭ<ofq=�p��p2�q��MKc;j��q�=V�;�U;Of�Y�<:���ջ���<���<xT��T������*
.<�Hb<G�R�(����_�A=)?���S;�o��=�k=���<�}a<�nL=�/�tŉ<��R��=T��<��A=X{���/�<0V8=��<��VR�<e���� ��#�������X=�}?=f_r=["�;T =�<�/=٩��4F=J�J��)3=�����W<6j<:�<uB=�ч<�vX��˼���<1Ъ���.<LE�<عf=.�2�V߼��=�综P4�L��<����><��̼NM;���<�Y�<�d=�Q�=ҿ(=��t=��G�g �4��u�%=y�<=�3���	=��t�p��;#�H����u�k�̓�<��L<�5����=�PG<��;<U�����غ�w<���;��;�f�;Umt<c�м�CN�Y
��4;3&_=��m;�+�pҟ��e�=՗ ��-������s���~����d�6��<����=FR/<��(=��<�	o=��=P�f<���9��:���4�?��P=RQ�#��<��:>�c��C*=Q�=��~<�.<���;8)̻��Q<�%a�!2�S[�H���[����_w���G<b-�72(=��=����	<V���ֻ�le�%����#�<;��e&�zT����E�vȺ�
��<�y�Jݺ=�=P��&X�<9;��^=��V;��<�(ݼ+����|1�Կ<�A����`�/��<ݖ�<��Ժ'�=Z=4��6^4=��)<���l��<O�u=(���T=��(=�q=x�<�RC�)��<�;���
�;@�'=�ZI��=��I�!X�<�
��"ݼ��i=ȲM�f�Ƽ-I���-[���=o�#=����(�׼�%;�΄��#�ʹ»�-�;�e�<����.Y<^��� �=[6�;Ejb� �6�<�D��_=;�~��1�;�<pP�;��=<P&=탲<?"�	�<��h��ϼ�{�;�\<���;�s���)=Lo�;����绻�}f�	�-��d_=��껡�;,�r�d��}H=Ev1;�}%;�"��P8�:f=y�;�{f#��l�<bc��� =^����LA��.U���)=m4=�4�<���;�鐻���<(v��n��%=2�1�2��<$��;�H�<EM���P�C0��RW!���N�Y�<A�����<�E=�AǶԭ$<��%=��<�=;[=��;�V��l���=���<�q��$� ���=�s�'�n��2J=+*P�~�9���D�\;A	=@:�;���<�3��y�==���7B̼�)=�}�=6��<�T�;��,=���΁= �>��U=��3=|
<�{����<|�I=��ݼ�D�;�/μ�ȻX�)������b��C$=��<=(1B�s�;�g:z�=�R��Z|�A��<T0��0�q=|��/�Լ�]0�?���/�-���O=.�1<�ۼ%T�c�m=u<Լ�cҼޯ��(=�'a��B8 �ļ���<p�6�S�<R4I�F��X@�;Y#;�ڳ���YI��⥼+��<q���3!=�� =�hѺU��9,�����l�o���e�U>*�ʭ�Qj�<;f��#%��Z�W]a<T=�Nһޱ�<�K@=�=	S7���8�S�<��#=ϳ!<��=�{<��<K2<�&��E�=vu��a��l�����=N��;m�C�w`e�o=���<&��7��<�C�����?�;;?<�[�<JIC�P�B��<\U��9���<��=�d$��V7�)5�;�=�Z�<�>�<�;���Y#=T��*ۼ�h��K����껊dv�2�:�� ���%���u�`�༛&=�6 {<��f<�&���I='�A=�V�ȓy<���eF�;��H�3�P=ƞ@���F=�UҼ�L�=E��U=���������s=3{"=T���%va��u�����Y$�A0T��&��g�@��G��1_�2�S<�\��Tv3�N�=�"�=6=.{(��~\=�ʌ�)䱼���ï��D-�Ѐ#=�7<4p�<{�� ���Ө<�2:�����pN=fH
=q�c��K�<�=S��<Ui;�:���Ǽʹ=��>}���6s?=�.L�30�Zt� ��X\��w0�vk(<�h)<��'M�����B<�$�u<����Z�\=��<�.=i�=��=[͌<�Z,��ӆ=a��j=�9�H}<V	D�P��;�ɲ��$J=;Q�<S�d�Ѽ��=tnG�`T�<���<Ⱥ��9�=��i�{�-���P<�E4��3ϼ��A=Ը��<�q=>w"�����׈0=@�t�GT;��p<Ӟ��R�<A�\=;.�<��Q�m7:�������w#�����<o�Լ�q�_�<����-���<��[=M��S�m��g4�8=���<�ܻuO�;�eW<;-=����3<+=�<�kY=�� ;�.�x�5=��:���.=uۼQY���ϼ@FK��y.��L�5��<6��RBK<�`�����T���̻tj=5z�Ώ�<\�v</zS�������&x�<��N���\=���;�w	��w==rK�p��<�7�;�,ỾzD����<��x�gI�;�l�h�_;n%Ļu���A���=�S=�x<B]��j]=&s�8;x�<=R��<,�:��v�J$<8O��K=	P��f�f�h��;*�M�i�_�i�x�c�м_�O=�1�]v=r�*1�;T��~=�g��c�T�4��#���<=��	�t�I�A �L�O=!;x��M�<šS����lM���.=��ļ?2�<�<��E�V��U(�n�R����"�Vq�<�y���A��*6����;S��<����M�5�����;��μ��伻��<H���C�9<1���~ʼܖT<25���A�<���<%�R=LkL��G켁^z<��� ��p5�=�)�<��G���%=�� :8YE<r"D=5*N����	�I=fi<��ټA����L<�	�=��{�=�e�<1rR=,8�<%�������M�M~��rs��SI��ڼ��8�U����;����=J-��ƻ��L����<�͏<���DR<�B(=y3=�����U�I+=f�:=zL��<5*���<}t<��@=�2=�i(:_m���;_�;!��;��1=Q1�] �<^��"u=Mt���z�mF;bA�;�9��LL����G�u���q=/��=�ʼqX<&> =t0;��C��t���_��]q�e���:m�t���|���<C��<�';rg���:Ɵn=h/I=z|Z��\�Σ���*�:;a���O	�r��;_#]�(�3�f4���S�Yp<v5\��Ļ������2��D=*�6<T���ҭ<�߆=�|[��L��Ӟ8��TV��v>�uɭ��N��W�h���<�]Y=��=�.=���<D�(=��R=����xo1=Og[�s3���=:�Q=���+��<Y�i�kr�;4�;�3��*?E���H7�=�c�<��<5=!J������?�<����e��M��<�ټ�vn�,�"��
����<�ٮ<�A�J�b=Z���񗋼ə�;��L=y�x=NM= �&<�P#;Rq.=�yƼ�-��8_���>=4�3�/7=?�+�;�t<w|<��M=��U���/��4�<��μ"�S<�l=�!U�販<�7#��b<p�e�Ksl=o0
���<�;�<3!=�}-;�]=*�=��1���$<z����^���;>�� �<���<S:�����=���<3��<��׼��o5�"��r#m;�[=�_���*��ԋ�<��7<oW��?|�<ޏ;�7ID=�pϻ��$�\9 <]F�<����$ݼ�H��) n��w�<��T���<�^���."=U�<�U<zD=�R�:V�+=Sy��d.�����O��:4'�O9q=k�N�o��O�;��8��`���=��W=��<8���� (=�==��0� �4��l;��>=��h<(�D<��9<%�5�1N<�Ř;oM�f�ϼ�-T��;�<�&�<�B���X=��=��%=��͛<�*V=H�P=ٖ$=��D<��ͼT��<Q)$=�᤼�0���=~�Z�uZ��iW3=:�<�G�;P<���<_[9��ļ
h�=i»��;�=bOk=��T=��<��<-I<=r�ؼ�����[�;�\�.H��_�C=8�A��<v�8=g#y�_�=q(��#p=��<=<UE<1�^��5;u�<8�)<��;y*=��=eC���p	=��%=`3_�,��8<�<=��=�RJ='it<�S=�����:V=y�#=���<��B=rQ����<p��y�<y�|=?.���R=���<�������C��i<�����5�<Y'=B�<�ͼ�1R:�V6=H�=L9/�$�5�-����'R<�,=������I<q�<��������i�a��ʼtA<m 1=4gJ�ٶ�<h.=�+=��S=T�\���<ӎ>�?�Z=�@��Ʌ�<�i���[�;�l�d��L���թ޼H3�6��<������<��<8��z^9wQf���>��'=�k>���=�4��f%=��T�fQ<.k=V1ּ
�<]����<0Ba=I�@��N�;<=��%=b?<07�=�q�<�'�sO�t<w*�;;�L��;*�=��+���=�м�J;��$�n9<Y��/\�<Iم��]=6�����=0������<�H�<G��"O=��D�u<Լ$�<�R=�'N�@d�<�	f=�CW�➟��8=��<�2j<�G�<��D=\�:'�
= ?=�:�Q:x���<��a햼��i�A�<,>�����<�(��?P=E�;L�=6/=��y���1���L�zw���X�����Y�<�_��7׼�̤<Nz�;�(��
�<#0�C�2=�=4����h=(=v��;�QE=I�H�mCu;��<��L<�D�=S꿼�f��PC<q�<���<2+r<";���Y=q=��<�����y4=F�%<P�2<%�Ż0�i;h0f��6e=�=?�k<��z=��=g�V��E�<0��<�Q���
h=�ZX=`=�4R<Ƚz<�p�5.S��N;\�<�p��e=$�:=��G=t��C��� =Ps5<��=k�
;O�N�
E�����$����Ѽ�¼,��������_�=Jt�'�7��9�)
9��X�<�vS�|�A=��9=s(l=}��:}�<��=��넻1�o</q(<yv��0�e��(V�V���`���<�z
=�1=k=���:���|��B]�I���/�����;9��_=��<T&-���}:=$f<N
�5>t=�]k;em0�Ș=jX�<��)=�|���]=o�v�:�м"-=�_��Q����:ꊽA�r�|���]7� .��H=�E=��ػ������x=���,�	�F���6�<or���W�<!J=�z�;Z:Լ.�������0=��8�C�b=zw�4?= U��}�;��k<Qå����yp7<�;�J���0<tԳ�P~$�W�<��μ%�<^�m��A�pe�<o+J��g7=P��<C�<�&8=#� �=�U=�G���8=�� ���=wa�j���h�<k�P<���<`>)=��}��,�<w=�I=7���12�<�x=��ǼƔ<=������g<bQ�c2:���w�{�<�c�<!�M=�tB=tc<9��<,�ؼ��.���;w{�<�Ҽi>I<+?4< c=�J���*=}xj��w]�<��Q2���K���(J�e�< D,=챬���Ѽ͓�;��<(
�<
��8�<v&�;���t����������ǣ�{�߼T����<��ļ��p<5-_�����u�༩�]�w��l��*c��h���ڼ<���,�<�U<�㟼nJ=���<��<\�>=�ͼЧw=�>A=��� �t�m���<��� ^=��f=k�����L��=֣~���=-o����<��<)�p�C�F��� ���@�EI;#c��z��4-��92��X9���]c�K��<T =~k=�p�;t#���.ؼ�`B���ͻ�$��q���i<E�O��:L���=ѧs=��;�=��!�V��e=��z=��<��¼Sś<�7r��o<��Z�p�n���(=2[=x
��o��2�_<~!O=�(`=��-��57��GM�?J=i�X<�0=*Ye���=V# �Q�=�e�T�9rB���=<��'��T;=�N�<���:=�6=�&"��ټ/0V�3��	�=v�g<�?-=��D=U�G=�z���y�5P�<ZB=1i<hI�J$�<�=�=8%8=U�=ɱ{�#9�=�;�<{wK�e�9��==�=j�5���ռ/�ϻKA~�
g�<���<U��i�y<\�=�i|� W;�+N���<��N�y�,�!�r<�i̼�.v=�*%<�� �b��< d=<q:��\�<PRS��{�;A��F�M=�6�<^Y�&=^�R�
>���=�b.��Q�����;Z��<���<�DǼ��|��l�U�R=#C=�;=�<�sI�����7кs��<5e=��仩�!=�	�sp�U�k<�:B�6P=*��<�N��*���ߛ<�(L<�����������<��(=�6
�C¼(p���*B=��1�E��<��E�|��;�0��U(<��+���;FB�<J^=l� =@#G<۸<&!�<�ܸ���=�6���z+=��!�'c<���X�W�=��F�<4D'�Y�<5@=S�H����==T�9�(��_���=
�O<_�ʼ���<F7��ׁ��ys��;<gS,��='|p=�^����,;G���G�<@�B�M�=[/=�p<p�E=1�<��/;,I�<�w1��h	=\�>=����A���Mi�ֶE�����n<�悽���j=�<���u[=	`�<��=t�'������X<���.aq=_E<O����n�1����<z��<~���&=�<�m�<=+����M-a��E�<3�(=���<�E��"^<s�=,0���y=�*#���0<1ϩ����Vμt��;&��;X=���P��<���V�<Y5��<{`��v�<ʵ*=�(=�����&�<�M =��\</g޺p���V�&�^�������'�;$>��%x�?
Z=ިc<�S;g�C�q��;;��2�i�]HM=[�=_$=u�<��Z���ۼʢ�<* ,�M�,�Ȅ9��̼$\�<��`=����;���L%�<��e��s�Mp;�,�A�F=b�N�~C�t��G�=�e�JDf<�C��E��PM�{h�<�CL�>�5=��<r�(�)t�<FV�]�<��@:���<=Ao�<����\H=�9U=�^�<(t�<𣂼�5h=	��Y�P���<>��Ǖ'�t�����T�LN ��a>=�u<��-=��G=^)=�N�<>�������=��=�OX=M�k��=g���X�<�,u�}IY�#:4��;�ާ�	��1A=�>�<��G=g_R=	:�<�H�`Q�K6\=�^���;�.��4�#�;��л�jk=Ѣ뼆�f�j�1=nM8�Z�.����;s�$=��ʻ)=Ԥ9=/%�;�Qy=Z�l=XC�<'�j=����-�<FG༪���tP=1�<uM�<Ń��gH8�Q݂�f�$��q�<ӳ��̥U��S!<(+�=5R1�nt<%s<́�<D�=�=�8�<�㼩���5';G|��B�G=e��O�:=4�=П�<5s <nfi=^,j;q�g;ު�<��<=��<�=&��=&�o�>=��<p솼���;o\*=�{2�{�A�Nj�<�H�C��	��C:�Gc���}=�	�;���o���<X>:��V���<��F�����wy=X3�-�<%}'=0���$�<_*=���
��=�!�ټ��=j��;���<̓�����6���\B:��<{���+���j=_s^=�D� R�5KC�z��<�����)=�9���_R��:q=���.���Y�<��;�{;� e�|�˼�rP<#�<��<��r=1񫻋=u=�V<[�;�K;d+S=d�<��<z��<�S=6I=� �=�@U���<��#=?S�gq��S=8�^=�~�;���=�����ļ�t=$CF���<:�Q�J4�"�A�����_ƛ��u'�l&�#�*=�X�<�	��	I�<0�"%=��D=G��uI:��O��A�u[��ټ�|��'{ʼkp%=���<d� ��З�����8^=-8�<�N=q�"T=.�%<a�~"=e;�<&)]<K�d=,8	</z�����; 6�;���;s�=���<Ž=�t��;<�IA=޺�<_�=��UC�9)A<9Ӽ��=|�:=q�=��%��`�<*�K��e����L���k=���~�X��bd=�Ab<���3`=��;�f,�l��<�>�B蔼���`X�8�3�0�:a�� �T=�8c����<��;��}=
�;+��<��<!�+�s�	<�?~=�������@�<?^!��=�;\B7�mN)�`,���=D���ʺtw�@�=FT��v���c�� =�T�W�=�;��<fxH<�bһ�齺~�,��{<��;�_׼M�N�K=�su<"�<|lr�x]���f)=T7<=nQ�=K]'�1��CΦ<�[�<<[&=�<=F켹=Q�{"�;��=��<��;\u���M�r�<�=���V5��]A��4߻F�$���7���o��=�<}�=�q��Ǉ�K��<'�<<�<��W=��&<�̻t�^�������%���~����8b�¸8���ܻ?�>�xI��0� �H_D<L�=%�)�Q��Qӿ;ˎN�IQ���A����<��%���S��	="p�;�it���<���;х�=�=� ��Y��r�<3�ʼ�K=�I������j<=��b�;zC=���svd�<H �<��<�#U=��2��p�_�H�*�����<�}<=NK=K�<�q��Y�O܊�'w*�hڤ=�}��7Q��K��I�~G=ƻ�;�U5��Z�;�cļ�=��?=�_:�f�&<+��~N=���K�&=�V��5��<AW`��/�+j�$`\��&e�1���$���*�S=�ѻ�̼�uW=�) ��w軡	�c��	��=	!=�OW=G�I���<�:�v?��]�ۻ��=�,=�rb��A��~�<W�(5x<[��<�;ܻؓ<�kƹ<���t=:}"<{:j;i�<i]�G����;��+��F|�.�#=�(/=�1�;�A�>�?<��`u(=A�x=��<�p_���g�2�z���s���<�3�<,���
�<�e��KC���?���,�欔<bt���,;/��S=R/�;g`<u"=5IU=����̻��=��{�=�m=?����H=1��<#1��O�<0_�<,g����E<H�=*����'�%��Ƽ��A=�1���a�w+Ҽ'��<6�D���(���/<E��<<l��<��L=���:fP��<T�2;��-=y+=�bF��]��O���"�ü�Vb=j����\=���<��=E�F=���;��d ���=Zd/=m�=����X@=�ܼp$����;|_�;�φ��+^=o#P���<����B,�����n< b˼d�T=I�)=��ϼ	���#(<#�b=���<��<�.���d4=9�S=I��=��r=�]m����<Eߜ�v��<��@�LCż*���G<:>:�N�<��>�p=�`=�Q=���;J�N���=��<+�O=^��;r��m�a=���<V��<�z5�8�_����$X���<��,��{��=�3k=�(O= �!<���9X/�?�=�B=~�>����<�ݼB^E�.�4=|9:������Xb���=�?$�f-=zl:��c<�{'=ޖ��`�X���?=7� ��P�-�<.���H^����<�QW;9򑼜�<���U<�=$;76>����9���;)<�h(�; v��-�d=����k0=r�5=�8�_;X=�w��=ȇ=�oC=���<kn�<�d�>;�H}=�?P�=�.;�c/�49=d�����&��?D=����5=ܕ����*��=	 $=��<$�L=cwl��<��<X�:�< =5j"=P�.�;Q�o�G�S�8�Y�d=��S=� �<����D=C�<&ʣ�����P�ݼi>�Qq	���}�j�G=o�S=GO=Hz�<�R�:bt;@$Z���ɼ�}?=�+Q=�J=y</���Ʈ�<��;�D�.�MW�<�E���<���<���E�;��ͪc=�F�b<=�m<~~�C�=��B^=�U�wح���e=�8<�y=ߤ�A%�^��Vf=@�O=���z)=�6�1=�|=1��v)��k�X=藍<���s�:?���/��<2��<��A=�V*�]�;����M�x=��<Gk=�;�Cp=WR�M��0�=s<�?=ɘv��4�e��;p��.�v�E��a!�u�=�iݼ�L@;j=�]�k�<��D=����7��;�I��<4�Լ�<�=j9Ir7�\B��.=��-=�T�����<H)=jwR=��"�rM�������\= f��;�G����~<��m=��;I �jt��u�S�y��<W�K���^�M���u<^��<��}�a��^)9<KR����=�01=��	=���<H�,=�Ƽ��09r��?A�r`5=�pi��=yU=l���N�<�_=��Y�<8\����j��:h��- ��\r=7J���xq=�ۛ<�=�<�4��/_<�
w<d��+?��Ҽʾ�;=�/��/�<�L㼒	=���;��	��{�<��<��O=�º�So=�s7��M<�@:����<�^�[8�����Bd<et=R�<�C<=Qe���"�:\�<;�^��$���O���	��<���.����Q�k���a�q�<�pA�K&�<��='������<!Z	��"��j�c��a�<9s>�/z�=���<�(1�JL�8	�+=�Aa�&X'=�⋻^�=�0�1���.%�yM�W�"���E=b�ּ��'���ϼ��=b��<�S��#��ւ�;�X=T�p=��*�j��<�;)�]��;w�M<�:5�co�;�_⻌��<��<��6�fO�������@ͼ?��I��W�u�ٺؼD5f=����*����9�B�+=���=�<#�<�I�����F������϶=;��p�ټ�M�4ｼ�'$�=R�=!#��iH=1��<caH=�B>�xPg=~3ڻ��6=W�5�b�0<�M���[���s�=�#=�c;�{�+=a��;�%=��`=�=3z�]�G��%���S<w�<*�;/i=�K���<W�3:ii�<B���<-������\�	�,���뼸�@����<xG����>=5<sF��;P�z��<���@����V=�J=g>:)�b�#�X=��;F�P�%b�w�S=a�Ⱥ<�:2?/�嚚���/�e��<[�<^����1��T%�gK�<��4=��a;��l��66O=-�"��<w3G�3�|=b?���N/=�M�{k�<�/=������<�Py���Ӽ�����r�F$�<��k<�p��8�\�,G���y=���9)?=��;�x�e��F=��=@>*=NV�8�����Y��\��;X�+=������Ѽ���f��<��N=�==����<�5��ؼE�ؼղ�q�<%�<u���)X=��<����"�;3$�:�.��s�<U�<c���h={�м�ɑ�9��`W\���T�*`@<�L�Ρ��@���8�Д'=��r�C,+���<J�`=Z݁;Hj��I��<πI=揍;|%�<LP�~}�<��n<w��<�`<�ި��[��TG�<��<Q/S=���<*�8=�5 ��-6���U����<}��<���<�j�nE=u�8=c�9�<+h�;Ht׺�M�<�)���&=�[1=s��:��/=|�=Z�="����<�FH=u%4O=����q�;�oj�!������9<�!
��9=��<�eB<�=�<�ed<��㼱D=vE�c3p��M=��>�����H`=����<�<�7H=���<r4��#=:�&��U=�:/=i/P=.��;5��<1Q<Y�ʻ!-�<�R�;�7M<$.o��X��S�t�I=O����=.�8�.����m�F5�<R�+��&=�lE�X,�i�K�"�;n�=�#9��6_<�nA=�m=Б.��Z�<��<D�<|��;��=m���6Ӽ���<9n�Vʁ;�.���<������L��̦��5<���rn�ۈ����!=p|5��e���R==�TĻ���@��;	�6�>F.��}�A�3�)_]���/��m'=9_�<�J�=
Wü7��<�T��z�<�a8;�"���#�9��;<P���5<rkE=ک���:�%���<�s�<�[��i�(��v0=>�< :,����<>��:V���C�N=L�<������N=31����;u�~���	�n�D=�E�=|5��&���{=@d�ܒ+���v<؝ �]���� ���=� ��C���d���j�F�lʤ<mN��h�i���\����;}!c��W��D��<*a:=��� ��<t�<��L�C�=��s��AF<]C@��8O��Y��+=��ڼ�H<�h=�[J�y���=�)>���t��i��n<
�G=ـ����<�8s�<IW�7���8^��lFؼҤ��±�<]q��/�����1�<"t_�էg��-=��k,��e=��= ��HQ={-��$;	����J�<=���V�Y3߻!�<bR���=^�;�'�<1(>�>�5��u�<8�!=�U�<�gG=��s��|��Z0��ݳ���=����,����;�B=��Y<���c��=�=�;��=p'�<�M*<p�
�֤G��ޏ<��<�����*��;���{@X�=�������MW=/�;�;(:�j\�)���=G�I�@�Ҩ�<bT9�lxu<.=Z7=	��
�<2��{=�&���<�+�v:>�_^=T�;������:	>4�ZC����)=>�=�=ܼ܈|����<���<�{)<� �;/�0<��>=�C��G��l1'=���},��Kb="Z[�l�t=�Ym<�'���4o<C2���+�;��l�9�������o J=�u �f�2� g-<82]��n.;�d:1ic�B��ϻ�f�<�L"�������R=��-<4�6=j`m=��=����_ײ<��Z<�j;�#�<��&���o=�R;��U=oŉ<�����,�ȥ�<���;��,<y��<��t��ƾ����= !��r.=��=�R׻���;��I=졮�و��&ͼ'��˭��^J��5H9󈷼��;.�.�ܺ�ۼ���;ϯ��tZ=�ȸ�IC�&�i=�S$=)E��T=Ą><>�)=k�B����Mм�z��"��Ȗ� �E=m��*�u<�>=~����<��Ǽ���<.M�<,q��XOB<5��<=�����X=l� =<�;<_=�;�+=y��<�0�<��;T��E�V=��O���R���=�3鼤ܼs�f����;P6�(��;�
�|~7=%~g=�.I=_�|���l���(=�}�#'*��P�<�ؼ�+4�U�]q*��6ּH#�<��e����(����R���*3�*�W���1����=P�@��ww;�K=fGN=a��3�:��[:�N����;�;�Q��/=/�k;�e�<��(=u$D���7�M��4:�<�P�<�o�#�<?�1�c�R��K��\='��W0�< �C�pP=M�==.=E�7=L�<>;��-�=�d*���==��	:<T�����ż�X��M����=i��� ]=R��;���.��N�<4�Y;;5Ҽ~|�]$7="xϼv&(�p��Qy��dj]==�<	�B�X);�W�Th����#�<(�;'���o�YP»���^���{����=��=�h缵}o=Ҧ���[%�������<6Rp=ϲ��@ż��'�t.D=����[��^�}�(���==�	n����<�Z�<�e�;�zw;�s8<��=�G)=�r=����<�0� �`;MSJ��S>=�����@����~ˣ����ucR���8=�!�<B�r��.p_:)�鼑�B=�<�m�:ǅɻ��4̼.$=|+��
�<���<�>b=����=�(=���<}&�<�NW�,��b9�<ԉ/=|-��R=[H=d����!�tU=��z�`�!��u	;���>O��f;<U�� P�r�V<Ю=r?=D���:s��E='�E�4�<zُ�!�	=�"=3V�<�%�~�<�j�~#	=\�F�;9�$&����=]l=�����+��x�m%=�F�<��=�v�;�ţ��Ѫ<���6NZ=��+�]r���<�Ke=�y=GE�<�W�9.\��ؼ�=S��	�4=��h�ԈY<��K��%8���(�g[#��3ѼJ*��wEq=�?�-l+=�SM;#o=f�=�l�!��r&�.p�:G<��N�<h@����E=-�V=���<H#C�^�^=$i�;a�K;I I=
��u�<;?n=)t=�s<�������=���g��<�/�<�3N��{�<�%=�T=n�=`L;S?W=|�<Y�ļ��]=(9Ǻ(�R�71����A=޽V<~j�A=%�E=�@�`F=��s�����D���n��<^;=*2��#=1��<l�<⺜��[�F��ٌ�k�o=�:>=��=�!��N,�1�Z=}6n��!:_�/�vΝ<H�d<���3���<-�"='�$=�� /�Zk='|��}f_��R#��d;��.=���J�5��<^,\�x2=2��<�=�#=S�Q<��Y=.:<{�%=(ꂽi=J���;w��D=�:<G'%���'�#a=��<��'���;=�؇=+e^<�L<�bQ�� =[Qg9�^?=�>�;�	¼�m����I��QY=JOJ=c��<�ʨ<� <�Ou��l���9=�y=ܕ<q�=�5�<]�.�R�0����h������khA=[�;�{Ǽ;�c=#:����<sz ��f༟zɺ�e��,�;��;�� �M�L=&�=��8=u|= ׼B"��#�Q��<�C�<.d=�A��oO���(���<�R�<���<ؼ,=� ��'=����<G�A���`�Y���<���;D�g=t�}��J*�_L�I�#=��1��q�<.+���;Z����/�%��ȸ<ڿ�����<E=p�.�F���&:��X��¼\q,�7����K<��:�q�_��KH�MR�<5���<�5=O{+<�wF<���<Dhn=�E�����<.� �@��=�&�q�W<>�Z�-"���<S:��</<�=�<�/=/�=5�=//=�H[���<Ӏe��Ǽ��p��<�z=bk6<��<2�C=�Ǽ�/��$m���Ѽ���<�0=�$="����<�&�<L���{����<�U<M�;�;��1�<�a���(�G(�ݕ=�/���v�<��4�o�]��8�ԇ�<4;F��%o<�)=X�f���?��[�<�A=�F�<!bJ���`=��=��4=ш�;N�<�4��� ���(�>�;�Q�@�@�$=*s
=^���d==�䳻��<�U4;�f5<�c��A<n=�D�ڛ)=���<7,,=��>=�f�o=��<��<WP��B(B����޳-�I��<���<.c=�J�<�{�hi�o�ȼ2��<늉<M�����=7�D=ck�<�q]=n�Ļ3A=��p=gx=}S*;������7��B���d<w���e&<�H<^86=>�=�D�.�S<W.Q9� =s�U���	�+6������?=e�M����X
�< �=��f��⛼�l�<�黮CM�Ҝ<Z:���:a�,�b���q�ż��b�4�=V;=���;�E=N:$��\�^����ͼ�/�:�);��v=KDû�)�<�Z=8^��i�<��U=ˁ�ܽ$=��H=(C����#<�wM�"A�:��=����\[=;j=Fz��5�<D4 �Gt�8��0=���Y�{=1�X=c@A�i]:<_Cc=���u�(=K*�*w4<ZQ�\ؼ���+{��I%�;�+=?:����0�$�
���O�,����AW�����=��i=p�ǻ�c�<��=6=KG����ګ�u���b9�ڵ;=-K�<�tE<H����/�<fۻ���D��ݱ���9��/<�~�;ί �cå<�m�<(��ʥ�:����M�<��=�l0=��A�K�<�Q�ٕ%���ż����dZ��G�}[��
��<hP��X=O��\�Q���9���J=i<a\p=��>�2_�=�'A�i��;PW�S�/=���<'�L=��<2��kU�:>w��s=b b;-u6��=���ꟺ9\=�/�;ty=�����;<�Z��J52���k���<�#Ż�TK��&�<Upo=�
�=Z�s���=�w� �l<X����՜���`=h�C�X��;�+��%��9߿e=�[�=��G=(2=�<�N�ޤ<_桼F�!=h�<�J���d���"=tB��Ԡ&��/o<R��9�֢�B���t���~�<���8&X=�B{<���<�
˼�_!=�y��'=�N=��^j=�z�������;�A���Z��hh�������<Y��<�Pv�b�A=E�#=��"�BC�#5L��U=�lX�`u�H�A[(�9��4�3��F\=��3=��h�܈���<�=C���N����@'�!�o�3=���!�ȼG<m=����`�<��c=4�Y��SZ=�M=���;BYۻ�=d��<|,6<�q�<^�>=��=����Im��c�<�ż,���)��p�3��Ha;���tu0=&=�<��b���<�;�n��S��=5���<\��l�2��׼�  ==���͇��6(@��z.=.3Ƽ;$U=��}���e�����mwN�
��Xx��H¼)�a=�����hK]����x��u=��<�;=�o*�GO8�_�B;�
�<3~N=�Z����x=+!���+��x�V�M:>c%=V��3=�Y=�
�=µ<��<i0���Z5�-���%|<6��<��1���
꼔��=dD�A��.*�\<�|׼�v�����.�ϒϼ���<y����=�A=A�=�0�<f	=���I2+=(1�N[==a�:���1�0�X�33<=u(�<��'<�n=*&�2�o=a���[�F<�M�<��=,���M����W=�kL<%��<�f%=W���%�H6��w�<}�;�g��A�@_S�6= c=�f�<��9�~�<&�u=�",=�J�j$=�En<'=�*��'ɻM;ɻ�L8�O�ۼ��w�k�p�\�9����B�<��ȼPLҼ[��<G�Z=Y�<�� =3y=��=��= $<b¼S�=�W��*D���Y;�2"��#�V�=�s�<�g�A���aCW�/�Bs^=��6���ѻ����2=��K��=�s�<m.=��=�����켮Ă��=�Ò��g=t�V;�-D���m�1�=��h=��(=lIr<���;�/W����Q�R�x�&=*�^=���<>5����A<mU�<�=�z�4�OxN=��;=;��J���q�<.��S闼�4ϼ�y�<6H�<��2<�\?�W:��&򼐊�<��";<@=@1=ꔻgC��}�<k�1��=ұ�~=5= ~8��F<�}N=�4�=J'�*����I=��=��������	ɘ��=�`�S��L�8�<�oQ�oqX=V��<�	7��珼0a�t��<�%^�yH;b3O�r" ��<ͯ"�qu$�O��/�<h�.=@I�� ;^�<-Qb���X�T�LK
;W��<������<?5=�>x�3K�cF�<����wk���;�6�!�;�W4=x	<�f��X��*���b����;å�<@�D��r�K'5���=���<@x<�r�<*==�>=ܥ)����<5y��M1��9��5�M=M�6=��L=�3�<���&�<�#=��e�k��-.<K��Տ�C�\�����염p����<�m�<!\��w=@�]=���Ż���r�?<G�(=s�L�s�ݻ6v>��u!��,�9S�%������ռ4��٫<�~<����
=������<kv�<F����U$��|4<��6�Խ�<��I=��_=�yv;N�e=����4����<�=�e%�[�=m�$=C��<��#<�ꪼ:�=�R=���<�<
=�=�i��C�><2�2��.�<N(����W�2_Y���.�{<�r����<��`��&�8��<0<��u�!�x�<�|j=�饼"���u,<�'=J�:��8=�?=��V�6_=�sj��k=���<���<�R!��y��9���=V�4=��5=ML=ʆ�<�1j��P=j+;s`���=���<~U���?�l�<��#<��/<���f��<���ᬼ�B=��<��5=`�����;ʏI�y�;RG�9"h�Sf%=�	=mL&=�p=��;^#+�Е';8qk=}<y�=��<;�*��^=�.�����<<VQ=�_�s
<
0ټ��}�c��;1݇<�n���4����<�<O�<�KK�"G�<��F�GK9���a=Ӽ�c�<��B=Bk�<a�q���<Tai<DiJ��=�m��<x�;Z�#d�/�L<��>=3s=��&�)S����]H=d�����������\=��(<NY�<f=�O"���o<�����Pω=�\��I��;g�Lк�N1;=��l���=#C	=�ؼ�+��� �=�m==�L���:�0<����/���g<��ݼ�����=�ǂ���^�� �u�;� ׋��M�<Pp=ܕ��!��]=�`Ƽ� <P�O���U��nN��2=<��X�|��=4k��\�n��=Q�y=����!=��<������ټ,�;�f�<�J.�D!�<��9�G�ͻ�<g���y�c<=E�����<C�ռ']K<���=(G=�)�<�-M<Ě���� =��;Sn=�f�<z�=#$Y=%��A�]�uxV��ai<8��:^>:�Z!=�8ȼ�Ū<j�8ʜX��b
�|�G=���؄�=������<=�T������G�ӻ��Ǽ�,�;%��<��H<(9*=�G���뼄�����-=Y�ݼ\�=�Ѣ��|����X�WlB=/�����ʺ�;i켆�.=kG�,��<�V=�u�|]�*�;��8<h*==?�<�̖���
��Y=�3�<#<&<v)�<c������Jü�ү<uV��k~=v�5������U������9�3c$��x�<��+�C3���㼳�v�ȱ�;��2�7�=�.v�D���	�;��=�T���<�r����<�p���	=.�<B�U<��<ɊT=�X���=a»��	=�x��F�w�@�"�ܚ[��r��c�;�w>�K��<���1{=��(� �1��w;�o+�	�=�w1���+������5= �k=�u�ؙ<UN2���9��%=NW��0�<�Ӽb�_��|8=�O�qLf<I�мjA=g捼!$_=É�=K�F=r�t	�fx��^=��<j����>=C��<z�<�=E�O=�����'�/����=\��<+��<}1�<'u�<�����-�&K=�RG=�P�<*QI=�>R=�U6<��u��0j�~#˼�����=�Z:���Ἑ��<��I��B�<�"=��S�9=#�<��<?��<9x$=.��<'c�J;%�ѵ�;��H=��i<=+l=����!�W<��=Y���b�<�F���[�b�B=�,���}=�lݼO��<,��6$<E[Ѽwb�<��I�C�<�=&�=�i�<�ѹ;��=�+\
��T7�W:�� �;��2=���=���<��N<�3Ⱥ�w<#�P=��@=�r���%L�Ah��,؃�m<�r$>�P1�68n<�@p=�"�<D:;ٿn�f8=��1�fEG="���| =L�S<�����J;s���=b�=`�F��2=��R�ї�<-(:=OP��������<T��<�؅=����b�	��zE=��f=�_�;��<���H}ؼ:d���%r=6��<��<<�1S�bc�:w:=��<�k�<�	=M�
�+�<T�G=w�>��-�<Y�b=����W$���Mj��L�;�L�j!8=�u���#��Vv%�4#ܼ������<r�-=�p=�b����=>�N����e�C���<>L���[X;HV�"����|=E�K=�Nü}�N7K��|��:���ƌ�<r�>=�J���V���8���N��ֆ�%�������(�m��A=Nkj� �<�W"=6�<;��9b�>5<Xh\��� :�'D� ?����
<���=6:+�ק2��ݾ�.Y%�v�.��'ۻ؏�<�2<y4��w�<���A=_i�=eY�`2�?g�2���H����5�-7=M;=��7��3�<j�<�=��2��D	���]=��=���Vl�(����){���?��+�b='����P��P�n~=Լ���MOL�,���26=R�`�c>�A\=������s��Y=�+H��P%����C�H(�>=�t�<Y���="���E<L�H=���74�/�<��#=Z�k�=s<�t�w-=�����w��G�=_h�<)�<���;��'E=���Ǽ��Z��o�<��!��Q�<`��|�v���l���<�y�;v��<��6=R\.=��8<hԑ��ؘ��?�<w;7=b6�;��
<P�������$<6��<dռ�d<DfE=C
q����;��;Ļ~�={���(�<�����,��<T���]���5=S��-�X�'4;��f%k<E�;<�Q=��P=r$3�Yh��M�=�W	���e=�������<9S�����0�<~���s;��%=�*�6��<(?2=�p=2Fż^�N?���*h��Y7=2¼����(>ռD��>3�<8���y��i<��g�
�������׼:R<���UC=|��O���x<@a=CK:�Ĥ^���¼�R��;��<�=q��E�;�N<�#��<�3=��<2�f�ɕԺ��޻|����!M;�n�@GP��l�E�w��i=�s�cD.=8�9�^��bd�� ;�J=�2C�m���Xw=��$;^V����<$h���t%=d�o=v�P�#�;= ;G�ԉ+��@�������=�G2�I��Hl`��Rz=�<��"�;Wf=�����`���<mpq=K��Ȑ��:<��;k�G=������V<�i�<3�<	�s=�֧;~R�t0����e��d�K:�����6=�O���������zE���缎xA=6$t<��=��<=V��m� �u����@ϼ
<�����=���&�=�^��<��?<D!;h5�쐑<KL=�a����:5��;-��<wy�I�5=��ռc���T��!5�S�;H}<�Ἃ�+��;���gX5;�b�<�+�;��j<�C����<#�<hk����<w%=-����;����0;���������
=���;�h�;×q��G���]�f+e�?۹�W�<`/�M8&�y��;��-���*=r����cC�\K��	=@r`�lI9���N���4�}��<�q���<d��<;�B�i��=��<��$�IL�<D�t<�����#1�������[=
���t �<�Б�{b<JOf=.;-�o�@=MjI�/n�W�<H�@<.�<�%9<������ "��D��ΰ�;ȉW��=�<��;�D����u<�i��+�&=���<OdM=������w�<$��<�3�:��ɼ&$���_=@m�EW=�o��L��;P7��f"�<��=dF=���&9�<�
�۪��3�_����[�<��A�ˣ�Z4[=��<҆8��C��=e�=ʲB�W\D=�<0S�M���˻~����ϼ�,|��%8��<����� 輕���,�=�=μ��7��M<iB��N�1=x�<�0z</mQ=S ��(r�w]<=�\T�F�Ǽ5�㼼TN����E�<CC�<0O��nĻ�.M=��<b��<L����E{�!Z��%�<�H=n}{���*�-5��&{Q<�&-=4�׼~������<��;cul=;O=o�� �<=�,s����<���<���;̓�</<#�%��7|}�m)=C ��e<BFA���=�ػ���0=���<$N)=�~R�w6���9O==<�L=̍�<��e<
�V=7me��Â�\�V�g�ɼ0g8=�=����;=����=>G;	�w���MGE���Q���^���V�,ʼ�*'=��"=��=X��<?\��NI=K�i��Q=fY
=c�=A(N��x��9="c<D0\=���=���m��<��G�w$�<�k��L��'�i��V�F���������$�u�C33�#��-�=~s=I�;�tY�-�=C#u�O�=�'<�J=��ϼ@�<�,=�򲻂T�<n��Hߵ<���<v��XԹ��<���v�=�4�~�;+,����<@�L<2��<�>�����9�f�����U�&��\X;LM绸2<�.-=�=���d���==~P��cxJ����;�?�<��D<誼�-�F3�mjT;�Q�;��;��^��.%����!<��"��&�y/=Hko=�Q=��<R==w�<�M�<�`<63F��E;��<��<$j<�����DJ=9]A=M�+�Xz_=)?_=^�<j��`6"=S���U2B<�jE�J�K�L��<�A{=��.=C'6��p=��s�yE�;?K�����o��F�<�i<�K��B1�)I=�{�<��<x݆�,LK;��O=m�]R
�������5<�8:��=�p�;��'=�).=�d�9�=G���'��p��#!/�� v� ݦ;(���2��<ts���p='�'�A��;)��<fh>���=W�$=��<��H<��1��M���I=�[=ʏ�;\%�<�z꼵*�<��<|�Z<h�<=���찺���M=��.��PƼ�Q2=hx=��$=��={+	�@9B!J=��;Rk=Z���Y=|i0��s�<n-��5�W;��=z�<�U�<�B��Q��ц���;r�g�Լ�Ҟ�W7���1��1�<!*�n	�<���:D��<���<䃻<�>m<:�-=Jb鼼w����=u�w���<�%2=ؿ<�GJ�p0�$��}\=�9b=~*	=�*k=�e=��<`�l��HK�]Oļ
� �/1�<o��<ˆ<e'�<���<{~U�w�麬x=o�N;�T���0�u�=�;���3��<}���陎�ɫ<���<�Ri;�6M=��e���4=�u�<�|�av��F�3�c�R��m@�/<�5��9=5���}�bZ�<̾F�&=żꠓ<��<Ļ�����AIQ�xY=�T�ě���=��i=NQ;�4�*=;�E=5�Z<��0��<]m
����!�'�=22=��'=�c��-&��=��y�
�Q=\�`�dWP=�7i�N����.��ݼ���<�μ<�5��Z�:�M=��?=B2�<�}�r����|���vLA�C>=SW<h65<���H=7��@�1=A��=�����E���e=�g�������$8O=�@@=*�D�N�����S=�<ޥ�E	]=��'�v�\;��C;�dF�K��AX���1�F�=nX�<�[[���ؼ+����*@����=���k�{�~1��J������u=�:�+�;�|�����2�<��;)� :��^�$�^=���;�[N=��=k9�<�����;��յ^���G<�v�<|2����� =�`������A��<�q,�|�?=�P~�A��<.g�<^�����=�;=�I�����р�&�=�����t�`5�<���;�$=��:�����uN=}��:w7=��K��l=I�<^�<����̺ȭ���:V�y�׼HB�<l�� �I�cD�<�l<�B=8<X��N <wk��j=3���?
��Ҩ^;=	�<[��=�7�<�=��=S�C�5 ��pU��*=z�=]�ʼ}���"=Uf���+&�aӼ�&�<?�=�-P=�|����:�)���<}��<W�"=�ڼP7���мv��=�B;`0�X�P�D�����=ܽ �μ����*MK=��0���=�<pL��P= �>��G�zb׻�x;��9=;=E��;3���]���^=�k��;=l$<9g7=��{=�1޼.�K��T'�����uH;9X���LF=;R�<��E�)=j1�Ih=��{=�~��W���d��n��QD����;��J��=��ּ��=2=�/=��z�B�M<Vq�<�x�H�<D[=��㼡��<��M�V�t=���9yn`��k�;3^�+�ٻ�b�<\�A����<���<8D=B�/=�s�{��-(=�qq��0=��M0<��8� qH==������J�޼�R���<�~#��-<�	�Ќ���F��Y�=������x<U�%��=�[%��q�;X3=��=�^	���<;�=I�2=uj5��eF<�л&,��X�|<횘<D�2�7�<��|=�.<�_�<�)�Z�8���x��n��6]����<aE=i=(��=�W<�	`���k��K8=�<��[ى=2(���܄�h"��u]ػ�=��=8��H��Ef=@�h=��&���м�h.=**�<��I��<�׼��<���<�.��o�	= ����N��v�@=vF˺��m�N��:]�
=�Z�;p�	=�����1���޼�=�f�Ip���(�Y0�^�n�!�n(���g=Rn1=�0;��	��&����<G�*����L:�<�pg�ff�:	=��=�V
�whۼ�@�����x���<�{*;"!<DKj<�<�g�<a�\<�CD�❨<��<��j=�1*<8��<N�=�9�f&�G<�<�;.��*��<�G�#I=�
=��w� �=��}<$�<�8=#K�<�b�D���6���7���	�cw�( =ֿ_�^CӼ;f �l��vI=�G�=ҽ�b_��r7�c٦��Ƽ{D~=e�9�D�=[
=EM�����J,<��g�8=�Oh<���<q��<06�[�I=���;7!=��6�aq.�L�]��a<� ����������X=�E�t'J<\I��e�E=}T����ڼ4�ۼ�6f<:h�<q�������2����l��[黔r=,���p=�#�;��$��Qs��+	�z�>=�!�<�S=��=fg��ʁ�W��<���;Ypz;��a�|�1< g���<�8'�	X���K��v�<�f�<�<��K����_=��<H�?���<A7<��S�;VD�<��= �H�\�]</v!=� ��F��M/=�q	��I=��<Jؠ;�:;�Ts��C�<n�,�0dƹ}�<x���#>�����9���n=:�*<�H�c� �^sE�����#��<kwJ=.<�Ӽ���dB=�2{,�-ZT=��1���9<K�ݼ>�;���<v�;"O�����<,w�<\�<mjG�mr»��k�@���<ߴ��d�<���)<�G��<���<����׋�;<n������%1<!?���$�<��U<Ԉ����8�.��<[��@UͻV㟺q�[;GnL=dXW�7?ż񏼀e�`�M�X�g=w,=ه�`k�<���\7��r_=��:)6U�9�b=����#�;t*��Ź���I42=w>廃	a�2��%���)�x�=!8����$=>E�<�D�_9P� >�[���&�<XX�<��<�	Q�[���IP���o<�А��-¼\�ټ~�U=4�<� ��.U*������{|4�	k�<����w��' =BK�<���0�<|K˼	�h�q��;j��/E�v������<��˼-�Q��T�<��!���<<J��]=앇�n�ڼ�.���x¼w�M=���<9f�<A�*=�o��=�^���=QL�`�J=xl�Y�6�\�M<R�%=E��L�H=���9�>=1	���<A��<2�;F���@�����2��Q���e\�/�����T���c�4O��=�v<���;�z;ټ]D2�`<�}e=�S3=ܡS=(�<Ⱥ<i�V=�m=��<�<}={�>�b$=�s� ��;�:=���Q�C<\�q���<�-��`j���.�T����~pI� $�<D4=[%=LFѻǈ�<��=Z.f��� =��� �3=�r��Z�;oOλ��<����8����3�ۻ A���S�]hV=�
w�ŋ=8��<���@�]=�r�<����y:�L�g��Ǽ�}E����hNB=_�μ�v���V��0�I=��!��SW=�١�4�Ҽ��r�?�hdy��?�<�[�<�,�4�m=��=�H��� =�;=� +�;[�<�G���g��D;p��<�o����;�L��T=ϢQ=����Z囼,7�<�,<1�6=E�o8�(Y�M�W����5���C������J=J�ֺ]�%=E,A�td2�x�c=�6�<����2��8���z��iM�}� ��XK��ۻ�F=�<�[��xR�b��"�k=9{;��u=�5<�vK<Up��J54=��s= CY��7|=RoM<״"=�0�������;(T=9�������G�w����(�� =�y�<�ü�c-�����B��<�yл(�»s =< =���<'�=�H[��!�;߳+���A=/(!<��)�3*
�A��)�=��|<��=e�g=�p$�?R�<A5�<��+=�F��`=�|D��V�<���;��O=[D<����H��^/=���=�P=�#E�Xr=4%�<�,=�<����@<`T*��(�<��=!=��:�k�=�ڞ<9b;���<�j�;�O`<��%��_���{O=K�D =���		�=;#=�hI��Kȼl�~��>=~��"���H�O��W>�cE�<�q�<���	d=��Ǽ֜�� ѻ,�<��	���=,I<��:r.a��5P�1J�=�$<�#<�����:��>=ڋ8=���;�=T=�#5=�����<7}	���;P&<�Xd=$� =� �9Q<���	=�~��c-=�g_=}|	�F�;��0<x*���A�DVؼh7=�F<K��< �<7/9�<pG=�_�<-_���ڼQ�9�p��H�?<�Q��R��=�e�;o9<�X�5/��%�� (=��;����xk<?�,=\%����B��<�=�<�n
�w4!=l��=�Z��"b�<>�<{�C�T�,=f��;Hj<,�g�<��;c�n=�8��'6=U��<��<l7�����*+=�6=o*�;Dͻ��{=�Խ<��=�=7#üo��<&96=�ht�e�E�Ou[;2�;O75��'���;�u׼��<������<7=<�=-�,���<�n=[��6B%�v+�K�S�w4?�!�ؼiHO���A<*0=��6��n�e4ݺ/�<0���\��N%���.<����d�<�^X��/���k�9'ļ(-�<lh=d�-��5m���Ź�~��];t�޼k��b�_bZ=V
�<�[��Z�<f��<Wq�t� =w�żEE.�O�^�t鍽8E��^��<d<��*���!����m�<в<��K������&m=]~F=����m5�w���%�<S3���;���; �j=@[=�@�<
����㏽���<�=hy�:�f��3j<n�ּ��6=J)=�uҼ@=�z�sT.��<b3=Ü+�!��<L-�< E=j�:=A�3�Sq<hw-=5=�$=�  <�0�<�
=U�:wQ��n#=��-�� =xeӼ�Q��⤼��n��J�,��xc=%kd��R��"���<m=Wav<���<�|�7i��ִ���<V��������C�YJo��C�<�����0=�s9�����!��Kv=M�������U��Đ�CU漯;&��Zf<tn�<g>��؂�ۚH=6��<q6:�����a߼���;L�G�YB<�5�HKZ=I��<Ӛ!=l�E��C��4�_������F�0#̼[�D=n�Q���;�	�y]�;�F�5ü+�4<Ey�;}�l='t=��<�V�<Mk-�r� =��r<�����ߪ<�#�<%��e7�<�w�:�_#�����>|�WO�<�=��<���<A�<=��a�y�=���=6�x�ⱁ��փ�`�F=0D��/9�<�=��i<��x���Y���$=�YS���=&=y����g=Pϥ<<&"=�}��73m;�zL����<x�J��˷���(�5�-=s�X=䝇=}$�Q =�.�)S =��N;k(q;Y;��\ ���ȼc�ڻ��-=�4��=0���=���R�<��1<E=�4��@� ɒ<���W�'�����<�=�V=o�
��k�<�=�uL�Ji!=zЋ=d���ݭ;/B�y��qA���X���<��`�b����u&��Z庢i=8�W��k4=r� =P��<^��;Ԍ���"<d1�]Y��m>�<:=��t�k���10{�%�<4;&��t�<��9�s~\=�L�;I��<�.A=�����X|��c�;0`�<�r=�Q��<�W��Cx�:���<Aɳ�t�)=��<�,�=�=�d�Z Լm�=��<"�5��Y<��%F�m�ؼj��<�&����E=�R�<���<�䁼�wI���>�o�`=t`�|n<ha;=n�o��W���X�����=��=�w)�AR=$�I�k����G=��ü���	;��=[S�<������<V`�<'�
;_��<�+�:$,A=��&���h<?�U��JP=AD5�/�h=ԉ-��	)�ĩ��n<����:�<��Y=�d�8�/=�u<(�;;u��T�����D��Ղk=OR�:ڷ�,e��&=W$����=���<O����W<Ɣ3=$�+���_<�q���z�<@��0l��M=����=N=v��\�<�=��P=�(k<��<��;��1��7;P;q6���=)��'¼��'��&=�ۈ�ƴJ=��=>\(=��.=SHQ;�࠼�7 =�k��Rn����<X��<�,8=ľ;��躮�=Ѧ=�)<����S<g&�<2�F=(_=���<(�<����F*�(�h�**��9_=�(9�V^d�:��'���$��ຒ�J=���&^=Z����L�!f]=����6*=WR=5��<S�=�}��M�<nt�I����̂���1����</p�<� �;Ε�+�4�
��9�(]�|)޻>ߕ;�=�yZ�|H���N=�ڂ�Vd;���!�zL7=|�T=ѡż	�K=�.)=xq2�
R�����8<Ň~�9��><8�G���l��� �Y��;8-�<:���ˑ�^-Q;��D<��<L�0�?�;Հ0=\��Z�ܼj�;;+q��J���@G�B3���f<nO��\�8���pjj�X�S��gH;S�*8ܳ��9�6��r�<=���ݼ��<j�I<�;��)��&=���:`��<e�D=���+\5=t�=<�u�<��3����<cӕ��}����<zc=������<!I�<YD���;�gWQ���k�������O�$<PW����j=������;7�<��C=��t�A/S���4�_=(�?=8�g��8N�<��z���s=v�+���<fʯ;{���5�PN���E��x+��v=N�U�v�;DS�<�3[=��9=?����;���<�r=�W�<��&_5<��=�z{<nBT=f�����,b��<�=YQ\�
;O<jՊ;�o7�,��< =:(��V<$\_��� ���`��l}����:i���ng3���*=YRo�(��<����цN<l�"=�����bS<l@H=��;=GZA�˰/�-��<Ee漳j<��=�JH�[��<���C�2=�A�;Q��b�e���=�m="��<8�`<IS��1�<�G<)�<����9��,뼴.<=�9�6P=��估��<b(u;x���࣠�o�<���^o�]�"��|&�E�:�ҙ=�o¼,�仏e�<��#;�~h��{�< �9�+��<C��[yŹ��H=D�L=�*0=�qe��ZK<�?�(��"Լ}��;�o'=�`��w6�Z=>�:<����<�=�e���K�<Z5P=�3{���}���=1.��;�e�"�]�_�8�9~Z=Vu�<�����WO=扆=�湟F�<�I����@�ը�<\Xo�!hL��ye=t���j7��47�l�=����nw��e�=4tb��$��7���8Z<��<�ͼ\(���-=>eR=��5=L�F=�g8��"W����<���<��=���<J�漨q�<LN�<e.#=��N���<�o9=��=O����<}�gB�`	�
�f���/��9W��y&:-~�<��.<q���m�9����\';=ç��4��=�M�<#"w<6��;]�U=.�+��G]:�#�2ܹ��
���=U�
=NP�ݪ�����.=u=}N	��M�<�Q+=S����p=`��<R,s��^< �t=ox;=3���m�^��Л����<�9�<��=�\<D\=zZ�<�H6��<B�d=�>��<A=%|f<�sO=�pZ�PZ%�w��{�Z��ʼ7�ټw�ְ=��=�e=�6=��;N�����＆5���?=�Z��B�ӵ�;����3�0��S+=�+�<�� =U���K��8��<��/=�iҼ߬���n� �5=��V#���hO=@[��ԗ��c`=w��9��FZ�<X�m=���v�=l4<Hۯ�@�H=/�>�֨?��`=ʀ���=.>=�x=�F<P���1����Q�;���V��c=^�8������<�.�;�~��м�p���G�J�==���o<� �¼KAJ�6梼�OX=�%-<k�G=X�¼r[��r]=�_��S��<{�YV���1=l<$=�\���G;A��q�
=!A=6Ɋ����˾�9���<��p���w<��B=�z;=k
=�o��T��a <:h)�*��<mW���B��a.;��;�ɘ���<����6'�;�a)���&=l2Z=��G�Ҽ�k�X��<mڽ��^�&���es<:��7 ��RT�<Uǆ<
�K�zW2=�=X=�x0���'� d8�<P=%�G�@�a=,�H��a￼�=��1��˘�ث��R�Y�Z<�8P=dfB���<W0��VU�<�����sF=�j�e����1=��-;�e�>����=o!&��5����h��*_=ji�<�$�s�x�0e�7�N=-n�<T��<FY��0���3�<\+�;)�=Pc4�T�<][=��+=fEL�6/�O].=�\K�j^���5=+���5�}ڹ[8�<�c=���U \=�@=��	=x�UY=��<�掽K��=�+=��/�5�":�>��靼;ޏc=�~p<G��<��G=�>���'ȼ�޼�U�<�ƚ;t�T�
)���Gp��	K=�+�����n��nK�y}�Q�=��6��bb��hA���d=���Q4�<I�����<_�4����7쐼&��:HxC=�I<=L>�� �W{=DU���&*P�,�y=o�'=���<�,=s�1�9�<�*(���<���;B>=^��Ѵ�W�#��Xz�.l�<���<*�<�9��.=n=8:��={�%�8V�g}���=E��<��D=�'��5�e<�@x<s~�<�"�;=O=B�z���-��Sn���Z=.<�vq)�c;=���;J�JR<7�=2�K=���<�+:Q�j�EH»�]��cη�@<\A�K�=���:"���&R=#���W�]=3E*=i�i=�U��i�i����
��#F��@��4+8�4C$�G�0:�v�읆<I*=N��}E=�W_=�hL����>�,=�,=f�
<i�X�ϼ�"`�z�b=J��u�	=��/F�<�<|;x��<a�<�d�2�ػtb�m�>�\���3c����<�m'=Y��<��r==���L=I��J<���<0w=���}�<n�)=|v��@<��W=;��<��=e�=��
=}"�����o�G]
={#Ƽ��;�&ݼ��߼�H:=����ӊ��[���ш�k�o=mڼ�<�|=p��<���<D�K���&�D|��Kq@��9���w;�=���<+�:�����.l�=C(=%9滅Qd����BL�����<_�Ѽ�([����<���<��<�th=�[==�χ<6a��@4<I�2�K�<v��DQ,;*6!���~;"�f=��@�;�8� ��<6�<i� <�W<�7=�mq=�q=˫c�r��\�=Qx�b�������{:D�4=�����_= �=�Sw�9K��#`��f��Y3��d%=b�<f��=n��:A�@��9��P	�U�	�+B���7=����뺽�θX=n()���h��Y���<�8�<�A����<A�B=�<�'� ���,G�P}�W��e��<P`5= x=�Y_���� ��_���7��u=}�=��ȼ旒;�����C=1�#��b�;B�=���<DܹB=����f����$���=���F2���W=@��[===�J�<�k�<�t<<K�h;�j�:��<��(��q�JVU=�ώ��;=���;'<�0=̲���4�4��|�<	�<�e�<�;�=Nvb�p�ռ|)�i�X<%�=T�<�I��G�
=a#!=��,�2)�S-།��<�;=��#���<'�I��y!=	2#= ���e�<����O�A��<?_=�q�<���9d\=��N�ֹ<`=�k�&�3���+=�w�<t�鼈n)�����k�?��\��[�<�x���Z��Ր<m�M�1w�D伖*)���:=�DżS�<I(j<_Z{;rB����=L�����;���;$������k<��=�!=k�4=��#=�*�;V��;�N<����=I�G=��=���;�=�<zy<���<�|a��
=<�����<`&������ Ҽ>j����5=s~x=���u|=-N��zm�WjI�w�żQ2=C6�$+P=\�*=��_=�<���9=9}���GQ�L����!u������Y�[�.<�.�<�~��#<k;5=���?=���<xK�<�^���=k*=P�~=�E$���9<F\�;�V�[m�;�y�%�<hP~�&�x=��<��P='h�<����?'�<�><�7��H�&i⼻i��/�S=����y�N���_ =ߐP=s=��,=�h�<�=��;C��J�<��?������ֻ��><���<m?]��s=lμvۼ-b%�6�<Z=�E~<_�+�	mW=K����e=8�x:��;wj����X���n��(������w���<�;?��gR<�"�jA����;�=-���������TN<`Aϼ��'���6��c;f�d=+�<�W��s��<3)�qm<a��<S���>=U[%�i� <&�; R��A)[=��;����Y&���O=w. ��v�<͵�<�`�_�F<�Iһ�2T=�w���u=�q�<Y㱼M�<9D�������u�%`��_ѼI)=@� =�t��<�3=4D�ʞ�<�b3��t�(��6r�g����&=�ŀ<Mh��y6��3�<K΋=d�=bƽ�W%���X���j#�簘�u!q��[4<X�v�OH�����<$N�<�=�w�6�=}P;:����wA���=#/�<�	��'��N'�(&��߭7=�*�;�7e���
=��^��;=G���><��;�GA�otP����%=��=~�:��[�&pK�%�L=�/=U{&�w�%=�M�=� �<4_�ȑм�Q�Wi=��?��O�>�<� 0���k<��D<޷
�>u�;w�ּ��O=-%�Y�Y=k�໼`�<zo/�+YԻC =-�t��i�MT��p~}<�ż܇*��g�<-c�=�i=,�<j��<iaN=��=G�Ҽ��Z=L�b=�tǼzB�����<�t���8��G�<��=�aM���=,b��$C���:<y��9�\; 5�;�Ҁ=��<�*�<s7�<y��;�p��]���悼#E=�F��h�=Ȥ=�½���D=�d�<ڔt�A���E=�Q;u&^<@ ����E���ּ��j=�q=��D^=�CS��ټ��Ǽ�n�<��<��=폑<��?=. =��:�@=�[�0�3B%=��C=*�l��=&=���?��!#=�7⻤���S�@U=��d���.�ìW;<[���~�<ӊ���0L��*���<��p=�3�GKD�aV=�����eɻB*�%�=��*���\=����`[=Nr�<��`<+8�<32X�*ֻ9t�Z�c=�t
���N�nk;�&=/�%=���w#�H���%�<f=8������;�������1��� =v�2��_=7��<�ʟ<h+=��<�+U=�+�<:;ߺ�H���#�<�?l;e%�:�<[�ݼ��o<{���A����;��O�K�h�'B�<�}�;e
<=��;]�!���5=�!O=�k�Rv����ե*���v=9
=K7��+��<�|��'���M=e����M��B�;�yƼG3=4��#�����c	=m�W�&a&=��<���\�����-���F=jK����7=�B���=L�"<Oqg�0<��E���<х&=h��<�t.�{����ty<��;3O���Z>� �.��Ŀ���<����9�G�<#��969�\����U���U=
<�x=���5!X���o<�kϼ�\%�/�<��\�����B�����,Pӻ6E=��~#�O:'�w�ż�Yb��#��ҡ�\�l�v層^��y��t'����;|!�]0H=��<0�'�N\ϼ 7;6�y<�\=�v�;�=)�>�^���=�EF=� 3��e<E�H<��6<f�v=� �!D=3���:��<�Lq=�""<����,�y�Il�<����	S=Ux��)B�˔ <��H��&<�	�G%<�Fw7�=�{�Y�����i=��Km=]Ty<ï����;�����q(��iY�����f:��};3U�<ҥh=xͫ<R��<W�(�_E�H�n=9�D�� =Y��<�;������;��x<�\ =��<�<<�xn=�	�u/@=AvX�\�>=���<>dռ߿u=ۥ)=����P�=)i=>�c;��:=�B�t&��y����?=S6d�J�W�����\�p<���
=��<�\�<�Q�<�A��=o�(=]
-���ջ(�9��=#�$�w�<�1��@9�{h;Q)= ��<�{u�}�<U���=<�����L8��~���<:<����G�XVR=�V�<w� =R�ԼB� =1�/��Cɼ��=�����=��x;����|;�]qA=9q�;v@�;8 .=`<7=�=�6==>�<�ٙ���ؼ�ɂ=���j+��P �6#*=#�X=��S=�.=��O� 1�o^=��C<�\�<~%����<�����˻�px�6g.�dV�<o��)z���#!�m*|�(��_�C=b_���=��W�"Q=g=+kk=�*���Vn�b6<��_�ʄ =�>�R�@ݻ�|4���h=�sg���;�Q=k�@=8�\�&�M=J��<S�W=�_�<�n�8B�;�<�4�<3����e�h�?<��S=�'=�e��c;��{��>\��,%=� �<l�a=DNo=Q�0��咼n�<���;��W=/<8=ZU4�*_~���G<57��F/W��,�.����0���i���<i�<�ck��2=`{���&4�FeI=�C�E��:j�*�804<��;�$�f$+�K�;� )=^%��$�<~u{<��<���<i����g/=!�=�U��J����,=)��<�rȻ_.���%�V�^�	D9��Y�<�>��dz�$!�$�=!N��4͏;��:�/bc<t=���<(R\=HB��
n��u,=�ǻA�R=�����4=!*:���ØѼ7��4�7;�g<�Y<Bi=��C�!�"=|r[=���q�.�=��<���<���Mi<�p滥
��QH��~Y�:��=�z�=�@=�鼈h��Jo�<��=��K�~]=���<4=u���,�;���:)��*�*�|�<J�ڼb՘�a"5�q�E���2��1�<�4<�";����d�I���P��B=HOO�V�%��p�<��=�Z����;�69<}�@<����(�+l=����8�ؚ�Fz�
vL�#�=J��<�u+<!͎<oa���x=�1S��λc�S�w���!�dY�S�h<�RԼ��W�d�F=M�=h�l������9�<�p=t�λ:�s��ϼ���<� 
<O�8=/�ܼ�K�<L25:<��L5=63��s�;�Ds=�h���<D 	��=���|b�xy�=N=��(m�;���&e=���<XV�<oG�<qHm=�g<�b�<T�F���<���Vϐ��	�<�t�<d�A��Hۼ6�S����<"@���h�<�g�<�;��b=���"�<��ͼkED=o��;mpp�rD��	�<	�Y�`�JZ<��L�Qh$�y�q=)6�;�ѝ�DQ��rB=J\w��<=�F-����u"s���ټ��>�&�<�<����nL���v=j�<A�8�F =�v;=�/2=gks��8y��5��b��,&=1r;���;��.}�9�v���.�ʲ6�f���X����<-���P��\'��O	�	�Y=�y�<h�ۼ"�=��p<�+=������Լ� ���V�<xż�L=VG=��ҁ�bq6=�=?=��һb��";�<� �y7�>ό�VT��B?��[��B =U�I<�B==U�<�D�<�0�<̅u<P�<%6"���&=�r�;�6�<ӧ<=��߼x�-�43=I�o<C�
��l=�=-=�І1<V�E��Ǵ��OO=G�X�*2�<�Ｔ��[�_=�u0���<����TJ�<��0=��2<�����P=�ց<P���!:�"�g��J==�:~9�3L��H$��Z�����t��:Ց�Xw_�Y���t;���<Z=d:o��v	< ���Q�<3��<7��;ܸ��@k��7�ͬ�<�B�;�q;�f�=��&�
=�<�;��H󼳴*=�g��;}��C��9=��b<����
<=oj�߭<� [<&i��ƆD��)=؝���=�/��<i�N=[-�;3�˼�)N�tg���r�BP*�ݮ�;R=��#�J���LK�=�י<��ü�7J�����=�X"�<2�>��N�;ؽ �0O������[��;�#��wD���j��;Y���R=>�%<�� <���It�r5�0ռ9y���G<���<��k=�W~����<VJڻە�;iw���g����>�/��?�<��e�<\�"=ay�<m<F6c=�"�f�ռ提�`�<L��h�G<�f�<���@k�1��耽v8=�\��S�d;-1t;vYj<2~�<lv���2ؼ�9����6�"���	\7�M�Ǽ�ih����!�=<n�=k"������J=1�P��u���S��s���ܽ��@=�wR�j�V���=�@��kK�)���ˁ=Ƀ~���W�R��<@��<��<��3=hH8��;^�I=ŠE=���/Q��}�����2e=�1�<��C�T:���6�<tG�7��;��H=�F��4��Ռ�<���<N	�_�h=G�=��<0nA�R�4�@��<��n=��p�8@T=�{J�R�*=��=�Ie�5��;��=	�e��#��F�}=$���m`k�ڽ�=���;�_?=�A�<��|�8�;�SW=��#���!�P�;��=������J/���z=���ɥ�&�Լ�I=���;�0�<;�*�8<l�e�w(=�4�mH6=D23=eU#=�N=��p���r����H����Ǽ�[�<�1;���+��qL=D����p��9����5=ʼ�^B=�R���^Z2=��*<�����=�q=a0N=�Z=�#׼U�^<��E<���ҼE��[
=�<B�:���<�l�<[� <,�9<?PE=�H%�30;��8<9Ŝ<����d=w�h
�<<B=��H=ѱ9��I(�6'�<`ӹ<�zk<���<�3:pL �O��<&�5�{���*ҼJZ<�hk=���</���G3=;Ȭ�F$T�V�[=zȮ<s�0�x=3�W�-�<<p�:n�I�np��U��:qO���S»{�/<M	8��xQ=NN�>�C���#=M��<X�z=��A��<9n�:e*=��N�d��Δ(�J��<��<z(.�M>��cE�N�]�|;=�V�Iϼ��=��)��d������S=�p�<��N<j�ؔ5�,+=��$�����J���<��B=�;=�3�1�߼��=G!'��G<�W=��@��nF=��m���<[~�<q�6���?�1V��;6>=.�<�¼Nc=�A=�0�����~=�U;�n����7;��)���x<_}�<;>==�9=+�0<4+���:ɼ�:��2�<���J�l<*߼�%����<HФ<r��;��D�C�<���	�<�a��==�!�h�nϺ<�\=�J�:�-��{Y=9��xK���b���a������; �=��<[.F<��f�E�J=�A~<{���gS=��հ<���<?�0�� x��S\=��6=�!�;�=<���'m�;�g�<�R�����<�-�/m��a:07����~<jE=;��AR�\Ȓ<��;�+���	􅽒�w�ª<�Э���<�5��*K;�h����ü��9�� ��5���û��@<'_���M̼%&)<�
[�����l��<1��;֖=�S��壼���<���1�<�@��L�<��<��^���=����^����i���b~��~X#����B�ȼ�-���\<=[T��� E�djp;��X�-]K�g��<fAϼP��<���d�^<���Z,��_�S;q���~}<��d�;Β!�֎�<�I;�=�da�r�7=+�ؼgM=��;��;��=�PF=^=��8�=�:0=C}�<��@=�s=a	뼋�=dN9�xP����R;x��}ֽ����2k�i+��	=�v&=1�U��/�<{�Ҽyn�K�<"W޻pG:<
)+=�����.p=Y���F��-F�~�=�f�7�+< �9=q���<��C=zl����'=��;��_=!0��Tb<EQкEb�K$=�(,=t�<t1=�\7��<��U�?�,<?T���׆=:�/=�p��Y͇;5e�<�
=y��BX�<��H,ػ�P���w<�#�<�Ev<D?�Bx{=�!=�o���|��R�<w�n�o=��.=��<<<G�$�\B1=��%�ܼ�;6<�*=��<�)�<��ɼ�H=��O8؋����D�	�N=s~<��<T���C���2H�FR�^�=&x����:
�(����E�Q=�5�����
]�RX!=���<�|۹�Mj<�j<]o9=���<�
�<�:=-�$����)�;=�W=���<�мCg=��7=�U�;(~�;�'=�z�Z�<-��<�\=�=�D������s=h-��U�<� ����Ex������y7<Nk�<2��<u(=���<��`���J��<F��<�z��s�W=UB�<uy<=��O=vo"=06�O�ؼ���<{N�=��~�=�Ѽ��;!8Z�;!�n�5���<զ�<9T���<�#���ڌ�Qi;��=|��<�켳g=�T���f��nf��;�;��1=�_;�h�:=y�L=�<2=pA<�t�V ;D���d3��2=ȵ<;�(�<K˗<V(8��;�������(���<O8=�sX=�֫���(=����]	L���%��+"=��<����x=�$;@�?�����ؼ�6=Һ=u1��<2"�=�<���;��6�J�!=�h��5�����<�%�<}2R�H�:��;L&V=_��<2u"��Y��ƫt��뜻I�=
R <����[L�L0�j�<�U���7��-�r�<o��fb¼��=𶄻-�;�6<�+�<��I����S�#=o;��=��;���<����.���_l=��:=	�;��#�fM'�9�ἰH�<�C���%<8.�Ⱦn�Fb=+h�<��=)�5�==>�w���[=��P<�^V=Z��<��<�����1�i'��O�;6�<�oP<�G�;�lb�	�ټC(;m�=�;q;��!���<�.I�b;��Ȗ]<[K=O�<fd��n1;u����O��D'�qv߻\O����<�,��enE���L=�=J&b<�;6���	=?=e���Z�J<�S�<�S<��{�3��<�?@=n�0�z=�;o=��*����<u�h=�ܻ,=�'��]�w��<<=��L�Ŋ
�d���	=�Pp�}��<�&F="�<#�m�Az��==J�q�x��;}�m����<G��<V�G=x/�⬗<�m���߼������(=PKD=�6; ��<Ol���X
<��=��<XMW<���<����o�/=޵=3uF�6xH����<�ڍ��(g��伇����!=,?(=DԾ<'	���h=R=k�T�w�e�$=�땼��ۼxt$�)I�-�=z�����,<J��<n�#=n�=k=W�ټ"C=K$=�8,=���[T=�?=#�d=��=��y=�e�<��;:� ;�,���|;��!�Io��ʂ<BU�����|�<��1=���<��;�]6=K!/=ɍɻ_ܿ;���<�f=��k=�|=���o��5s�	H���P<57�(4ټ6_=�x{[�b�*����b�X=m�^;I����U�S̼�Z�<�+�<vNV=�X�pD�����}.�;П79C���b����5�iw��{<H=St��2*=�Q�;��I�Z�<h�n�U�<	3�g�Q��-�<�I���]�;Z���Oq��J������t	<��#����6t��̺��A������ܼO$==�y?=�̐:(=�{f=ڸ��N����3^�4o=s{��lq1=��%<���=D�:=��<�D3<9g)������zX<�P>=��;8{�;����P��<�E=�����w0=�%N�����9��Ǹx=�:;�^-=�&5=�_�<l�=j��<�v�<z|<���<��D#"� c��l�<��C�3!=��o=�<-�-��<��<���<D�<�d�<��Z�y��vE��C�+�����I0L���,�#=Y�f��%����<�t��|�-�U��<J�� �\�d1$=B�<y��:2EI=������{��Qi��h=J�O����<��U;b+�h*+�A�\<Vڟ;�3���y=������~=��2<�+@=��9=�˭<�><2�H=��k=�<n=��<�=�L����=K�=��;�ф:��"=
p��4)9������H��-:<Nл�r�|7=���;\e�<�)A�D�¼&Aa<M��>�Y=�Ƽ����ó���?=�� =��kap��ہ��W|�M;�x=<�=��Z<�5���06=��=�y�?�C=�%�<�+?=�3/=<�i���}=�5 ��a:<NZ��}�=Ch�;�OL=��O=��{�E/j=X!���S/���=��?=>���d�<f(j=��<��<�=�l�{;�<��n��ޜ<�xC=;j|;��=��"�R�j=��:�<�ח=4����QE��z�<ur�<��<�����\�t��<I��<dμ蒡<$=�kB��0�!�(=J�#=�G
=�/<n=)�<v-？�5=)2�=^�Z=�`���ɼ5���
)�;��(=j���=gi�;��=��Z=��ռ��h<����Z�<�X�9��F=|�O�#c,=�)��I�z��!%��:=�~�98伻�=��=������<��<�=>fc=Ce+=�%=y3E���<ʧd<7�P;��b=6�>�b�K;�0O���<��W=f�t;����_�<��=��=�.�'���>D�V��<Q�<�\��< �:�<x1��TA�����h=��F��>,=*Cf���=�� �C�;=F+�Ol2�9������Tx<�w;X5�<����3T=3�>���L<����Ⱥ��܌��1�ie=6��<����	{~�0f��mܔ��&a�֦�<޻��m�|�+=~3ֻ�D����?����;��_=�C1=�pI�>��<�ĸ�j~<��:�M�;*�=r�F�E��U�=�\�<-`=`]C�4�W<K�=��o��AV=�*%=bԿ�]�e�\�.=�%�Ȫ<�ݼF���\��<�9������<��<��
=z2=�,=3��{�J��ׇ<mJ�<b�Q�2A2�a\B��S=}i��z����x�4��Z��)V��L=1�ܻ�y��X�<���;��ϼ���v�3=�_��>*�'������<�;=V׼%A��d�`=N
=:���a˻�e��)j���>���<Em�<�
Q��U�<���<ľ���;>=�/�=����$=�t���[<�pk�v ��bټt�*�%��qj�< ���9�Eː=�N��9��;��<�y�<W��<n�;�?,<.��<�J��W� J�<ml�<��(=)}�ث��6@===z�.�<�Nj=*��B]�Y��+A�����Ƙ<�Z�:�<��b/�l��<n<�U~W<�	����f=��V=$|��ͿU<A�,=NI�<*WμZ�<*�j=^�`<��	��ޡ;d=����u��l׼o0X=��z<��f�X"=�9�ֲ�;Rb^=���<����m໒X�<�㼇�弍�J���3���;��<=��+=��=^����A�-�<L腻�zs=�
��9@=o�7=ꡮ���X��<�h�<�D����<un(<�����r�M{u���<�@%=�Q{�+�^��S5�]}^�5�#��]���:��$�<m �g���z�=0&�a�z�ޅ=�DK=�M=��^�bA�<蓔��K=z���W�&=��F��D��a�=�<:	�<�XH����<d߼P� =S�<�wO=vi�<�nw=[~�<�)z�rs=?�O�ݕj�b3������=���P<���� �p��<�W�<��/� �<<ja=� V�8��wq=y���O=d����<.����~�@�<J$�<�0v�����P=GiH<�E�͎]�h��B=�\A=Ԣ�9/[��g<a0\����<2(<D���Xټ?�����:��5�2t:��܈<��7B#=��b=׬��-�<��Q���1�1l�r�u�Iۭ<Ee����<+L=�<�ɼ�&H��q�; U�:�׾<���;�>μ�d=�#�<e@=zYW�_�H�؜�tE໶��2 ;�K"�#e2<���<�7�;�2�t������� �<r. =�g'��a=~6<w�[��)�<��*���&���H�"����ȼ�@!=��Ż{ �̙ʻH��:���	q= U�\�V�Щ.�@b<�F��u�e�F=��<�z��]S=cB=+V<�/Q=��K=(���MD=-���=�Z�<4
Y��&6�������?���O�<���<�P==b]�<�Ў�@b��ӼR\$���8�	�=_�,=S0��>��<���=ό;�¢V���<�wG=t-=/�D=e+<NӼ̵>=(��'����e;�z<�o�I��;�"����Q:�	�;Hm������y��<��u<Y�=�S�W=!E����β�<٫=�:ֺ�)H=�S���B�qO����μ���:]`Q=�};�� =������}���#={w��q�<^�Y�b�q<tQ=嘋<��%���g��Ѧ��7��+Z�����s.�ㄻ��ɼɌS�b?�;�c"<ob�]a�A`�<9����=�r���ڻ~�v;��mS��Ԛ����y�L�~:�;�'�:�I=]s<�E9@�мR �+�=��X���F<���<��=���<d�O��6#=v12�G��	�[=$>1:@S��C�$���m�#r'���S� `p�7|Q=�u�`
=��.=2�U���-=�+�����<�*B=����d=U��<��P��7�<��G�	׏<�q{=;�H��E=*+T�x�X��6=G{a�{�.=I� =��3��9D��ɼ�
�b8?���s��#�� nh���d<��{<1 =��K����#K<��/� =��3�����<xF��
5<�r=�*I<�*��;��<r��h��X����Є<%D�=E-_�����z�<�2��==�|)�64�<�D=��`<�y:=�(<�l=�H<V7&=$[=-�\����<R�B<�ȿ���9��b=�4�%7�<P3=�m;'B�����</<[��;�m�f���*|=�>=��U����<��ǼFz[�A�.���J=�4D=\,=��
=�R='JC<1�"�^���V5�����"�1=t���HM���Լ%��<Y�]=�A,��J=jF&=A��;Am��~(`�]Y&<��"�tB+=W�s;1#�<�(=�aZ=CP=���<X�弭�=�E�9E�QJg�ef���G���<u.}<~�<h�W=daZ=cz������/=Ŋ���-q��@������<�+���<9������<=E�y���M^���D;|-D��v#�F�c=,�d0�����t9=�=1��<��&�f9=.kE��=*�.=��1=Q�ƼI;��	<�;�8$=��-�R�C=�_B��%S����;%[Q����Z�<J�,=��(�<U;qo�z�ϻ�լ;?��<1�&=��<Y�<\�O;LՏ�%�.�A���g;R��g�<E��3&\��=�<t� =�,�;���'�=a3����<YԨ;/M�~���9�Òں�P=�����v������<�u�y�J=��3���<��
�jE�9�<�R=9��<��C=-�;������:=*��O=��M�#Z���3��D��j���뫼�O��E��
=�(=\hI�~�9$�y�a���><���<��Z:͋D<��l���l=H�z=_R��
=a�ּ� l�(C�<��?=,�:u�&��)�<*5E��[M���C=����μ�,�VA=�D��"��Y�<�ui=�`���8=rͼ�/�� �)=��;�=%W�߷��!����)z¼�D�I;����6?���0
�/�<��v=6�M�߂C=� ��%�+��䏺.��<+AE���=Gm<��+=�@��5�<��ѻ��<,53��ؓ��mW=
ve=��F�B��{h/=�+�,Xp���^<�I���*=� =pa<]W���B��aļ�U��g��;���,��+�<˼���<
4��N��Y=S=���<�мu�Z=>������;�b����<$=B]=�!E��/���e��#�_����"=�ޤ��0�o�U>j��h»��ӹ�`=&hC�G�;�����`��d�<�E=	�=h�<k�i:�!�<�Y��)��<!���V��8�B��A�<ߣV<��<�X��2B���j�����WFr�
���c;7ϻ9ş<��s=�GT�br�<�ه�3�;������<�]�<t�ϼF��<��<�?�;~߼8%�*��-D8=c=��;Z��<�d�<�i���@=9�<;�N�C&=�w4��>O���6�Y0j=���M
ļ+%�<��[��=�4"*�@��<�G=$p=x4=e��<���Y9�<���<N��KzK��0H�nr�7)��㵱<\/�<VNG=�D�T�Hѱ��/��b�8
�Oq�< %=�
P�z^[=��`<:dd=��<ݩb��Q�<��V=`=��Ļ(-�җ ���<�(+=�ie=�,(��X=?�=M|'���f=��[=_��J�<�"��!���<�<��4=��,=�}R<��q���0=84�;�XQ�B�D=�pt<Lw`<�?W�^�;=���<�=�;=Dt�� @��{9��Y[�;�V�)qD�O����;c���s�N8�j�;~��\[��]J=�=<�=Į<M�ż�`=�ڤ<�&�<�6<w�:�_y<}���H�<U�<�3A=)�o���=�H��&ּ��=V#���x1�&S�;�@C�%��#�k��bC���;<=K�=��=}wJ= ��< �����=���<�����<�S���'�;@�<`�<��O=/y%<�SZ=�m�3R�<G�M����<;����:ƈ�z�?=T�;��V=�^�<�y�=7�S=f�Z�7wO=�Nﻙ�༩D5<�%<��<����f`0<�^:�.�l=V$<��;�1D���(��}@����<{�/��  ���<�}��P.6�ޟ@=��`�c�伲�n�wO;<ݐ=�r�<�I<�@V=eh4=>>(�ҋ�<���<a-D=�Ǽtb"���P=��=	��G
��%����<�Mh=��=�,=7.0�~���ڔ�K�=��=	歸�]�;4U�S05���Ӽ��<�&=�,<��-<)�<��<�T���B�9�g��'=��<'FN=��l<�)�=��P���:/�
=P��<+�v���<��6=&::���<�r*�j\y��@=<R=G�z�4e�;YZ�<lV=��-V���`�4M<�B��Z=<�\�w�!�;��<�{9;̮=�W=ݻ}=��="�<>��Za=w�̼N��~꼇w&<�!�'� ���޼r�.���"�"�U�3sI=*:�}����?:
&�<�6=!w�Y��;��
=��a_=�8R=%ʛ� 4ؼjՔ���=S����=�%=}��<�<�T7������a�<�ݤ�}��<������|<xo�;mL�<����GM�;�m<
 �'�F=����W�u��?��pT��G�@��G[<�m+=�/���y<:;<@�<�Ƽ��
=������<�6�9�D ��Z�;;ּ���<{��:߼��	�01�<�;�������;��=�ֻ �^���ͼW@�=��A=�O���M�Y�B=LE.=��=�X3<V� =M���}� �Rj�<�x0���-=�����=^�=?��2u��{����������<ZlH�c �<\<�'�˼���/���Q��;؈�<[d�������1�<�2=��i=j�H��;��GQ;�UC�-S<�x�<�=���^�<*���qi�Lv=�8=:C;�==1���8[����ȼ�O��e[��\%i��� a^��H�<!�ܼ��S�<���=�Kh;�u�<6�<��)�1�м��W=�+m=���L�9<��ܼ>��ۗ<BP�;����z=wn�]K��<dO���
�4�H;��<��ͼ��'�1Z/�!�E=O��=p#�<���;���=]=; ����<�o�<-�$=��Ҽ٪�����<?�.��*=�WZ<��<zZ����3�T:#��<6.;��+=n�Ƽs�9=�: =���<���<Xg����<S�;_b=�d�<zG=���Ɗ���V�{�Z��ꇹ�Ѿ���|<�%=b�{��cR�.�"=�n3�m[~;�s^��q��k�)�����;�v��<Dq*=-�<��<�� ��	=�������<A��:�fd;itX=�1$�O\� �'=3�F���<ʙ�B�<Ω꼣�＋��6��u��
�Y�S���;�<%�]������BEK<'��<.�<�P�ql�K�;�F���1=�2�<��,�o
=���=�м<_�a��=d#�
�.�q=�� �ʪR=�����C=��5�6)�;:�b=j�=�o=�a=�Eܼ�I=q ����M�4hY=�z[���:[�tO=�iV=(�)�o==u;.�g\;�'<ɷv=.��0�4=F"�Z���6,?=��`�%�U�w��k'��=B-;L'�<�=Y���|�<�� =?NC�����]R;��(*<�P���.=��E=�&�<����F<6*����=�ɼF$�vJ=��8(^=4t�<`�>=���n
o=�|=n+<ظ������NF����±�5Y�q���[����7=.����I.���������g�N;����nڼ�Uټ�=���=lLE=OH�;gD?=G���A=k!��z<���N[c���:�Z==���#�<�{��KL��!���X�-=�,�B=�(W=����g�� ��<\D���O=�@=�� =3� =�D�'�
�T�/=�П<��D�2��:��+=)e=����8C=�Y��W�<z��<:#�<�5�;?=����B�-ȼ.ȴ<��}�x�]��c�2��<��t<sڃ<TEz={�<ӱ�|�N��-=.$=�=�04=}�1<5 ���=c�= o)���S��~Q=�$�*����=@�|��<ն&��Մ��k<3�滓����O9����<;�<�={�E���z�@EH������	�<ĵ���==��H<R ��Z7i=:�}=��m��m���+�<�~;�|�<�S�0�1�Fi<.�!=3�<�q&��qY���<��<��=W�ļ�/G��nȼ�Sļr��{1����<z�꼐����=+%0�W-�� h�(�=�"	;��g���a=ln0�!��)�����L=�B!��b��(Ƽ��&�Z�==Xi��y��)RA�����@��w&<��ƅ����'<��>4=($C�!<<v�:4�Y= ��<�g���#��N)�v�̻�˽<`~#;�l<=�Nu�&𻾔A=��@=��߼���T��<�T���)=qO�uv=��8�A�BM�S�<�����9Ո��۫��	v=��@��ۚ��5=��!=9�<��m�"��W�z=�	c�,Pn<b��; �v���[<��4=�E�;`��<�$<2S��T��<ڃ�n��<5�;��	d���)=>�!=S�<Q��<d$�~�=�뻸��%�0��`)=)n:<[�%=�Q�<@�=�3�;�sX���|��?=�^c=��\�_	==>W���3��UAd�I]���,����9�n=��<��U=1ۼ���˹��lx<qo2�N�=����k)=�H�	c�<�W=��e;�ɼ�(����<7�3�����@�~��ފ�V��<�N�<��;�ms=�R:��P=��<<μ�x`<�s{=�j��:�k;=^zI��8��M�<vOҺ��<� ��=��+=f����'=�x7�[{����;!ޞ<.���=��3��	=֣s=7�<J �<��[���t�ȡ
�J�@=�i.��.�<c���]�W!��#�������I;d��ߪ<�B�<����Ŭr=+��y(<P(s=<����@=��/=$���#�;�n��<�z�<�=#�׻�#�<�V!<p�J�RJ�E�+]μ���Z{#=pu=,�����&=�����>=�	�آm��z�<I�<�x���Ҽ?�I=<�*<���;sd�A������ꅫ��~лg=�[��rG��^�=�"C���n�}2=_�=����s�:�uq<�A�;kc��%y���Z=��?�>��5 O=�C�s����5��nO=�ռa��*�w�s@;U�=O�V���\�|�=��*����=��<�=��q=s�H�r5O=�x�<M
��vռ��ü�5�6�00h��0¼���;¨<[�_;�N�f�t<@x���{�<�?(<���G�*��I�<��?�����=֫�<"=VyQ��܊<�K׼J	�@+;��	�ї�3���k{�%�N=$��<��<2p�<�?�;�a=��Y.=?#����0]>=��j�]˼]�4�^=�E�<�5=?��֞<χL=ą�;V{�u#4=jx�K�@�E�C��sƼ��'���=��(�[}ܼ�]O=j�<n������x�<�M�C��2ɻ+*<֒*�b���I���A8p�7<�b2<5�Q�B�ü�U�"Ԍ��m6<��L�Nr=:1��%<a�=�Z�=o;R=d�%�F�'��30��J=��C�q�L���?;�/'X��1�<+H)=��=��X��>g=N�=�<C켔�T�2r�<�=D�A��Su�D!s=Q�=d��ץ弈J=�5=��;�M=������;����`�.�H=�?K��B�:�Z;�-�b�B}�;�w��	��,�{�<O�=���<<����c��R��<{J�M�/=
�<��<��<���<�)=[B�<�A�=
��&<=���LVB:��������g=C��<B'��xB��ɛ<"��<����\#�6�<������.=�+E=po�<����R��O<#��%�r��l,<���oL��O�<s)�<2��:.�K=���Q׼��=?v��	����)�8���qY<^D<I�d:e#��_˼�׸<I�j�p]<H� =niM=���W=q{�*@<Geں
���V�<�I��\b�X�O<�Y=u3=��ü���l���S�<}�<��]��1<��g��,=�=�H�b��;BY��H==�K��(�׾�<B4a�+w�,W1<|���0=Ґ�:6����s�u=���V#��
�==��=g3l=���n�=�
�X=��Q<}ĺ4���}����z������<�<�#=�!=}A_9�=��5=R<���	<Iw��	�<59߼`�=�CJ��F=��_�99�o��5=�V�8�߼Xu�^Q��E�=|˛<�ɼ7t�<�3=f��<�-=�L,=moH��]��3�<��S=�s��-=@�H=��=ec�;;i��O~<凑=7v�ʴ�<
�;ʧ`��D��H=	@f��&�<�"R=�V��g4=8V��M�;��_�U����>?5=�eg;b���f�d�������;�'8L����?���Y=�!����@�<f��<�ۄ���=����p��< 5G=}k�:�;&=�c(�΢�;�d�:0�#=
�1y�;kxa=�u=T˼PMr�d� �E{�:"���R�����X�,=�g,�4LƼ��<a�<(|�6u@=1����m������=�m�<&��<�U�(:������Y���{D��tD<a�=b�<D�&�ط:<��\;��Q�#p"=����Pp�{�<��;9�<=N*J�͑
=}=����{{=d�<4N��3߼���<R<]�滚��<��>=��FF�<��ż��O�7=ӕK�b=��M�f1s<�H���y;G��9�&��� ���7<���(.=T<�B=獱9Y�Ӻ�Y�yjO�"��<��'=�.���ml�0���1� ��:���=��B�v��Ϝ7=��]��P<lp��TՑ��zQ;�Q=��,��o���6 �3r|=)�;!��7���t==���<'�"��7?���=5�/��n7�b=@�b[��0/=�=�s�<YyX��	>;�ȼw���8޼��z�9]=z�]=��9�
"�;�B_��#���
���$���<`W=�~�;>�6���=tz�FG:=��<�̥��Fu��h�����b�U=�3�LY=�M�
!=�/=(0X�a<8�&2;O�V=u�����|�<�g?��&��aas;�򵼆�D��z=��r�Mƫ��*.�yT�<�����Ի���!��:4�R=\��<�����ؼ�|-�'=2��<�)��-���6���/=���n�N��ge��)0�Z���Fa=%]�<��
��� <Uk�<�Y�=�A�<���,��x��n(�<��=x�w�ʻ�9Vi�:�4<$
ļ\�<	�4<$j;���<�<�:@���08��j*��9��o(<N�==pMH�Z���P���<W����4=�/=�`��lļ��� 5���=�C�;dzJ=9�=��&�_����<=��_=@.�<�-D�C>�
㵼 �һ�+Y�Z�'<w���o'�O�#<b�0=嬀<td�<_fZ=�	Q�����O= M=��Q6��<p=�}%=�c=��<	oH=� =�!��<��P�B=�X����;����SR<ϳ���ż�h@�J��=k�W��Ý;ـ<�탼�,U=�qW��E伪�P�ld=/"S=mѧ�C=C|<���<]f�<�Z��b߼\�<oX/=_�<��Z;��s�A7�I��M��<�G<M�`����4m=|�;�,W��s�$�,��y���=�:7�<v[��d=0^�<�B���Ї�k.
�8[9<J�R�Q)�&}�� �i��jJD=^�=�[�������������D�;t���6=R#=t=�e="�V=8t�Jۼ-f��U+=u	���;�z�=�SR�����32�'P��I�<�<ֻ��X�7J�<(�X��kj�Pg���A!9-�7<�$�f\�z�����<V��<�6�9��!;>�7("=~)��<��
��Z!6=�3ȼL�h=��W�뢹�q-�O��:3�J=x+���2�5ܼ���<�aT�¢��;�<N�=�lk<��8�-��<�a=px��pe�<'�\��>�<���L�-`��6*=�s�<��¼�z���7��r=m),=tiE=y���A=�yڼ����ڏ =���Ϝ�<8+ ;?�\��HJ��d"�H<�U�;=�+<��@=|r =g}�<�]=dV��z4v�r�Bȁ�-�g<�2���%���R�3��;�E���<�=�9��_�<}�8< ��o�5=�7�^ �8O2�9��<�R����6;
B�<��T�y���f�������t=�q�<��!���8�� ���|O�����'�<�ļ=�<�C��2�^;��4�ߋ�;4��<�y���<=9�W���<�Jf=0<g<\�S���:�B�]���#=� i=)-Ƽ =n��Y*=��
=���Z��%d����ϼ���:�|ݼ/lû���,(<߫)��T!=��c=)���g����=Ʒ$<�?>=��2=.��<=�<n�y�K�c=��7=y�<]%�� X���I�<wI=	����?�� ��!e5<�j2=�·�����3���l���=?8E=Y�-�3��m=f<�bY=��=�1_=bXe=^��<5(�<��x=��=73��	�?t�����9o�p�<[w)��W�4Bɼ?�#�?cN���5a��;��q�#�<�41�̻Լ�>�<]�*=G�<R1켰z?���q=�~�<�Xͼ7V�܌��xF��=��.���A��=��^<�
ټq��;���<��B=D�;�6��s�%Q=��s!=ϝr=Dg������O��<Qj�<֢�<L�r�`%̼8fV��ܳ<�24=8k�@J:�*a�:������<Nk�<�8�1<����kV=�t�<-T���c�������-��#�v,&;4h��=W6��):i�F��H=����?�o��t�<�M༬}_<?:~;T�:�*�<�J�=�F;K�=+���� +=��<<Dټ#KT�阬�g/����=��t��m]<LWe��)��n�`�
=��R=�<&=��+����<n�2;�PZ=���v����QU���ӼXK=:�]����ͽ=��~���m<��H<F�)�י�<{"@<����Ҹ<�n=�"��fU�UH�<~�G=_aU��Y^=f���*��yμyż�s
�`�ؼ��<���9��	�v&<�t�f��<`���o=�����
�$"]�Rp����y������<��<���<IG��[Q̺��=�N�<����O�v����<��z�_=^e�;��0=DQ~<CC<)��<+�=�V���ѼQ�;�ܼ�ϼں[��H˻_H��s�;b�I���%=\�ؼ}N$=�:�<�n��*�>ѡ<�kC���<�wĻ�@d�z�;*���1#+=����t^=��1����<�?��¼�_F=m<�l<6=�&3<�e��ٞ��k׼Oк���*=�$Z=,=o<��ɼ(�)<q��;M�6���O�ü�ꁽ�&�ţd<n=�?���@=BG��d8��j�<��2��i�G�W�/�=B�޻�U��0T=�{&��☻_.K=>��<�h$=�>f���T�x��o�	��;9�>κH�N�� �P�=�W�<ˏ���"=7|��sT�Gi���=��;rz��@���J<ˑ�N�j;��<�ļ2�7��0��&�=�Il=PkI<֧�e���;�j����D=��-�sx���C�<Xx,=���<0&����$"y=1+O�7@S=n�;�g=�)���<mP�^X���N=��=B�=��<��2=4�==k����4�n�7��[�=p!�~Y&=�<]�:��=R�<#�G=��ʉ����x� ��E����1ݸ:���<CG�<I��ʬ;�Aüᤑ������3=zm��=��M]J�d�=��=I���m���c6��RH=\��<�o_<Bj�<�=���x�X9�<��;v
4<�pʻ/^��{����=�Nv���#=#����7����c<�o��?=Y�(<��E���弴(8�J�<b�=���;3��Ll(=V�<���t!��}��[�������:=���<��l<���<�Cd;x=Ι�;��;�����{<�rﺭB.�q�<�#=�Ɨ���<K� �5�=���<�#�~�#<	�E=�E�;�
T<.��<Z�����<߁�;M�#=˥;AϞ<��Z=��(��R� ��;KMQ<U+A���B=ܛ�a�=�CK=KV=��Z=O �&�ϻ��7������=^�Z��J���'�;h�i<]=�ԫ��[ϼ��ټJ5=l=�1+��o��c=,I=�B"=:�g��y�<1��w�}�
�;ߗL�a�=&�<!Zc�m�!s�ĕ=/��<z6���F=ڵ�=lԼ�[P=�J�Ԣ<����%6U��\��,���њI�N\����0�6�H<�N�<F3/=��T�q��
����:��<�dɼπ������#�֥�z"��94<��.�-�<��f=�K8���<YF<j
�<v:�<Ɇ張�G=V=v�<5#�<8/��=+	=�A$=z�<=��<�F���4=~Q,=�\=6�b<<�^�;��:�1�>0��f{+<�
μ=�<�ۘ��.O=���C��y�<���<���`�컆=<�j"=|�Y<FRb=��:=)�!=�F��Mƺ���xƼ�_=�����@�RG�n3�G�o<�)8=��5�I]5�;�׼#'+���~;�����I<Қ��J=N�%�ۙ��P����j���<u��<{b%=v3A����)Z
�����3�<��;� �)q�0|0<Я<# A�Æ�<ٳ�>JD=�%����Х�<%3=�h�4W<=����L��X��Q�ל��&�TG��x�`��N���V�<��U���ּ���<'��<� =X��<�9���,�<�귻d�W�ϓ;�J���9=�VG�jo�<��\<J��9�>=x󏼔|�<n5F�\��;���-�k�/��!M=�`=ƥ=H�<�ͼ��!=(q���bF�͈=�@S���#����;{b�JZB�ԑO���I<숼�$'��K�;z��<�?f<T?ịJZ=�Y;\Nͻ��,;��F=�sY<gA�;� <�/��%0M�:ǹ<G�=����<Rz��<�r��`D=��ּ�$��q��<�I=�j3�&�<'ba�H�=���@9�<0y@�N� �@�h;^1=I�<Z�����_�K[?���a��h�<^���a�Y��/!���N����<6�n<�	2=��&=l^3=%�J�ؒ;�H�;BJC���l=W2&��J<[�o=A�:���;�ؼI^�<m�'=�ۏ<cE��e���=���<b=���<���g��Gש�R2�;�Ƽ��<\;A��h��v�o�r�1�3�\K�<Ȏ���S�<�"��<��6=�=�u���0=��Z<�(=�����}-�a�_<�>=��<D+�<��<��	�R�=I&��=x����׺�&�:����|H��k�u=��μ�_l�5%��n�&��5\�>�h�,]=ᣦ���a=�����"=�A#=�wI���[=ڢ�8J =�_����:�t��z	<�!=9=a�8=�MZ<�?=�)�g.�]~f=#y<!lg=�;9�0�<*$����<X}<6)=6�"��
=�i�<�>��3��<
ǻFpO�d*�����c:��=�cQ==᛻�O�o�8�ڼePl�||���ڼ���ןJ;p"���k<մo����=�&�1>?����c�<�c[���;�B�K�=0k0=��<�嗻�����u�O��΋������#7:Ҟ=
5���=��ʙ�)���tI<��<[A?=?vżW0Ƽ�'��s�Q��;��<i�(����1@�0�b=��T����<���<F&�<��<��i�B��������۪<:?u<��;�)Q=*	
���2=�]�<�y�B=<�=�+$�pg�������ڻ�7�<�X��V
�'�O���Q�.o�<��L=CO��X���<��L<�1�/�:��!��F=��ͻ�����,�w<�=O�<m�!=��P��2<:�t=d��<qcҼ���bi=E��<�"���<�Q����]�v5=ݱB����<�ӥ� �c(;�rR<V\4=�s8�%>&=���Q�
�^8P=��(=UԼ�-X=\���;��<����LF�=j$�ai.�E�^=��U<�F<�-���4<�9+=���<�-E��R+=^^T�K����<�/��\߼�u=T�H=��==0
=pI7�)\/��� �1 �K�k=[򼦝м@��5�n��b=�M��d�;4~	��X=t�<N
�ş�9��:Ǧ=L�"=C�<�!=�	N��Ǽn	=�����\=2r-=/G ���<����6�<�м�q��h����<μZ7j=�"�<�V=Wڥ< M,=ZI��|3��Z���U=�!��;==>r =;Q��&�<��H�-�ѻG����r���R=��=�l��h��<R�w�x��9ԭ
�F�v�X��<�D�k�Y<����K=_��<�Y�<�Zs�`�R�x�0=�3�l<.��һH���u=��\�7w*���"�3�R=#h׼��@��6���hl�E�F����D$=��f=�˂��?:=��r����<�c��Q�;�~������2�λq�;���<�}�<��X��Ñ<�t�U*F=&��<�b��{��@<�C=�������<=g�<G"��h$=&%=+G=�)�U�.���>=�ņ����������<:��<�~ʻ�l�m����;5��=��;1ⶼ���<5�=��d����<�Dg=c:R�γ��z�='@9=�&X=����C�<����4�/�J2p=��U�n=��< 
��{�<��(=S�P<2^�;���<�.�<k�c�->��&���TN=�Pv���>��eI�2GA<=*=0��N�<cс;�5 ==:8��:��"����cG��P<b07��c����Z]���<q�����ݗD=8�=+"�=H�Y=O�g��q}<?�a=Y�N��d�< �Z��B���i��-ü��<=��=�����*ͻd�;.�3=���;y	\<�"�<�(<��=�_<���<�%=��żm3���B=#��GPq=<2=��Ƽ���<֦�w=p����=�_�;�~2�����T���Ik���D=�s=Q>ͼ��+���(��^z�!��j �;>��T�B=5�ܼo��9������<5<=1�==�iħ��ĸ�_}D��<�(=�ĕ=�+<�Pr�C�F���(��/]�0�<�Y�;���z.2=\���S�;�͊<���Hҕ��r��y�"������=�P�!�˼O�?<v�3;�¨;U�^=*~���s�h=��]�lSc�i>=�5-9�K�D�#�m�����;E�<ɐ[=K4����!�;I�:=�N=���:x�ϖ=�����+fQ�?�<���<�BZ�T�`=o�N<e5u<�"����=r�<������h<�]u<�sL=oD)��z4=�n�B=g�"=?P!�PB�)=?z=��b=��<x�m�]������&ût�9= 1��[ �<��1IU=�=ܸ}�i�l<|��7;=(>J=/�1��#G��%e=pr�<\*	==����iû�ő;�}����\= ,=�E ;����:To<�c<����+�����:8=�&<�V;d�=V6=F� �l�|AX�8�2�W�$=��<��������/<���xwT<8�C=�_=Pǆ�w�Իi4�0���TN�9���<�u������=�yl<�y`��BT��	�;�kk��n���<�j�<"m;�=G7%��I<��s�(��x�<��;"�¼o@)���w�gy	=%�;<�e=4ˋ<�#����g�J��<v`_<G;=�vü�x�>���C���^��[D="�u<:�m<pA���$3=�E=��¼xZ��,=��P�cq�<��=;��ʞ=Du��k�%{�<|);;8�+="�<W׵<��$=�*<��t��@<���91���|<K=x=Q��Q�����<�N<�%.¼��һ��	=�����]�<�u�v��P��d`���m=��U=�G��uږ�u��<�b+���<jyB=0"=\�[=l_��(��B4�<E��=��
��w=(/�畈����<n��<��;&ڼ�2K�uc&�'Ay�L�;F�j=˰���y;�S2={���?[=�����~]�P=s��0;��<���=޼Y=��Ӽvq�<��}�f��<�=f[3<��<�<�<"9=_]f��K=\���m�(����lp�_��<�ȃ�Y�s���=��=s9�<�9?=� ��t=��<���d��<���;��W=�f����=�D�<ucüv�%<�ʐ�� <k&��=*�<�ߐ�9o��h�x��L0����<c�����ʼ�)b��I�=�Q�;& ?=���`n%=�=F��N���D�<`��sZѼ^y�'󦼙�z��dj���\�:`z�A¼�D=��9���<�e��s=�U=����i�&;�to=��~� �==�N<�<=��v��<#���L"@�ѻ.'��*=��<%\;ƕ1�6�<;U2=ʧL�->\=�<;i?��ub���Z=6�0�9�%=l�B=���R�
=@R;5i�;$=]4�<{�*��JJ���G=M�_���s^k=��<a�q���h��#�<!sW�\�g��Ҥ���x�� =��^;Q��=q&=�/1��S=�P �0�=$���߀�:���<�1=��p<.�<�<͈7=���:���Q"�4��;��i<-�y<Q;�B�=�eP�l�w��"
�f��<�����<W�3�wF-=KL=k��<���_X=pQ=�_�@n(=o�r;?�����;5��<ͮS��g�<М^����������p4a;J���tX#=��.o_<q�(��<*�=�C�<aؼQz_=��=�O<�M���m3=����m�=����Z�<*�2���0�ڒ<�����Z<�-	��/i=̚k<��;;�<;�� ��Yp��P������05��T�����ǈ�H�t�	��r�~=<V��aQ=o�V= �<�j�;C��<�-Z�?O=T�j=���<���;�����μ�=̼���;������M��ݴ�<�v��b?�<'�ź�뎼D�V���O<���;S�V:,\<=��u��
���=�@�3~T<+Ď=0�
=0��<�G�����;���;��|=���g~�<xͼ��߼������Y��<է�<X���x�jk�6X�<ZW^�ay9=�y�ǟ=� �r_N�8<����f���=�s�<���c���-��zG�e�<]ꅽl���)�:����<��� M=8�L��I�$T漪�8���=��6��<�����*�X���(�;���;�+�q��g���(�=�z���Qy�+�e;��#��(����n�e'�<%F'=W�$�������F�?$���<;��6�;�%d=q�e����N�:=�3�<�B�<��Q=��0�<$z��O�p�u���=k�=�v�<���^�7=�T�<r<�G=�(|��5�7����=�s���L=��<O��<}qҼe&�<mf�<�l���(��{�<��λ��ͼ��<T�!<�V�<��,�@U<�=<ü!����
=��L<�-�;��,=�0�Ϛ/�H�S=K<�{V=��3=o^[<��=�8<4s%��(_���=_o=��L��g=�ە<y�7=S@E<zIE<�0.=�����=0	���/���<���:�<U�G��K��x=��B��)=5�
�G�;��=\k=����:�X�V�p9=�&�<����� ��w��ˉ�<�:�|?��9d=�L�<"}M=X|z��;��<-�;u*(=|a=Q��	6�i�Y=)�<-������p�弒8�<��o=�e=ӊ��{�a8�L�&������%��?;��9�
=�g�L����:*��ʼ5����1��=���g�S\��b��*��ʀ=&�C��;�;E�;Ih�<�e�ٿ�<rO��_�<���<�d=�8E�Rl����?��<b�<�<O���Z;���b�4<�14<+4�=e���E�	=���;e7�;��̼tҼ8�̼�R <m��2\��q�&=�<���P�!�мmPպ���<}$<�Ƽ�(9�ON�=<���7<�Ũ��9=�8B=O=L=M��;ÔW=��;�~���ŏ:�ȗ��W�;�4�?���l���}��<��B��l�9Ts���"<�F_���5�R�q=�NѼ0�!��\�<�W���%�X�+s�<�~'�A�˼�K3=�㢼>�F=� �*�B�q��<�y���3=�����'�<�?,��X<	����� H�<a�<��a��Q=+�S�i-��2@�����Ӻ��N�ħ���V<H��|�#=����J<�*��Ż�oռH]�<մ���D�(��;�<1�@��E=��X=�5�;�����@�<m�<�;����<+��b�~�+%=F�<���	����P=��Y=U� �3��<o�m; ��;G����I;��ռV<�<�E+=t�p�6R�e��;X�<�F<j=�d=]y=fB5=�8��������j�Zw=	&�N�<ӏ�F�»^����ûY�;t���F=����|[<?.�<#�9=�&=�p�<���<K�t�����z�;&^#�̆<����LN��=H�P<�;�X=�� <�=���<��d���(=b�a=tg���;.�Bm=>)�<�nW=&�����!�.M�;!�<sM=5l=�^ּ�G=xC����ɼ�&<���<���<��Ҽ�G&=�q����=������	��<Z��<)��<u��<�S�P���4=��<>"��2|�u�ͼ6���=�6,G���ļ�Z���I=,��<��A=e��<���d7�+q�U�y=��L�e=ī��g6F=o�<�����g4���;+� G�
�R��h��id�<��;� =�k���l=���rJX=k��	�;���_=[��<f둼�Ҡ�t��;��(�*S�b�:�}$�`�,��Ax<��I���B�׌�<Wp��Y�;@���<���b��k-�+����&(=S-�<�&k���;�`��Oø:�r<~�μm$��5�zd =�K�;x�<�<��Ͳ=G��<�`�z���|;���l��X����<C(�;eFY<�N����⺔]��C8��ؾ<��<�$L<|:�+��<��<_��S!м�R�<l�I<\�ؼ�A�ڈ=��'=�<�io�����߭@��S��f>=����+�O��<m:5<�ly���ͼ�Pa�u<�.<<l ="�	�%!�:��<b%9�xF=W@��(u��h�|�T;��g�9@:=���0i/=
3�7x��V�ڼ�a��Ws���C�_n,��㊼��p=M�U�eh7=dq<<�Qp<]	=�=gY4<�T��5=�� =��|���-= �����4�Ѐ�3m;-��<ZMd=�w�SZ�<��9��RC=r�==�a���=��t��*�CP=&`=}EB���7R���<��<Z	'=?�R�ot��b`�<];5=W���o׹���<ҵ8=�>S=s6�<P=���<_=݋"�8��<n�ݼ>�=�.T=e7?=�\�/��<�BR�X	��= ��,�<i)=mh;�ï�I�0=l;<�D�%��<o1_�UTS=�E��@�r=YK=9����<�����R�� �c+=g�M߼�-#=��~=h�TH�<PxC�z =6F�w]V=b�z=��?���<U7@<��<�"��<� f=�A��[�wH=���<�>d���X<��W���<�Ǿ<
�c��Iw<�k������'=.�O��8�<��#��6=� ��<v=c=���<�l<�Y@��YI�@I=c`#=P��<[<�<�Y�0u <�=C�?T�;�G�;r�F�S	=x��<(�Ի��;ɣ���(�j�L<|� <���<[�&��;#N��e=��A���]���t��<̑�^�=��F�Q	�<BR�	=g�<c�����=���<E ?�q��<O�_=;ҷ;�t̼@z=��
=Y03<�k���8��6�/;ᢊ�UzּR�=mV=�J��\/T=��=�\=4�Ƽ��k���=�(���<e"n<�*�*Ǽ�8μ���W�����(��c����0=a^��F9��g�I�<�O�c�=���<�a<e82�{����=�?�:�7
=��<���<�;Q�8��<�am�,�<� g;��Z=�@���;4�t=Z���&��O�l�=��*=K�A<r�*�V��A�À'��G��yP�q�p�����"����w=�?=jD=s;���S�<F�4=�)�Qk�<TBA=A���<I�X=�.= �w=0uB<�9=���vX�[����<��q��#r��{;�a�;=����@���Zh=���<J�0�o�N<`�'�nS"��F�<�*���PA��+f=,`�����_!�&I=b�<�ĵ� h=F0<�ϡ�!�4�A�<��O����[¼��;�g�y:�g��`�<�6j=�O=���<w��Q�*���i�1�j���e���=G6�<�-�;��b;4\z<�G;���]=y��R�=?ڮ��-<�t��b=L�:[�l=�@<��<��D�71�,[S���c�SK�F =��O<DSĹdѻ�
f��!��I��+�u�Ҽ9�=�0���;j�����A��u=����������I=^����Q=�%r� *���V==�&���6�P�߼�ź<����|"=��E��QE=��E=�,;��������p��W��.?=�����HF=��R�x����R���AS��l;N�p���x��=cFؼ�$�p�������<�><s�E=X����a<��ż[�(���r�tf:���v�ni[=9/���Q=t*W���?=`Ϯ<�ü��w=� =F��+�x+_=��<�v�<��S<] B��=%�Q=��6���}�;˼5he=�8�;�3=�<E�=�>��h�-���;���<��;͚:8xn�L����3�<�=�'=�\	�w}<��`=Ϩ�<WzӼꊽɈG�5T=�5'��n�.w��4p�����-{<�=�w<Q&�š��G<x�:=wTݼ�҃�*�����<�l~=�,�<<#�<���<S�;�+�$S=��ż�W��'��)=��=P����=��=K�"�m�L��~ż,��<]��+S=�}��{]�"[�l�<̻{�<�=c0@��r�ϮA<�f���
�9�7=�y��1�5��@X����<	�4=h�;��`�C�^��.=���=������;�����z�V; ��U��R�e=��!�
�/���8�NѼ��{�(=HcE��Q����Y�=���;�h���@���ļ�g<e�=N���g=��=��'���~���<�@Y<Օa� ��;{��}=�;�G=��
��,I���"��F��4��,ǎ��)�<3)=�5ʼ��$=%�\=%?k=9�S�`�s��;�<�&m�^b�p�Q=�rw=b.V;��]=陼�?1:��Ѽ�d��ݢ;�P<0�<�A�<����\H;;�1e�Q�8<<��<�����k��� 9;Y�Ӽ,J<����2��=2t��G��~����s�v>=�d�<{ŋ���Y= I!�p��8'�����<a�v�mA<�0g:֋V=�H�"�IE�Wi．�S�|w��v?=2��I�<��&=�~/��d�;qͦ<�)_=�+;7$P=��D=K�"=�pW��黙���.��e<＋����CS<�k���c=
�Q=	M<�f=�.����������w�K���=�c�$��մμ,�=,QI�Ua�TO-�]�ȼ��d�m3��+ł<ZU?<2"<<$�<ty�<.W+=�<h�_����5�R=�ɼ2�;��ڼ�{һ�ꢼ��.�WY=������<ՙ$�U����,�6cY���<o�=:�L#=�Ӽ�9����=5E��wO���u�WP�(ud=B�=�n�<�u�E�!=P�����������<�=��h=r��m0�-J=7zR��(`����<�����h=�\�V1�1�1= �=]����<�	W����@�;�2g�<��0��F�<@�<2�=�����+==0�3����<�L�f ����"���n�w�^��1C��G%;@!=�++=�)4=��u;���<e�����;�e=3H=OP�:��{�B �<5ƒ���V=/�<�u=�.�<�Z���N���=���;� <D�	E=E�
�	�&=o�ͼ�v=b�=�T<~�A��{ �y=S�=�e2=��S�q^�>$=}5(;�K=�3=XӼ��'�J��*�1={�<��=��~����-1^�f��;�o��	���#��nm;�U =��G=�p�< �H�$�ϼB �gx*=|�/��j�2�F<''��Q-�L7�<As�:�9�<*K;ļaĖ�.�s=��$=�=�=<P9�?ʼ�ŗ���Y���Z��S���=�h<�uI�/O���_�<[�=�1'�'K��Y8=Y�5=a��:�7�=�)t<c��:��P��
/=��K�ޖO=�qG����<e����`<���=�ݫ<�vQ���r;2���wQ'<�jk�"����<4"��U�=
���'b
�?�=v���ߡf=��'��Lz�1,1=�&�/=j�=��U<,�
<==���ZS={ֻ�Xߺǟ�<�T0=��q=K*�<�����G��)�.��]�&'�$�-&�d���ՄL�h�h�j^޼��<������<N��	e�;�`��*�9<��<�Y���=(�r���Ǽ,���z=q=U=��0=�)���x�<��<���<S�;H�h=�	�0D=D���;KI=_}W�g[;�6�<{=���t�=��7��/�<ن�;�S5�@e=E^=9"���Wf=��<�ۍ�N�=4!׼pY���D=��L��(���ϔ���<��D=�ck���f���뺼3\<k3�;
h�;��=�gh����<�,4�\K1<	�C�<�(�n�����?=d�A=Q+=GY�=g�Z����.c�;��ܻ�><��=���޲E:��/�N;���4��}FS;�ua��==�I�"<B!�H[���k��h\�e8k=��/<ԝ�;��=��3��s��DM2=Ul_�j$���2=K't���|���ֻg��<`7���<v, �?�"=m7�ן��4�<�`f=|�f<%+�<�lI=��C�<� <A�9=y�=�3M�uV�<���8F���@<4����,=m[=<�q켞G5�:}�EW�����"��<ZdE��,�;�Ց�Y�T<V��<�=99<��=�ᗻ=��<�=e�Q		��);���¼hQu=�J�<0ʘ;(�b=)�='^$��S���Z=Iy=��<-�c<��;��W="=_�r<��=
����?=�f=�
�<��_;b�;�S�F=ab����&������==�:NeS<�����R�(�8�_z �k�
��֤��&<̠��ٛ����%�`ZH��zH=Ntk���<���<'{�^��<y�=|�B=ҜɼIK��8��&����<���<&ʁ<(�T<K<�h4��~q<dʠ����7�<N20��7�ԗw����<=�@���L=v� <CVü�C=�l!=���<_+|<S�p�>�W��<<�D��-:<86=��l=C�<���<4ڌ�����=C��<��<DG�v�"<���37=ӘD=3_~���O�{M�̲_�=�6��:�;;�"=�t�<��;[�%=��=� =��k��;�;,D��\�<����Y���tU=�j�O�=ޯ7=Ɯ���4=B-�N��<p������������A=0K=�+����F=}�=�n�����<�}/�>QM�!7K�V(�ݣ
�H���g����P�͏���K��F�2g=fX=#	���N<>��E>��9�\��/�ߦ�S�'���o=�F
�J^=�/���c�<�WA=C�F<zg�}U =VA���#6=V��<ض3=Tx��7=#����V<��=�X=�m#=]-�����.��<7W=�_S���<=�H!�Ђ��!�F������2��)Q�\B�%��ർ�{�Υ0�����=T�]�=|��<���;`G��F;��)��>:�2��;��2=�:=�K8�m�:�[�<�q=�p~���f�VZ��-�=lь���(=���x�f�3Ի; �(=7a=ˎQ=�<f��H�:+�b���<ź��6>������u��Rj���,���x��G=�T��м��6��SؼLM�:�S;k鮼�X-��/ż�j]=~�=�Ӽ�,��2F=@^=Q���t�<q3�+y���4�3!��^D=bh׼8H�;���Ĵ�<ר�;�zA��z=*-�<9��vZ9�� h=��[=� =^�8=�t���iL=��?<Y:ۼA�;�A�<�b��!�;F,<��I������dH}8-��<�sg�n_+=&�@= ��GF���#�<��%=~=.��:�T<��]��u#=�[Ƽ��<� ���
=�������

�]q�;C=��o3'=��{�Ql[��<�I����<H�<UgC=��c<4y=�j�:��j��S�q��qʗ�Z���ۧ�<��d�$�=r:�<LW�����qټ�'�<����k7=�3=[������<4�=��"+���-�QBp�+�;����Zp�W�k=�=ɰ�<�;P=�J=%�h<c���'<~��=�ج�9��<LU<H>��0�Y�c|=�J"��J =B�ؼ�R)�鉴;���;L���7Ӽ��=�3����?��+<`X߼��T���ܼ�0�[:Z���ּW�;o�5����;�銼��z=�v7<�\J����<�C���=�*�<>,����$=�S��J�q<��мB0^�s�0�a��<���$�2=Y�^� �ִ�<Q������T<4+����<Q��<�a=�R=�̼��8Ի����pr���p�4G�<=�/�<��<5=>I��A��i��iV2���l=�J�V�=�36=$�c�B~m=�MW=zn+�*�����;��:2�a=U��Gt=4�G�0�?=�\��K��Y��i;<�(R�\�����<2�����=V~u=8�<)5=� =	^�;E{p�;=��������|�+=T!=��"��v4=��B=�n�<x��tE=�ʫ�e��<�R�:�"0=��U=;�<�4c<���9==B+���o �Q�;lE���=�*�<Ã8=�҃��2x=Ҕ��>���·u<"!=@��:�ż�HS缵^X�cw�;3��n�,���=w'�ȏ���g��m<	�)=��=�D����F�]=+֑<���=�<X=Ӎ���üe����B�;�I�� �<��6�Ղ=8��<�%�Ti=�0=�UP=޽E�a �=,"�w0��Y2<�o=�m���"<��:4��<_R=Dj3�R�h��$�;�4�<�/�J֋�8[ȼK�S�Sէ�7=t�g����/=9<�A���V=�&�"�1�����n=�p/���7�۩��`��<��/�Fx/��?"��"���=�$O���ټ^j<ͧ�<tm�;E��:�<('3�J2��ʻ0�V�R:��,=a��<���<y��<{Q��}z �����2Q=��F<֔C���p���<Q�	=w�<ʰ��Mh�;��m��:L�4_�3U=�8=9�B;��=<�0_<s�]���;�1 =A��<��]��/H=��<{�e�5�*�BL<��(ͼ^㎺1
�ly^<{�^;��D=+=5���En�	H=��;�j�<|�8@E�=�G��jM=f=0<`��<0-=��2��=��2�>+�����P=��g=xm���bJ��4�_����%���;��zF=--�=窲��uＨ�g�є>;�����D �&U3����<��F�^@=��h=�"1��Dc��q�< Kp�[	=�b=�T�<Q':<✻���*<�G�<�?=����x���ۼ@�G<��=�4�<�Ɓ�
�d='<0=3�A���k�����j;=�(����=�-
=�	 ���$�ti=R�n<��?�!���xF��퍼m�=�7<`��<�=��><#� ����r�<Ǎ+����<@2�<*=��+<��<<�(=)=)�,��j��P���!=����<��G�Vf�<$�����������-�1=��;�J`<�]<MCD=����>G�����`���a���<�D-=�1_�P2;�q����}���0_=h��l���#�<M�<ѯ_=��<�{'=ܞ=���;W�I�V=��w��n&�f�B=L��;J�&��f<%�3=�>��~$�<�׊�KM��R)u��M=�.r��J�<쫌���.=�ϓ��=H�A=z뼓pI�?}�<�W:=�Y<q3��a\G�ޗT=��I=�S�qp<�g<su�W�,���q�|V��mo=�?��gG=�,=��<y�d;)�<�iE�߬\����o�	S=�ʻ<�=`��i!Ļn=S�=�湼� X=lN�<̜�:T�޼�J=��<A�<.^��{�;ԺH=Jέ<a>�;k-=�k�<Ǧ3=IA=��)�zF)��"<�޺Q��<re=��s�;ln&=&ч<�����i^=�<qk����:��<3妺����.=�.1<xF4�z^�<i@<�e����U=.�#=�� ��<�r^�\<C��<�0=$��<:�Z=�`�<�0�p���ü>�%=��;�<Z�;�V���gb=��t=)1���b:=�/(=W{S���=�`=3uY��u'�]�0<����!be=��<�<�o����V�=��f<����<�����=�=�S�<M�=�A�<��P��U��8<��R�r�_=���2�^�
�e=3�R���I�c��<��V�bz"�k?3<wu!�����P3��f<�[4=���-<~( =/�6�tv<
�< �g���o��.w?��U��'W=l�,=h&=<Өּ�ȼ�vD���!=�QO���U��##=�G�M߅�Q��<�*#���<r�P��K%���t<�!h=@	=��<4�<�S=�=wq����:-==��~=G*��==������+=t=�R�LaJ�;$=�-�7֔ͼ�d��]��[�_O��<�n<ޮ]���ƼVץ�h*����_<�7���&���=5�<L�<��A�?�e=3#�<��K��3=� ���b�G��
<�<�Z�<ڋ��x��;��;�_j��k��<(�=Wr�����^e]��{�>�]C=8,���>�<^��<��;=C��:ռL��<�;=�8w<�E<=�7�;��[�X��<�N!��n=�ר�<E�>�v�	=��r���+����<���idA��磻���BH�<�e(� �<�=̺�$�4��:O`(����2��d:N=W
`;�U��h:;�:=1� �(�3���#�Y�c=C����4;�o$<]��੻��:=�,�:	���2��HE��=O�����ze=��#��`q=���:�-��CB.<�e�<�W
���"��=�Z<�3�a�<��<��<xq^<�#��s=�F|=N�=!�U��ū��pd�B7���A���p�պ�ዋ���#=H��}ޓ����<��
<90(�?�B�er=���<�=�#�O=TP�<`��3�ؼ�$��J=Y��	��kZ�� ��=p�@��<�1��決��$��A��.� L�o�,��=�L��#�R�Y<B����<tNa<l��<n�o�UU���'��������~�k#�<�3�eVF=9@�;�u�}�=XrU="F�<߼��`�����޾��2ti�RZ=���Ż <N��D3=�L=�[l�P�ۼ��~�$���-ڻh�H�,.�=\7ʹ��μ��]���L�_]��RJ=&Ma<컬<��
��&���_I�� P�FA�<�B�2�F���.����:��N���<Es=[��,,R;�:5=�=����=ּ%c�h�u�|;��"�<#~�:��<��'<ɟ�<�'�<C�%�����yX=n�=NR�j��;ˈ缼f���>��-���+��Q�o��Qm=y*���ݬ���<^��<��W����~]�q"A��:=������j+<ѐ�<��=K��$F��U�<Z�d=9=Q�<�Ｚj���E_���;9���>=/�M<Q�X���T=7��<�ӳ�&�?<��n��TW<�YM��K�ɰ=T7��';���%i�<Z�G��GL=a��;�D�
K=4��<�o'��f;>�!=.�U={�d=C;��ڥ:��<=�+�����<Ȇ�7	z��8g��V����,�U=�A��[F����=WY	���<�� <A�r=�(����=߁�<�YL=t?X<ޢ�&�G=���<�=ߊU�`��<���<����W�=��,����~�=
22=�2��=����"=�
	��1��5?=i����B��X��.4=�&J<���:B�E=����s�x�w,}<-VD�&����X��{��� =��W=�Y;��<�r �ɥ<׳�<4���Z�:GCQ<Ĝ���O�<p�k=��-=7���'v׻��<P(�8 �<�+��=ѷb=+�l=W�;n�e=��ƻB���æ2=�=)�d=�%ݼ��2= �=}�_��X�n:="Z�<��q��R:�~�$�3y�<@� �ap!=2co=i*I�o���AK=��S�� ���M	�9�`9�����L�;���<O��;��x�<��@;��ʼG�/=��3=�T�<�t�<,=��T��
�<c�=��"�)=�<Y=��2=[���?��<j5ܼ��=4�����L=ͪ�;G�=t�ѻ�����i<7�R���<ݟN<�t<��=�Ju=�Ѽ�=�5��^��A"<��<��=�v�)x�<��=��]=$!�;)ij�Qr:=����L1�xӼ�%��#,�$��s<=���W==�Jr���e�N}�<FҼFlɼ|5#=3 F�ԋ�<#l<�D�j�F����<��<��ẑWB�)Mr5�ZY������(��5 �<�#�<|C���o:��5�(�)=Ra,=l輪���yG�rh���W�9��<ܡ=�s�H@���<z��<ra0=���?�F�~\����D�G�4��lU=/*�r8=�]=9/���`=v"+<$�-��~�;FVg=3$=i��'��l�=�!�<�^=|*U����X���z4=J��.�V<���<�����D=*N=�`��&�<�͟<s��;�7.<��<�̔���O���M=1g=�4��:�{<[�.��?eȼ�@=��a�~�=>f��<�y�L�߼���;N i��'q���~��ݭ<u���n��{���<��𼰠H���]=��2=��q��O�������V����m�C�E��;u8=fh=HSD�A�H<��6��{e�3%�Z�9�f���!<��f�U��<C4�<'!D�Ȁ�;9��<V�k�?WA����UU=L���н��+༶`f�$��;K��;c�$j��Oڻ�\����_=����ļ�S=�8\;��:9G)��=a����<�"B=>�=�W<��=�=t�;?�W;3u;+*�wu��SZX<p����ʍ���8!S��J�,l�;I$=W��<|�\<���<���I�\<ɣ�V�(<��&=��`<V{�<q�;OW���Q=U�Ѽ�1p�m7����_�$h��]ռ�v�<�r�<�A=z��<QC_�đX���^=(�U~
��!=�i=2���y�<w��BM<��E=K�h<�e=̮��!�3=i�����;%���tm��]ip����h��<���;+6E=�=o!P��~=�zμ�m��X):��t=﵀�7��Ҋ<+t��p�뼈!�<��Ѽ5E�� ����G=3W'���=�j��>
h=���)���$KK=��=�$=5�r��C��
���Sż�/;)!=�l";nlg�v(:�v<��=.����=��;jz�e[E�%�d�q/��n���To�<?�h�v�^�X�s��u�
��;��J=%�<n������ �=cs�;#V6=f���OQ���<�w���$}��p���o�=3��=�=��q��R��5��ٟF��I��V�<�V��ڞ<����a2<� ��P<��=�:�����y�=��H��IP=J�M��
�<+� �ʌL<u�8=õ0=Nd�=[м;�.��K<R= T�ht=�᡼���=92�;�Z6��ܼ�[�G�5��N4�����Z?�B�=bR"�O�Y=�\<7�=�A)��Ｐ��A=�0 ��Bt;�d���/=s�=zMc�^���(L��,��b�@Z� BH=N�6�1�<�5�C�00�;l��<�&��;Y=N>H=�o=c��2�t�b����<�&�<:��<Z���$B<s]�;m������,�M��<P�/=���<�SF=�4]�A7=��;�[�;��L=k�༊x=bt�:�<���=`�T��N�JG=���/�;@�F����-O#;X�<�!=��;Oh1��Hh�n�)����s�R=�p��8w������4<�_`�C��Sin���V����<q&`=Z
�<%��p�<�F���0=81��?
=��'=�T>��zмHf<�t<ƇA��D;!�)�&< �a=w|��C�^�7OT���3)�?����=�R����Ȼ\AJ<�ټ/w<��P��~�<Z\��
���+=����A�; 5g��D�<��b=��6�����C��3�<�g<-v=iB=d�7=&z��x�<HH!�j�7=�P��Y�;D[�x��
�Q�5ڧ��u�;ā�<sr��f�o�<i� ��*=�'��ĺ<�
ü!��<�i7=�:��Qi=��c=�!�+��<�fo�E i�乪��k��|�*=�/����`�:=� ����h<�u�;��[�ޙ��XK�<jh<@���}���W��<?Xļ�u=)dI�~��<ߢ� ��<}q=ށ�<�|<�����D�ȕt<�<;]t�����;@S�<��+��q"�D<�@���-0;D�-=�i=��_d=�|=R�j=�Gt;Ռ߼|��<����j�M�/�C=kۙ���:�a���b�������Np��09�v��=��S=9�?<d��<��V�8�<ٗ8�3�=�;:=."<|2��^�<��=ilD�Q�m=JB��Q�1��H7=<H�<W�ؼ�ǧ<�U��1�P@ =AK̻w�y= J��r)=��%�6���c�Z���?=�0n;�n�<�U��	=��1��Լ<o>����]��q�;��c�=�4:?�؞乊*F�#.=(b�,�;=R�R�];-=q�H�/�p<l��=K,#���&=B�<V�0�-�<�N��=��=d�7������{���zH�j�R=B�>�&����K�D�k�.�=f�9=��<�
�O=YX&=���A�=���<4@=�b&�Z]?<�3+=�2˺�n�<���y�=	g�<�1<=f&�<��<�x<%��<@�h�-%<��<��o=���=�;�|J'<Y<�m6�<�he=�kK<6�T=N��<y�=��4=~i<=��=u*2=����=��~����<�W=?��<�f=��<�+=�k�;��h=|t�<#h�Ɗ׺�eռԗ�<�Z���!<��%;�7=	ﯼX=��8Gӻɉ ��=P�G��HI=����I���a�kJ��V�#=o���)��w+!=N"=x�=��\��^�0�4�%�$�=㍀=x��;�/���~�;��w=4i��n�<�d!=�>+��.��=VwZ���<���<�Zw�*�*<�	��N��\�&'�<`�����a�=d;�b]����<ט�O�H���5���O�v�J=�-��7��<��R�AC@��c!�$Z�n�<'b���Ҽ8sI��J��������6�<�������� ]B<���t���k�<�P�����<��<(��<L-�7ƹ;�/=ZJ�7�;|�m���6S�o�pm��Y<>�<n����`���<1x��w�S=F��;�17<ky��K�<�EY=u3�:�=�1=�_S=�Z2�G�X��:����л�5��Ѽ�<� i��@A=#�=|�e�f��y�.�ts�<��4=�����;����M�<dV�<�:�<�X��c0�nH<�)&�u�D;�^;g=�X�����Y��y����)G�fF<,���qt;��=�÷<��<�Cx<Je�;�f����h`=�}�:�XT�3X���v�ni:=�g���՝;c���C����,=��&�+�ߩP�5�<Mz=��<5##=CL=�j�=�Q=l"4=F��<��6=�n=��g<"�<(Ii<0��;=�:�;�1=�'"3��%����X<��R��{=~��S����9=?=>{:�\9���a��C󺩢�;��0=kA&=�.�<�^��\<���<U�H=b�I=���i�-�j�g�{@�;0��I���l��L_�<�Wn=�0=�� =�=@�,=1�;D�8���W=���� <R�8�	'�:H�e=h3�@�7����H*��p<�%�oo=I�=K6�<ob���=*�P���F����(=�e�p���El��찻v_�47m<�!=9�/��=�;���;�h<�N����>��=A=�f={EC�a#�j`����,�j�=F-˼��W=r�� D�7~�<�b=x�'���p�u3:�m���������BԼ��a��q}=*�E�V��%v漣 =p����(>=LC��FW�������_��O����W�?��3����q�I��<��<��w�u<8���T*=S�=��<vML= �;.�<�x��n�;�AT����;je����~�
=����t�Q��<�<���<WO	�ψ��<uټQ�A;���<��Ȼ�И�����-xe�Y6��!��<[��<l�����#:�q�P(�j�H=��)����3��(=��!=��;��� k<���<�ݼ�
�O���]#(<��Ӽ��R:KOg=�X|�D�m=S��<�缉�}=�y�;'Һ�[u+�w'����k�*�.=Iq(��<���B=iI=f{p=�б��1<��*��=��[=�����eK<2�N��=�Q
w=���<٢<�v��F;�E~���������G;/�F��<5�¼Z�f=!�=�˳<s(<:gU��E=�3���Ū<��<��%��c���<���T-R���޺)�L�l�,���"��p<Q{K=jRj��_X<IK+�۟�<C|��9x<�J$[=�sY������̣<M`�<9N�;��<�f��u�=�ì;^��<���<H� =:�0=_�b=�^=(dG��1��Ⱥ<��X���< Tü���<��	=��K=��<��<�^�;ܽ)�pQ�;��<�h���>;�+=����n�����<g,��j�����S��j�%i���G2;��û�x�<s�+�C��<T�<��@�0^���=��#��5��h)<F�=�hn=�eB==�μ�b��;Lݼ�Z��[�[���μh���l�;,RB�����#=�(=��>=�1�.gм��U)x�H��?T<�P?���=��Q�T�R=V�=�Q��z,;o�����O=a�t�ׅ��gn�����S�;�5w����r<S�j���ۼ�J��O;��Q���0���ϻ��J�;�\<��u=7U=�/<^�F=w�Z=^=<[�ŏ�Rr[=��l<zO߼1=��1���1;�h�< ��:��=��w���	�%��<��G=>U�<?���@,*��@C��%A<�G�;"��`$a=,��D�|�C=?ɦ<�Y$�F�>���<��%=-,����<�0���|9����<�B=�����_=*&�$W<�B�y=kl�jhD<��I��9.<�f�1�,=Y)5=6�X�������/�8<CW�bv���ǐ<DA=�+�<�����M�]C�<��*=0����d<�3�;�J=��x=���<�7r=�c�``�̉`�TU2=6�Z�o�����=����l����<�l��h�<<F��g�h�:�ߺ<���:���G���K�l<���<�qP=3��N���8���d+=<f=�y�����=EX�;�e��T�=�F=��仿+ڼ-��gǝ;Y��G�;6s�r�f=�z=��*=�߫��� M:���q=h<`<����S�c���Y=�T��G�}��*û�=T�E�	� <��X;�p��'�1�N�@�d¼<�y��ڃ<eh{��7&��y���}�<;=ק��<($v�m3�<���;�f��:'�<z�=��H�C�I=��ܼ�Ѫ�H��(�U<vޡ=�Js�ę
�.p���q��(1���S��;��ٺ1�B�n9+�Ȝ=?@`���=27Q=4$e���F=�,$=5K�)�<�U=#�;g�_������߼�Ҋ��C=3�S��{�Wy�=�}Q=�~.=�=�h�y-���e�<���2X=bBr<�b$��'���ʻc4H�:Sh=��h��F =ҶN�h�~�0N޼��A=��;��gƆ���Q��j=w�1[�<�7������7E=b�F=K���@=W'^=�O=+8J�i-=%Q���^_=����	=���<�\�F�Z�
��<���b�|�L��<�/=wB=�@���>�U��<�'<I�h�K)!=�r=�N=oc<}�;=xP�;A�;��	 <�/�����a���Z��� ��<R�Q�|)���n�\�>���<�m��;3�D���D��j�A�<�#E=��#=��S���^��B�u<��5�e�-=���<�̑�����t�3�:���f;�;��($=�,=Հ����<Q;~�<_X�rz����5��<��j=;W�0j�5�b=xF�;n� =��3�-�O���<q�=���#*==��+=��w=�y=�<ݘ&���@=xs���Ƽ��-<�ok=�4�Ay�=���D� =H<=��<����|�ʼ��l=Řܼ '�<���*v=Zp'<�w���Q=�$9F�0���<驲��2���ʻ0�=���<7:���e���h=�x������H��7�=�m*���'=�W0��=��D=\M�]�`=����=��=v�=+�<;#YT�S��Ξ;���<���泙;Yh\���::��8=Ͳ����<A��<z)���������!�<�&@=]�9�IV=#���	=��p���Q����E�Q=�]�<���䑽�)(=�w�<[��)��_=s�X��0I=��;�=�; �Y<���#M�H~"=*'Ӽ���ܢ�=0x�<J=<׈z;�xm���q=*�ͼ��;ɡ=��=l=j��<fs=DN��h�-=�l�<�U��!��V>=�-�����Y�`�@���x`�.`�<�l��	Ɔ<�1�=�� ��<~����g�<�� ��E=梼�D���;�X� ��;�����Z��sA=f����	��=@ڼ�7���8� M��=
ȼ���*6��Ⲽ}�f=��I��:�	\�ymG=��G|Y=eU��Kc=63߻PNe<��ȼ�`o<���M�q��8�<��=��l<Ħ��o���{y�;�f<~�S=[>�-֭<�\a�3)��򊽺
:�Y�A�.=|��b�b@��R=�d1��a�=��q=�;� �<Ā.���f<��=BZ2������=j��gv��*�3�6�3{6<�I =�T=	��%9����\DK=���9��<��P=���Z�;vS�<������9�N(]=���<|��q
�<L��<in#�ړS��0=�ג<����I��O=�]#�a10��b\<�,=��G)��E+��(��cX[��KV=h�E�|pܼ�w;�S�;�i��������,�<0==�����^�-�=�F�;�<�G��Vg<�h�<��=vC �
��;�)�;ܓK�d:W<���?}=�֛���ܼ�S<�P]<�!�4�t= �;=��]m=�,)=Ww<J85=�E�=:��<�M�<����n=�4=¨Z�;��1c=� �H*��Π<�0�ore=��c� �賻��[=WU�<��¼�?�5���=Kė�������=�P���kƼf�5=?��<|�<�6��_9=D?�<��I�_��@�<�zH=Ҽq�=r������<���VR�<~-��9�J���ļ#5����E�S�>���-�~,;���<��;�EJ ��j'�t݌=�Mݼ�q=��=*�+�>���J=ܟ��h��<�[9;<Lq<:��<�_=�=Ot9��J;�{�<T=�/W��q)<������k����<fR(���ݼ�,.;Y���2���7�<5P4��&μZ�b�%��<?=ˤ�<��E<@ 
='�<
C=.>���{$;��Z��t�<��=�S<"94���6��6%�քO<��[=*�%=u"��a;0���u=.e,�{yQ�C���X,��X�d��rX<ߜ����<��<\�X;���؊��-lۼ7�U���-�ެU=�Iv���q��C��}Ӽ�9=��r<T̼�Yм6�H=MI-=0�<���B�׼�dE=����9=�X���=��I=s�1=\��<F���vW	=�`z��@��V(<�_�;�D�g�f=��8���*�����V=��<6k|;��Y=Ԇc�m�1�e�5�����U]<=P@��`�����<c^"���M=��"�*+�k�8=5��|z��>/���<� �<xMͻ/{=��y��
Q��Vл�1�	�o<���q�;��<g�
���^=9P��8@�Q�̼*��<�lM<J�&������<�.�W����l��<��U���;ħ�4U��뜼��:���;1��<��:7�§�<��<Q�/=��Q=��J��)��� g���[���  ;�,S�dL8��ݨ�&��4��Rr漼�=�����m�oPҹ�6=�rS��>
�E�i=w$����<��]=����5�k�R�j�!5�<�r��9�J=1�=b�<'�;C׼�S�=�| ��)�=�zb=�<=2����<u;W��Z�<+^M��YY�v�q=�/����`=����� <&�Ǽ\Y�<�X8=`F1=)�<�u���%��-�<��;ԍ�wY���t4��&<p�'=H(G�W�<��%�M���@����<%#=K"�<O��SA�H8G�����=��;��=)�g��=F�b�~j<��O��:���5<j�V���)<n��M���]<PKy�y�'=�WV;�oX=ӗ3��&T����;��C�u6���V�[
<��}��� =x/�<�OX�H�^=>�D��O��p�<N�@�B�@=��9���<+P<��<�5�q�߼={i9�����p~=o	E=u�ܼb=�Yy����;a�<�‼/S��.��~%̼.'Y���Q=�Ä=(DI=�I'�k�����a+d�~�;Q�K�P�N=&ټlc%�3��<�����e=��.=�=����NV��J�ө��[�5�=�3�;�A���<��%=6_}�Wo�<C =�FJ=����51��=����_= �s�~ć�]m�<@j�<��s=��n=����/J�x��NI�����P��<���<�䲻$bb=+s��ٙ;/$���!�g�=��R�G</<���C�Ȼ4��=r^w��7�A�=��H��~2=e�<2JF�!��<mL�<�;ei&=S\�{K�����[P��p2=ԹO��.Լ�(g�;����:�����Ez�^�<r�~���<��=2��:-8�<��N=>��;.�!��<�3*=���
A��U}�<QkC�϶X=��<}6��G��WB��b�<3��<G�̼I:���<7}�: 2�_����<p�Ǽ��Ҽ���<�������<��0=ō����;�ؘ<���q)<�[P;|=��=��B��в;����t�<;�=�L ���/��'!�0N��&~p�9;:�->ڻ��E��S=i�i<�z\<b��fA�<���8�8D�b�,!;�x�<���<��ü�;ɼ��v=.��"�����:u���<����K9=��<b��<�o<��P&�[�<wo;��R=qGü5e��ۂ=w#7�H<<��:�(�<Z��<!�c<�O6=�z�<�d���YӼ%���5��6F=�_�6�����;�<�y=n�
� ��;I�-�44;'A��D����x�P�F�5=!���g!���<�����N�.�1���*=$x\=16y=Jr�< P��	D	=�Yɼ�r<E�U����ڡ�<>,p;�F=z�n�g����2=~aJ=q�ܼ&�(=_y<��=_'9�\Y7�u��=i$�6.��󏹆v�<hM���0*<ד5=%0&��u2=�n�<CB���<�i`=},���ٻ���/=�8ڻ�I{�N؍<��;<0����0<��=��HW2���2���<@�]���:<L�Y=��/�ĸE=�p@��D=~���&ۼFԘ�Q�:�{�<b�M=Z���*D=�\�#i�<�#=U�<�YG=�tT���c=O\�;�j@������g�bM�:�Ν���a= ��=��<х�<�����ڼei��`����"@=7�`����<����`��<�3=<-<I�T`</�H�c���z
�ԅ��t�;1��::7���<'�<�m���V�-;�O <BPC�>YK���<M	=��.<7�@��׼��"��V�=<�.8��4�9�=�=Z��\ݼ^!.<�� ��=>!Ƽ
�1�
|�x"�<�=Q��ԀO�	�����q�?�<<J<�<��sC�:�9=H���=wL��z�<D��<q��:/-H�&���oP�v"�=��%=/Q	�4~<`�E���Y=�v=�X���=]<��Ҍ=�8�<��=N�R����cy�<��D<B�X<��= ��H�X<���ه7<Iw ���<�26�~V�$~���=�=�ǳ<F�>�0�*<yڼ�nS;�겹�㨻��6�B3+:k��J�ڻ�A�:R�I��d�ғ�W8�<�,/�0m���;�R6<����N9�w,��ں�Xc�ǅD:�����^��?��@��<�r<=������&=<[R��s=�5�;<�<�ե���7<���<˿�a�
=
Cg<�
�iP�<�_B�A�!��������)�L�=�O��Q�<,�U���<$d�:�߻�'ǻ��<�}<�~=ڍ����=g��Ht!<R�<3��<�S�<O;s=	���ĥ��<��;=jg��)'�7�<q%�ۮ(�X��;�(�<s�G<2:=�}&�/:�Ɏ<=��_�����<�/����d
&��'=3g�;
O��"�D̡��k�=��ܜu�(�=�MA=��������^=U����y�7(!=��W=��=��<؃ =H�$��1z=ך;����k=��;�?=����3��b =��ɼ}�s��Њ< ����q=ՉP<��.=��	=6��<0.���I&=�=�塼�諼�C<�U'=��I�(J=��$�
܎�*a=�<To�<��C<Բ�<�P"�:ͺLw�NM���2<d+;�p��<{����<{�U��X칿⟼��ӻwD3=
�n�!�^=I�+�*��x�+�<xI���;��2���=�>�<_4��b,�ot2��oq<�[4=��<�)�;
%L���˼f�	=�}����:�Xļ�yϼq���)v���)=#�4=9j=�KD�0��U�d�r<�Bx�9&�9�n�Sn:<�R��A<��c=� ͼ�c=���8�N��z7�Nw�<ʧ��1��6D��V-���!=Eh+��茼~�C=�T='��X�;��� �T���AZ��^k�)�&��N=��r=	0Y=��:r��<����H=��<�Pᙼ�_�hD��߸=ނ��F��'W�ȇ <[�"��[=��v���R��J=�<d��[� =]3μdȕ<
B!���<�{ɼ�B��g4_<���<ς��Ҟ?<$���$���<E���1+�طb<���<��)�=mv^��ܪ<'~<�P��@͜<$@������=E�=�f<=r�.(/�H&3=�fZ�|0=ښ=����%�<=D�A��s�<Ymy��k��]�-=�]<�6�X4�;�%�b��H�<�˼�y���<n��`[���(�J�;n<|'�<�d
=�vp�vL<f��<��(=��<,r�j�=���<�k��ߛ<`�=2��<�����!=�dg���>=�û) ����<=`3<�棻�j=�	=p���O<{��;�ؼ�N�s��<�O<T=���<ʌ�iq�<;�b��J<�*a�%����F�����4O[<��"=�M��@���*���ٗ���<�?�<جU�="�$5����<���y�=Z_����(<����~;-�o�7=eD��`���� �W�ļ����N�9<p�/�h ���N<�T=<���6��=�̱<�0��G�;�x=K���j��:�<�,�:���<-�I���z<�<=@�B���ڼWm=��<͹A=ޏ0=�!0<�2���<w;� �J"�<P������[����`�=^;�8E<�%�;�H<Q
)=5�<�݄:=P�<�Y=�V�],;�2��58��=c=�iR�i�.=�Cp=�)/��C<��*�iIT=��(=�E�<�mͼ�/=�,I=�W��㑼]�!�.��=��V�!$�<�Q,:�u޼qYܼ%}�<��<��໵C�"ûfW2�l�B=$֥;��^=B\=���:�(�<2��Wqc�=»E��<�M:���E<�K$�s �80�ͻ�G�X>�3=�5�=��'= L˻�0<�qJ��l��r��o:�<y�^��&�<�������3��W^�<k�S=�a%��F�<�$=�Ӽ[����h6<K�!<$m���鎼�c;���Ӽ�?F=E=��0�1�<��m<�~=�8 �Ly$=e�]=�߁<��#�rP�C�=2|��T���(��&���=�9��<�+�<��<�'�<^}&=��/����<۞�<!��<�F�<���;��=�q�;ub=�����У�#����X=��z�o�/��뼃}溦�B=V�ټ �0��D���h���y�Ie�:�s=�e�������'�E�a=����k=�3�9��	=�����=>�J���w<�R=X;���>���|���K=m�<*�9�y[(=c^�A��<}���]S��U�c�d���P=t$=��`��X<K-����i#4��0�<��<��&=q�l= a�<�P�v0�����<�;�1c<�����W� ;��Mڄ���<wl;�rN=�X�U�/=��㼕c0<���h�%=�;9�]h��i>=֤�<���<��	�=re<>�=Y�'=�`��8T�m��<$�l�L�I��9d<�:	=2����}�l,)�>e<�>�<�(b=�U��8o=�;t�`��n=Q,E�u�ü-��<�D���F�<*ŧ<^���K�R�Fx>=�Ѐ���&<�A=���x!i�W��cHR�K�4���s ��1<�uY�'��l���f�&�}�==S�5;S�`�s�����<v���x���"���.�翫<~f[=��<E��;�'d=Րu��~>=ܚ�_�L�K�V��#�:=@H'�{�3=+����<t%=�!�X�+�c��rv_=�K��K�;�8D=��9P>L<@(= �<��A=V���,%=M47=�y<WB�2��U;Q=�󃻂�8=S|м0�5=5Pn� ?j=�qp=)�ü��廿�4���Z���S���6<	p�<o[0��D=��=�&=FW�<]켃IJ�m�"|2;�l=���+=&�P��6)=ǘ=�w�;�a;���Ӽ�}���CŻ��Y�m�<l1O=�
ɼ��?=�1=U�9��F=}	���R=q]��><�t\���<����!<���]rV=�1�K<TDR=h�\�`�2=�</=�]K=�p�<��=~�R=*bj��˂;���fD�<��
<N�����_<l9�-a��<�S=�~���������|af�~V��U��z�T�q�X�bWD=?X=(��Fd����'�P��-=���<�~=�^�<Pw�=I�<i�S=�Az=�?<�+�<"�H<��39c,v�n(=���V�s�����e�@�<~8�<�-�M;��Dc=S.�;��7<��q�5=��J=�*��F=�,ļ�Y�� =�#�:�}l��G���G���<b�O�ִ���X=�~u<�m���{_=�DF��m���<T*x=�P�<h�ż�k�;�=Wٻ�Y0��;dh���:��t���U9�����B���4�<j:�;�l�.���b=��6=:�����+���`��"�<��f=g"g=��l=9�<�aA=�KV=R�=rC�<�C�;0.�0<=1\=<�N=�=�Ǉ���7����<���Ҿ��t�<߇\=��<��@�)C��|��<@_���
#<A_%�K_'=+3<e�:<��'=�'ϼs/=莼��2=f�^�s=`=�&���Bü�i�<��O=���N�]=�|��yk�R�=��7=�~�;�y��"�<�Np=Y������TA;��,���<!��<�ݍ<��7=��W�.X׼ ��<P��M����Uq�%�ۻ�w�j?����ܰ����kn%��c���P=����y=���<��C<�E=6�;=S�G= ����e¼���<�۽7���v�%�=0����qw<U����R���7i<i@�r&�=� J<Pν��x=11������ż4_e=�� <��� C��7�(����`'�m�|���O�}=��)��+w��!��!�<��4=+\�:e���� =i񀼲�V�Z�W<�"��$ֈ;�ҼT�a����<�ွd��XJP=�DV�Ҿ�=�4�PI�;��8��;�a=�7�Q�;��� �<q@���G=`>�A���G\G=[��ט�<	���樻�ְ��t<���W�4�Bas=�5��A�_��:X=��<G�I�V��<�A�;���<I�:a��<rD*=��H=�fl<ŎZ��� �<�z�<�S��Tǐ<�� =��¼@�[��"U�!?�<��c<!zD=��G�8���U�$>;��;�k�`�<��=-��<�`=�C�V�ӹ�ϻQX=�S�F
=���C�M=�/żIs�;�=9�!=J�»�*<k���z=��=��"L��<��Sb<	�ļך��陇�o�
��%�)<=0.�jF�=!u�<�\Q���\=�䁺�E�=���<��RX���7=�&��8O�<WƼT�=�QU����;��gDW��)t=S�=%l�.
=0/q��ב<��Q==��&=t�<��U����Z�=��==j�=��L�<vM��N=k>=\��<3���=�a<Dd3=�T6="���JWؼ�N=!	�Wz�� e���=+LG�b�,�� J��W���8=���f��;�\�;v�'=��W= $=J�Z��3��x�;n�,����:�]��%q��[i�D�<TO��e+]=������)u'��� �<L=�K_�����y=�(=	��;�HC��hU��i�;V4=�}�tm0��L�<{�<��A=�`�0ݜ;8�û�&���2���Q<:�-Zi<9eX����j\�l��cm����k:����<?#�ʤ�<�6t=�ZK���X��[�	,�a�i�u�<�q���kgܺ:��<� ���<i�q��m�l��	푼z�ļ,�T���	+��O=��>��w������'$9�4�@=��<��o=AnO=8�켻�8����<ނ=qiy<�#�<���:V#�<�<=��`<���>uw�6���!�T�DK��hf���4=)�F=`�<�C=�t������a#�<���K='=G�9e�;F�0=�]=E��}xV��t�f=�4s=x�!� �<��T=��w=���~�i����ͼ��q=6�S�M����gQ:=j6�D�=���<� ��!�<��C�mhr�y#n�Sџ<�o�\<ӑۼ)|i���m�ݻ��3h��u=RJ1��Y%���<�) �ho�<�r�<���<|<�)&=\؁���T<tL=w�=2	�<�6:�=&w��*��c���,��<�-`= �=.�=��Ǽ ���F�VV=IW���=�f���e����a�<�l�;����j��&�X���<��W<�,��μC���b=�fn��D=f��<t=�e
=���4m�<����L� *üDV�;�bm������xA<��=7��=ea�=-����ߵ��F7=7�}�W<�	=I�;4=�r<:����<=�<4��:�7�o�<�?�;f��<��%<c=i�/�u��:�*8� �=;�+1=�j�<G�<�h�<�G�<!-=���;��=��3=<.��߈<z� ��)+�c�O=(r��|�m�,�����Q��<�c+��xʼl�A�I
=�G�<k����+<��K�]�=�q=�P5<�(�������9�����
����������Zʗ��3s=<�#=
=ݣʼCq<�v��=�-<l�)< �<5�1=$�G<ϋD<��=N3��Fv1���4=:�=�r<�3x<%���;o��q�<��F�7�o�.Ӛ�y����<z_�aO�<`ہ<�V_<��<1�o��k��|<	�`�&=�q�5_�<۴.��@�ՠ�(���[���<�p=?�S=^�Q=�}�=Z:�<Q�¼L��<m]0���ݼ� =�⦼)*�<�7����;��Z���<b�a=��	=(%=v.<��e����6=�����<��9<r�B=��A=��=��v��0=�#T�[�����>�)=���o�n� ���X�<1�S�;<�P���k��:35����7�L{��b*�jW+<m.<�Y�Ux=�oL=�Uu= ���a��ԗ<�"�r��=���v*T=�=�l=s���C��0�{�5�:?=#,x�s�$��"d=o �=�=�N�<�n�B��;�ƺ����2�=$r�;By��V��[��a��q1���A=�HG=�IN;��������Ӽ\g=z��9��ټ����A=�{&=�2|=�t��J�<ҥ�ϋ�;y)���<!�<���b�;�.=	���^����+�rV�� :x�V��f�|�<��@�*�<f�3��I�<�ە�=X�ߜ��Je��Cd��>����<+�;�d[<�w;�4<�cI<GOp��ߠ���3=��<0�=
���*�:<��2��&�=�\L��/�<Z=Jy-�N����= �l=�H��˻��.�;�<�@=����`=��?=	��<T�1=O�F;h�=�>�ǒ�<�w������
6�����ӍC����&��<7H2��[G�:N�<n�\��.=��Y=����,�麃�����	�:Ӕ=a< =��^��Y���=����<�(F�,`�<�A���D��@�!=݆:����<�<�[=�3��q]��)<��<��<v��<ջ��B/ռ��=����U�<b&���D<Ѽ蒿</:=��===2��;P�<NC^���a<%����2�j�0=��};���3=m�ź�є=�*ʼ��Q�D.ۼ��I@=�4��=@���JI ��ԁ=T����\��C�<��ɻ��j=��5�_��<���<'�����;n�"< ;���<R�,���M���L��ռ<&��*�_=�
�<oUּr$R�mL&=��l��G��x{1���x���=�cs<;�"�<��L=F�<鼐<���<.�\����j1^=�F��Q�Q=P��:ꨭ<��5<��+�u����_<��?��Ǽ7x�O�K����=>�B�m�<'�=�*_�Q;�����d��|�=I}b=ҟK���=ri��́�nQ���0<�qe�k5S��l��&;�e5�
:�<[�>��s�<��4��V><�=��o�|�<$�%� ������O=ɇ��E�H���B<�;�1�<,�<N�߼��F=�	=���'�נh=ӴD����;��K���6=,=＀K��^̘�'��;F�l��C<�g�;%���$�ϟ��d$=��G=C?�<=�����ؼ�$p=��%�OF{��#X�[��<��\��崼�P��m��	
��,��^��.F��<���;bf$=pP��l���B<�<P=��;{��<��\=�=�v=<��=	Er=eDܼ��:�����#�<�cm=�Id�Kn��>]�(��-��<uf�<m�<񀝻�(=�+�<�ר�7��<�;�<�)�G����=�!�-=��P<����	n�����ܯ$;d�:�d��T���n��<�5=���<��<���<5�<��p�<oB<�}=�N�B5Ļ80c�� 2�
Zʼ�
Z�(�U��.��H˼�
;��L%=T�;F�<g�<�(=�'<F�h�`��
���$=�=G=��3�+.|������׼��-=F���d�B���'<�)	=O+����;�]�;�*�7W���#��ļ4�D�B�R�[�����;���<�_4=O�Z���𻖮==eo<z_���q��r9<e`�;j��0E��֎<�A���j����9� ��B�:(M�6.�m��=ݐ2=�1=ߘ<L0��z�<�6<,�T1W����]�̼�gD=j�r�����[m=�Q?�0G�r�=o��<��O=��o=�ż9G�;f�A=���?=��=��X<,��<��Œ=��k���z<B�5<�A��i$=�>��`�V��c1�Y'��D?�����y�γ@�V�c<]�����<l=�K�<.V�z�<ȶ*=�(�����rH�%�<��=m�N��ͼ�"��)�< ��<>ϕ��(=۞w����G'G�:�;Vw,�u)F=>4�"9�<�^�<L˼.'����A�F!�<����'�;�`��2=��9�1��;�m�w�<c����И��bU=�^Z�<jl=��q�7my<>� �;Z��=p�$=�W=o�A��9��U�/Y$�[���of����u�k=�{�<��ƼJ=�g�<^��;=�X6�w^<���|=<�<2HP=�C=���*)�+i[<'Y��G=C=��S��Q�;5��<�����%�|��֨<�E���6���<,�b�8x.=Drb=nV�:�	=�#�e�<]AX��RJ=Ɍ�=�x3:��ҼË�QGV�R��XU=�>�<m�M��Y˼;Rݻs�`�|�=]C,�2(�=s	��W�aw1=��ؼ�,������g��9=v����4B=�Z=�UX= �:�q����\��;<G����7M�̵���?�<�F=6�����=WQ �{��T=������G<Y��ݞ9��=�������<
�8=3��;6�==���v��	Q����<��i=S�����Ģ��B><��#��D�&�>������nB={�Z�(YI=g^g�w=�����ڇ!<�J=Xa�<	��<�-a=_[T�Eg��S9�y��;�P��9�<�T*=�\���(=�=��<�/=Kl=��
�e@�z:=�f*����m�3;Ŋ�=`\ຟE�7�]�+l;j?�<Ԃ=�H��۽3��m��������< aZ=�~¼�כּ�`)��$=��;�;�;q�0=C)j��Z��KX=���f�� L<�@��/J�<�E�<��켏�=1�F���`=E�����:<�`�#!=\t�<M�9;�L��V0�:�Y�l��\�ؼ�+�U��S���]�I�=po<_�9���Z=��E����J�<K��;i���6	T<<'���ƻ�
!��{�<��ɻp�0�EO��(����<��D�Q7����9\�<�;ʻIl=�㖻 
ϻ��m�bU��!X��<��Q{�<�jC�j��Ӡ��,�<o����L5�>�<� �<3{*=Į<��c<�$h�<~���=�=ck�עB�F�<��m�8<-<<d_=< .�$������Po<���<�5ɼ�A伆Żͪ6=�K3�
9;����C=�Y@=���A{�1[����S=�c�ɋ�;�,z�R-^=_G�<��<�?b���%�w|���v=3�8�3Z�<b�S���y��𰼐�l=��4�=�\=�gq<;�@�d.=��F<�~<�'9=G��2��ۘA=�+��'�<AP;�lU<T���l�<}d;��T��?�������R��@��[;~e9�,� ����S=o�#=�b��m[�C�<�Hp=�k�i����kJ4=���<u�E=\�h=�`;v�`=�}�<
I1<�R�<�Z�<M`�<$X�I�<�J�<��
cW=��9=��A=o�9<�H��e

���޼+3�0%&=�d�e�=��C=�D��H<�CV<B�H���<鿼?:�6{<G�;��z�r���j�:�<�<i4=�ޥ���<�aK=��=��1<�v���4�p4T<��R<��&�����=����������<��I��	�/p{�&/C<��<�Eh���̼eN�<�8&=�]T��X �qބ���t;K�,=�@&��`N�~�ɼ�8Y=Ld�;��<��=�Q�;�/@;p�/<A�:�&��X���;�\�<��弴�<����?��u#�75<��ż��ؼ����� �G��Iξ���t<3�<��=_)Z���ż}�<��"=��K=�m�<�6P�X���K�ջB3=A#H=�B�BO2=��(�i3G� �&�q<�֠<3��=?:f<���a�<n�=�6d�]� =��>=�g<��=* M�"2H��ƛ<��'���=��<��<<'=9
�ms!=�������<-l&�k�&=T�?<b��;��ü�NE=��=��<��Q�4��:5|U<�ƼR�5�uȮ;��<�D��9=]V�<m\�8�4�Mε�,i@�w,�< j��뎻f�)<� =��v��r=D-T<Zk,���/E=�A<�`�=�D8�\�@����&�\�oAF=�k8;�*���	�IE��خ^=�@��'���U=�M���򼮢"�گݼU�/=�hh;�vS��`=��P�4 <l5D=}��<�G�<d&��6M=���H�)=��4=�x����=���<���<`��<9f�&�\='�<��.��`p�ڂx��0=�<|0,���f��뎻�@��9+<��<�� =p��<���;P�+K=�y���1=�G��=�mG<" <ڻ�:��<�%�8��4=��:��3=�=(i$=n(3�eT=lDԻ��q��a=�2��`<��9�o����<z\�<'�N=k�X9�Sy��=7>�\�)=�%�E̝�-�+�X/=U!�<��
�(�F�Ӧ2��Y=���<��9�F;�;�J<=R­��=��p�� �$=�q�<>�=����</�i�F=�*=
��<�-��ӹG;72˼{o� ��z}=�&=��<���<;l<~-=��{���X=hc'��X=�A�YiC��Y���K��fX<�Ү;�Q,��p<��^��� ��\"�̙.=�C�<�k!=N�=F�<]���t�P<�^��.=�M=����������<��k=u�A�<=�o��5"h=��;䂾;�(�>
J�z��(�'���k=�림jx=�P�N8�<�X��*^�0i!��M�<�s�<���<L}^=+�<��ۂѼ_&=�8��$<�?�q�=�=,=����'8��6=�밼m�<��@=@�ۼ�p��w�`�>=r�/�]Қ�Y%�,]���軮AI=�A�nD�)ec=�U�<A���J����c��U�:aW��.�<l��8�;�@T<3ez=�}޼����E�M7���;����I=�~?<��<=���<����՝���}mb<�$����W:#��;�Fa���n<4�i=#1�;��HU=��A=Vy.<��D='8�<��=��T��w�\��<[�K�3@�v�����}�����:Z��;}�$<�3i�ŒD=�>¼�m�<��H���=`�6�n��^�<�8ȇC����`>p<�bE;�+B���M�E����ŧ<�̙����=Y��<�1�<� ���d�<��d=q���;'=P��󸕼����(��C�<t��<ĩU=�1���RC=D�9��}���==�,C����������<dvI=��F</�<���<!�	<��B�ݴW=%"�;�2���ֻ�c=�H�<2j�<�D�M�5='dt�!^`���?;��"�����L<<t`��\�����B�M=$P���R=��C=y=��(�+;�,0���2��D�<ya
��3�^?=цV= ;q�?�O�<(�_��L2=����0=�&�<�7=�㋻\�籃<���<�S��%�<���<�@+�N� =�IԻ{��RY�<�|��G=QAP=DI	=O58�Q9���!�:����RQ��/G=h�k�)��.�-=���0c�-P�<��߻�s<疻�"=�	����#���b9�l�;�`�?b=��/��7̼�"E��F�����<�S�=DF	�v 2���C=|����1��B��J���9>b��sJ��`y�'�=ZT�3j�<'���<�d�����[��c�#=�����=��4=��<�<z���VN� ���B��[�<l��<�%<.0S�E��=�'�<�'��?�}�#=mPc�[=-��<���:�kM=�;�4W%=��=^��<u�P�Q+�9�o=4�
�\�=�,=�|=�ގ<���<J<��d=��_���%��U�<�e�<�=h!��� ��YTR�T�B��+f=^[=�����<Q�U=��&��<T��;��������=�1O:?�h�nڧ<f*<>3cX�+�<%ˋ�LS��?c�=�ʈ�+̠;��[�B�MwC���0=��=�X��4�N<hOp�|H�P�_=B����D��JܼCU�<��4=�:g<.�r���	=���<��a?��=9H1��i=��<N��;��"�"�#=�X��ջ��_=o�<$�c<���~��˖�A�L=NS��=��"�����l)��h
���ɼ�=q<�<τK="0v���k��8��U�<�9�YQ����q���Y=}7�<zW=���������;|<�`=Fm�:n�F<��$��`�<�d-=S�伥�=����4�����8��q=A��<��5��$�U��<ɭ"��W)=�)�^����<�;6H=�%<OC�}ۼ�@���_���:h腽n�%=-�*�iN.���}=T��m���B��P�Ł7=�� =V�<𣙻pV#���1� �Q�_���{��s����Q<!�Ҽ�\!��w9�	����;�>�:g�D������-.�6��<��=Y�<|�6<]�ֻ�1̼����l%=��-<��o<��=��i(=�|):��;`_�<6p�jF�<�z�_��:�t^<��Ҽ}z�<��=Mg#���%<:��na=���Pk.��C=����x=�L=}�L�]�Q��<��A=�h?���!=��J=�o==/pI=�=zB���pF=w�<�����;���:���<l�
=�t3<���;�:�<z�=�B�ys�;�+��L�����s=rG���8<7UD�9 �<9Ҽ���<�C��l\=�<�	�����C�Y�{=tU�<>=�&	�]��8CS��`����Q<�_m�������/�hB�W="nE�7�0�"d�<���ꀽ`d��9��tq=��/���&=H��;�:��Q�=T�N�6�=��g=&���jծ�r
���+���e<9e����J�����0�<�Ë=�'�<%�̻S�#<ޥf;��=ٙü�5�<��;�I�EѼ���=��2���k;|�;��<b�S=G.!��}�<F$���9=c;w<鉓<�� ���=�=��<�y$��Q:����Ǽuu<H�뼭l@<��,:=�y/�!�ǜ���=��~4gh�<<�J= $=Y�T=n��l�Ӽtr�<�L<�dO��U��7��
$=�a��� 	��Z��S�!<F(=<�헼�E�<����5�˼�T&�",f;s��< ּ�	���[F;�b5=(ga=PoO=v�V="=���DP=�ݽ<-K=F�gt�9�O�<�n��������M=0��<��9=��/:���m�$�����S�h=}V���-�wy�����死�~~�uWH=��<"�C�pg=���<��>�0$+���=�j(=�8�<���<�A��O���j1=F=��	�.�=�<
-���id=�/c=ܹ�����ށ��'�e�"�p���n=��w<�Q��1�M�ؼ61	���Q�Ub�S�g��<�K=B.6=oآ<M 8�/c�;̐ =�&��Ӽ�k뼼�6����<y��;L��nYq<�Eּ���<���<��=|�J��]+��Fm=����-��Mh�|��<x
'�4b�=�W�
�!��,=�j�i���I<d/$���Ud^�$���Ͼ�<]�4�:A�<�=�2=~)��C��ޞ�� c��粼O��<�� =�9˼,w�#�$=��{��l.���]��7��/���<*�H<�nH���*�9F��L9�wX�;�F=�=�����<��=81s=��N<��<Q;j�Д;E=���u�I�;^�üIۼ��<�Mʼ�[=Cj�d[ռ�	�sj<�5���<��M�S>��Y�<o=�*Z�<��<���ul=��F=!� ��4B<�/%��A�� +{<�}=��.���<�λ�4=e1S=�l�<$� �H�����%��sP=Q~��%���OV���_��G��t���_7��{=t�G��S$=Hm�*
��ِ��/�5���t�<oX=D�	��M=[�<�,�q��9� =��=�2L�4CI�ڮ��m;!4N�v�#���X�ǅE=�fq�j�@���y��)= <sZ�<=�O�SH��\6=n�%=k�q=���i�V=+b���h=��V�#L)� ��=�[W=��,��<D�@���I=��_���1�jfK<�6g=���<��<u�<�t��f�t=ۍ�X|==���Φ:����m!�@;�<�<(�g:���<$�<d���C�=��$=�S�;�8J=Cl�=��O=4�U<���u�X=�{Z=���<��=�#�<֫�;ÄK��9�<���<��.<�!>��Hj;�f�<��B<ϊ6<o�7=R�(��0i=Sv�=��¼��� �<?8W=Pq�<�����a���=ѵ�<��ɼ�lY�R�/�5=�yp�E�=c�<0X=�0�<�Ǽ��B=��>=���<+>v���<>�8=��C�Fv�:�!�)�3<��@�a�d=̉^��£:�H�=2\��Er<=��<�ҏ9�_���� ��^=PA�<d_&��=_	N={KӼ򘜼m��<b�8�䬛<�}d��L�Ѐ1�:�=D0�JL=t�<�tM=�v=̀=;솽=���м�Q=����x�;vr=�����{ =�e[=�m-�
^�;ԍN�W��<β���*<݂���ǼBi=J�����=�8=\Cc<=`=�v�<�4<��;�Z��L=������<����jj���g�:���<�I#=�GZ=zU����<��̢<\Ƽl^5=�7�;�=��;F"
���7���<[�2���D<ǶD��-n=��P�J�㼡�=Bk �<m=\(=��;YLD=���9�&=���<U�?=��.=\�Լ�N=(B=n�Ӽ�?���Z��=�=L�S�3F��R�:���ռWc�%G=xUr<PT:�-�N�4�@=�X=�g��Y�;ҝ����"=��K��='��<��e���(��o�<$fF��<5a�� Js=�@�.2=�q��8μ��<�-h���9<B<�h=*V�'2���<=*h)��5�<�����ɻ�p�;�j���zA��5<�n�<�#�<�W�<���<$9e=��=�fW�eʲ;7~J�ڒ���պ壄����C �L�9_R=Q�J�0=��=�-=�c<��6�+G����:��^��N�4�aW��W(K��L����<<���c2ʼ$�|����Vn�����=��<s��=3+a=0�&�6U=y�=Ǿ&�9�$Y�<�ּ=�5�� ������U����Sۼ��;�L��a8��z�?9�DO<�ż�|���4={v��Sʞ��L}��(;P�<�?=��J���ڼ��g��*��E�O=�b���Fɼ�����ڼlh=V�ѼSA=��񉑼�4i=��Ӽ8��NE�;q���8�<���;�t��*d�I�!=��8��<�IG<��{�I�<�v�=-~��x,N�O�?<���Y�U"�:�tb��޺<�ο��<�M�<���<mDA�=&��}��9�ͧ<�-�<C*�<�@�<W���&�<`�<]kn='���=��$=�,��X=H=C���'{8��<'�d� ݋<n�B<Z��$[:�6==;` �ѝ=��:1�:Ѭ1=���~~�����T�(���f6��L!=&(�^�伭�b�_X�<�9Z��AE��"�:�z=9�H<�O�<h�= ;<Ѓg=��=��$=���=� ��"�<�t]���N�<	�J��3�%��:�� �������^�����DE�I*=��Y='9��z��Q�^3�<��=n����l=�����fX��+�<���94m��P�X=��μE��� =�;�n<���;����kF<��P=e,��q��<���v��<Pa8�?G=@i<�>d���x���%=KN�<����a5μ�c����_��i� Cb;4�������S�;��;�5�<>�+=��;�E��zF��o��d2��M�A�O�eA�`�,����F��G��侼1�nz��Dg�I�<l�S:��E<���:�[�߄W=GM=���є<a�S�0�B�TU)<���;�e�<+_ �*�=�	��) ;�1z��/<=�����j��\�< Q	�Y.=�_ؼ2�F��a�<��B=�(�@|,�ˀ=tU�<��0��/��a� wr:z�5=�*<�l=��� =��<E��W��<[�D	��d�L<�n;��n<��I���!� 枻��y<����=�T3=��z<�g=��h=p�����<䵋;z��<��	=�ad<?(����<���l�5�(�=�m�;���Y�"�*�Z=��L<���;�ƴ�aJ�<j�#=�V�<8�=���=.8M<�Ǽ�2<�SI;��[�FƊ���ۼ��	=ھ�<c��t��;��_�dj==��F=k<�r��=�����b��Ո;_%�$��׌��a�<S��G���&%=�<�<��<�D>�H���HQ]=*a]=x0=<�:���<�=^�.��H�=�"�曆<�vU�`���0=�Ȅ:��;���<К��?���n�<���<7���`w&��Z���,=���2y���/��$�<��<*-�<�<�e$�)�I�H�%�DnX<|+=��;�(�^�#=��;��<�m�<P�:�����<DTf�z�=~�?/Ǽ��	�A=,�	��:Ҽ��=0�P��\+=���;h��9;�1=��<Y56=���<.=~]���]�7�*�x��O`,=EB<Έ����̼/��=�K�r<���XQ�<�A-=C�m=02�;�
����~<��<���<l�7=�F-��l=xu�:
��;��<�o�7q9�H��;IR=������?���6�R#�#(��]?�8(��r�<D��;!>¼�Y=�z=��<�R0��i]=�Dn=b��<�tI<#'.=JZq��ty=�/����=�8�S�7;������;H�=�^�6O�<���_8¼:�<���(����Sȼ �=ո�<,�d�)=l���G�I='k��=	s��6B:=o2����3=h�!�?�=�w�<Z1�<aN;|�����G<3�N=ъ2���;��*<��=1Ȋ;���<�4T��@��<	�h���¼*�Z=jl)=	�J=���G�)=rY�������<�Ι�d/�=�ؐ���<�Z+���5.,=�ꂽ���<eU=�b��s=3�R=��.<Z�z�m����u��P��<�"��<�<�k��+	�-�;9)=�����-��<�'���:u�<.3d;����uR=~|6��;¼Do��+o&�Rv<5p=��<�����R�;�g��$/��!�<~�輓�p<e��:�ĻR��� ��Ϲ���:u'�<��ռ�(6���[=��4=$��<z�Z��'@��b�x�6���	=(��;U�=�r�>��b]���i=uE+=$���X��'�#&=g�;�d1<�P�cN���J=��5�����?0=��L����w4�\"D<auG�_��9�E�}?X<��>;�k����<��a<��z���ɼ�=��<Ԓ�<����oK�Lr-��V��;m.U��=`��=����H=t5&�0d��ń��$����*�;��I?\=U�c��ѯ��"<�U[<b�
=Mǧ<�=��<L����=1�W=�ʘ�0Ý<ʹ�;w�e=�v0=�N��3�e<��<�l=|%=˲��Y�=0,����<o�=��R<� 4= ����}��da<)P5��0���o�IQE���a����������9���z<���f<r;B=3�� Y�<(�0=�"$�����<�l�;S8<Ih=ͪ'�N)����3Y=��J���h��E=����a=��+�~+=���m) �z�Ҽ�:=@�7�`�!�Y=z�	=Gw���<fo�_��D�&��.�<�DV<C��� 8<+2�����<C��	=e*@���}=�	�/��<n���B�=�W<��@��_b�A��;#ړ��[�;�<���`�������L�_2=�S���[V�X�=�1H��ʼ�])=O� ���v��?:=�	��ϟ;�'�e2^=ƣ&=��l=���*t�<�8���ո<��P=�7�a�-��� ��`�|Y=)�>=�Լo��<I����H"�H軝/-�V�:���<c�;������<�@M=���<��˼�Ҽ:0������>�h���C�j*�<0c��嵻<��!=�ú�+O=,�%=��"�t	�<���:�
��p��:�t�k�B�&� @U<�P��~���üy� =�����lb�2%�;�"�It>�A^B�s���~�M�����v�I�+Y=�B=���<�4;�~2=)Ҽ�=ʸ'�f'�=�L<5��K��<��=#���2;f(���<�R��d&3�V�G��|�;�ֿ����<�(0=[4=���<7²�W���V�7�E��㩼q���Dۼ1$<�lM=���,�E=�鼾����0��T��+=�j�D�-C=���<��m�/^<ɋƼ>��G` �%��<�x2��=$�=.�\ ������<;<9<�O=0?[=|7�G���p��xD=�.���U=�J�nػ;Zn+=Z�y��:E�<�eE=O�<^�D=Og=T�<
��:s�D=18<�jA=_���X6u<$=ۙ��}ݼ#�(=�%m;��d�"*<ԡ<;�������<�<�ׯ;�'�<NvZ=X<<��<*6b<�[g��c=+�P=�))���<�6+=�D�<RuJ=��f=��=D�0<�Ҿ��ѻ<Wb�;�ĩ�&m�:�ڼ$B����<�<2�Ȼ�q=�����8�t���[i�{��VnI�=*=b�%=��<q�=�?=hm=���<�˧<<+J=���<(k�<��Һs��Fݼ�<�{d=���<�N���jB=L�m�:1��ns<L�B���<���<�d����ֽ�iՄ<e(�7�-��xS���o�ڇ=�E��������<�Df�v�=�������%�\�Z����<ԧ���uX=��#:�@!=����!��n�<��<\��6<��y��׼<Xe�<��;�ё���绦<���5�<A2�<�~6==B�<��<����(��r���ɕW<�ֈ<y�<�(��
;�D�;5M"<Q1l��8=A��8�l�<S�);
DR=}dY:�lN���w<�mB=�(����P������T�>K��/��@R:�
H�;>R�<u�<=����v�S����ѻ��m<�
��%��CLW:Ѫ=\�N�Z`s;ǳu�匼�P@��{����"�k<��=<8=��$�J=�)@<�H�<���'a���w>=���;����λ�E=�N� �l<����s<��=5bP�v��ӗ<����T7��ZL=��L=�	=�L]=�[�<���Hü\��<}��C�=���& :�{�]=�[?=�g�<ֳ;}Ӽ���дv��M�;�><�T ���!;ON���9�@�D<�(=�(=Vq=oZ�9}H��i�<ba`;�j	�D�Ӽ�p$���=�<���]:�1H�9T��B�)=y�$Ƽ;�K��۩�P�;ѱ�<E}���K����=Gi=I�D���0����Z�5��b=�\6=f�"��==�AF����%t=F��dz�;��=߀�9�_�(����;�����D<_�<̙G=O4�<{=��^<<~��X�R=(��	�!=�Y��rm.���S���;l�E=Y�=���<�{(�A덺�!�<�����c=	H=�f�z?̼��Z��^=�[w:[|<4���G���P�_%��漽��<HP�<-�B;#�<�	K�d-�<�セ�g<��¼]��<GJ���T��<�;�9��
��X���@=)w=nA$=�f=?�<Zi�<,�z;��b=p�(҂;�0=1ղ<��H��,�;\�>��x�1^�-G�ҳ�<]�N��\=�_?<cN=��<�#����;h�S��#l�Q�2����39n�φ��N�;��Y=�>=��<�J6�I>=;Լr�׼߶f=ɨ5��=?=N�b=��<}2=2^C�_�<�7=��	=�H��N=��i��OV��J�A��<{�_�Xg�#�Z���¼���P<&= ��C��-M=��a���T=K6C=��<�[=�<���<��#<-�<2�H=��:<[�+���D=_D/�Y�����4=T���8�:�Y����)��>����!=JE�;��m�0��G��e�����(�Q�I=-�,�VG=0Q=*��<mpn=�(�<DpH���T�����0d���I<3؄�'��}�Y�h�K�蔂=T���o=�D=.__�J�.�0���H�f9)�i����p*=\&=m�9)���6�=P�<�K��y���_���=Cd��ic<�������(�?�{=a0=��m�5��iM��CFb=��<\N=R��KSM��삽��0=l�H�cb�<�'�|�輭�7=�ET�*��6@:!�{���k�.�޼��˺����
q;���<"���%=F��<U*���!��&_�<����nF����;&&�<�m�<�C��Z���g=:3̼D�l�g�&U��"�l����vd���5���*=��
=�I�<CD�<	��<e�ټU</=f3^��-��0�o=*����<#q'��=�g�i�ຠT�<	н����<@?B����<_�������@���n��
���<��4�r;H=�=�eM��%�;�r��H|=L;;���<'�a�Ā@�ڢ =6P���;�� <��l�� =�d=�<pC�\\'��N��=���4k�+ܼ�'8=}��<��=/Em=�	I��8Y�
C��N+<�һk73=��Z��*��g�<ʷ<��y�/q����<�E=�Bû+d1=z
�<�N;<���<�(�e~�<���EP=��*=�k=0s�j��<^b��W�	2��<k�Q=
�S��Q�Q!ڼ#�<��=�e�<�05��S$�9�@:�F'=��<��V��y��<�6=j��<O��
�߻�b�����y�@��N�2��N�.��\=�u=W��*wU��w�On�<�ϻg`��+ü`�E=K/���4���I�#�:@/1�ͮQ��Q=�G����;��j=��1� �����"=4O=�%��5������<C��N�μn�=�=��G<z�4������;{��<��;�p=�K:��]�Ӄ��1�<=00�·[=:�=$t�<�]<�I���9&<%�,��?<�3=IS<<�<�V�>M���:�=V= �T�W1���=x"�ʙ��r^�c�<S�<jݞ��q�i��>B�e��<mB��
���d)<��<����q�_Y�;��<�N=dy�;eVA����<;����T���M��)i<��<�4�<J}n�A<�Ҽͳ(�4�=�=׭<)Gr=��Kc�	A=�tG=��<)���R���TD=9��<�X�<�+G�+</U�<rs=H��}R�;�O�<э�<,�;`^��G=:]�R`=�����U�[E �Lλrߘ���4=��C��Ƅ:D�E���<�b<0.�<H}���غR5<LkL��Q={����2�����])=Fᅽ8Cy<�i�<�L=Lx����=[�<�/e<Ϋ����;��ϝܼk��>�~<�?��A<o&M��(��ث�T+��8�50|<l�x<�͔<fJ$=(�M=�㞼߫=��g�zD��K�|�<�`���hk�ǁ����/���5=�Nh=`-R�*;P=�����5���{J2=��/=�`�<��<�U�Q������h��<f��{B3=H�g=��</nN=�����μ�-�=��T��
�<:��<�"=�#�(r=�@V�\�A=����B=�6�:$�<�@����U��S�8�e�U��ڼ��(g��h��:�\س���W����wV�<`u>=�[��=~u<��ަ��Լ?V��#��<d��=��B�l�A����;��0�s=Nؼ����2��	F�<T�<bE����3�)�.�w�[��G=F�[=�@h=��G���`=5m=s�}���;�?ɘ��D=��=���<�K�=�c�;be1�K3�ڈ�<;��<�7p<�~=T��=��<�<��8��ټ�U=��]="<H=��$�)��u��Hg���
����:�L�<�=����&�=�|'�(a=5����G=UB=��t=|��m^�<� =�N�<���<��W=��=�=jț<�8��\�i<G�g=�@�&�Y���b�w=��t�"==	����Ըx��C;����<S�=ہ���<�.P=9���#��<�%�<!q�<�[���|��+�;=^v�psL=�D��MZ4���G�w=��D<!%�<Ь=�����Kջfm~<�`=H�<i>=�P�i�!�����*�� �� [=�C=*=�	�<f=ӱ'�@�����7��M�<[�/��!=/b���.�R�G����Ct��D�=�=��n��ؖ<�,=Q���m<��;�UT=|'!�I^={}�<A��<��Ҽ_��<��B<�����;����한�i<��M=>f=?�U���?�ٴ$����Ep��'�<�`ɼB�s=�绻%D<{u��a+��أ��~�<v�J�� ��"s=��=��N����>�6=P�F<Ч#=�������<l`}=q/м�(���+�NI=¡t����ٞ*=4J=k����<ƪ4=�?=���<�W޻bp�<���<v�X=ήe=�h���d=j�Y�E(�<��N�P_V��\�v���?������<X���=��=D�<�{S��t��f�;L�=�I�;����6��LD=����f�����=z,�HCd�m�u=��<�"�e�ͼ؍<(��<���=��q�����]� ��O���]���=��<���<�==QL����<I�J����;rr���]:�7	;�\	<�8&�_�5�Y��<jF��KW�ێ�<T8�<�O(�(�K=	]=n����=N��=P��"�����<�[=8��<j`�4�"=~{C=�\=\l?�8p�<R���3<��ǻS�<i�n�ԬQ=k=���<�=�/����~=8�]�HS�<3'�<�� <O�<ѥ�<��<�#���t�W^�g�T=��=͹��GJ=�=<fOM����9ZS �q�h�j����<6�@���F=�AD<�{��͸<Eم�n�5=2q��ZO�R�u�X�=q�����;6���}�:��=��ּ��2���4;�Z5�Y=�����L�;��y��>�=<�;�7=ʑy=t�<�%l��g���<,��;�j�W��<�Q=�ar�?��< iO��q*=!�=�j\}<\���
����+?"=��O�����l��u�<�wm=�9=B����4.������|=;8;��O�E�1<I[l;��<��<�e��i���9����(��<%wN=O�=fJ��� ���L=�(��U_=�\c=h�:�aj��F<�?���߼��5=�];=�E�<��E�Ƌ���p=�+`=G�,���l=���<$t�=��3=N-d=��<��'���=��׻6�l���=�û���g~�����<�}�8z��FJF���-=(��U<�,B��4�_�O�fPc�2�a<�8�;ӈ=�=�kH�q� ��wD���=J�E���1��<ʵػ���<ô<�{�<����/�i���V=��=��&=8�=��^;�j=YfD=y�<V!X=|�F��z�p�0�v�<@�#�迌�;s<я(�ՎN���d<4%=�񶼽��A�'<K{4��|9=���<�+������Y��р���=,ۭ� �I�@��=m�B��C=�
���ҡ;�K)��c�<��;���$�T8c���<�=�,x��Cü;�~���h=�=%����]��a��b<HH;<�&=�]�;Û;��X;�3��g�:�Ǽu(=�@a<�#�<7Ϝ�;b�f��Ņ��l+��*t����=/}�@L}<��*����<A�x���S�e�^�lg����߼�]=�yJ=�7���Z�!�y<�dW;�HF=�������<����h<Z=��<�L)<n�<�d�K>=x]�;���<&.�4��hAN�� L=�z����<��1=�t��y��<�;K=HI<��`=c q�0a���"=�3�6�<�j����v���XY�K����-��V=4ܼ�(=��&��^���qQ=p��<(����ż����5�;kn�='�6�ӂ<���;��<2�=���:�==4���<Ӵ=+Pc�읟� "�<q2��x�^z���T�<�)t<��伕�S����w�'=�O�<J�q<[���V:����<�3=�<�B7=��<�]\�Y8T��k�<ŀ=�7=LL�<L��<�6�^o,=Ռ?�Ɍ.=�?����<8�	<X*��@=�?K<}��;`=�û;�!�)& <}#�<=g;���;vf�<a=�l7=�f/=������1:q�;s�=�W����K�3�T�@�5=��<��H=\C:J��<+u�;;��<��C>%=��<�Ѫ/�E �O�����_<W=Z+T=]�Z=D��9�r���3�����Jѕ�B�����<w�x<�+K=
�H<�H=z�K=��<�=_=O*�R�ڝ<���d!�N��O�&=��Z=�|�<��<�ws=k�=�+�;�&Ӽ�8�K=�m=��<157=�'����<����L�<��h����5R�p*/=��=���<�W�<�b��t=9B��i(���M�۳���U=��<G�=a����q;9	���nZ;k��<�k�4�6�JbZ=�M�V=��ռͅ<��:#�m=8=J�<n��:�7����=h����=?(�?)�U���Ĝc��\�VV��;��<\����,n<�����l�W�e=)oF=X�<]����]���̼�7Q=�+;����=�0`=I]�<l5=�t�<�(��&==S=mi=!�5=lk�<�[���:��<���;A�={h=�k9�83����:� =�36��<| ?��1�v��<����j����6=j�6��K�<u#�=���;@�=��[<)�Y=�n��,�=��vm��T���l�v;�ż�}üj��/�N=DZ6=c<ER�l���ß=iO=��+=	�ż>�3=A��H-;�(=5��<��T<S��Q��x]��D�<���C��<ҿ<�Q�;��M��V=j�a=�X�'�+��'�:��,<f\H=�H)�� q="��<E��<��Ea���x=�޵���������`=˂>�mSS���=�5��PF=j�J<��;/{%<5�U�|�d�_g���<�=�l�۔��O�v<=ŵ�q��6��ϧ�=���<㝼����<
�9��ZK=�=nܺWxx<K=���<�����wڼaV��[*=ì;�=0=��<�.<��P=/�=D	9=y%�<�;Q�\E�B�;�K"��������<��=m�=p1�<��c���D=�18��X:=��:�G�<nqA=��n�j�\���k��N�ʽ>��s��1����=�U�2H=�:={L=��[��;�H7=UR�<Í�%��H���$; �d:��P����<�M��D�T=Z�лG�s<��N=u2.=Ϳ�<���:�,��ft<�{=�i<�L�<С;d���k8�����+l=��0�X1��T�Yp�<Y.ټo9�<5ܠ���w<l�_=j\�j1Q<D�:=q?�/����k���M���L=q�K=P|�<X1&�������;��=@V��2�<���<0�=��/��ц��i��;��<�=d�i��e=n�:=��;K����Tb����<M�#<>��<��<��4��Ջ=��;��^�(;�����c��<�恽�);~E= �ٻje:�$�/��oq���#�1�P;�M�}��<3�=��<m�M���d��x=�m=�짼!/�1�7=� Ի����-uK<���\Y�;WU�;/�<}�G=�' �
ou<J�w��TJ=�G$��;=����<B�?<�=̬���K�]�*=-c�<p�[����?<�.2<�4=�N���������=�y=�K;�n�=&j.<��=���=H�w�y<�����8ƻ�S=�p1���=;O"T=�K��p<ߦw:�,�	�C=��<sy{=$�=8�,=�%"=��C���$��sH�����{��V��<b�L���%�Ӆq���<�c����M=�Hk�I�4��x��j�6��»����UM=�z=��:��_\=?n�<;��Ţ��^���ռ��[�\<0_��5�:چ�<��B�R��<��I=K�˼��P=��9����r�U�(�<�`}=��}<��V=;�<�1ۼN.=蔋���_����'��# �uJ�;@�1��G�=n��<��0=�`����)=r����SѼ���;ȡ��6�*�<fc5<�-=HCO=c^��)5G����BԆ;^aʼ��o�_ݼqp��������4���A=ia��^�G�:b a=�vp=݃�������:���a<�N��8���<Q�;��p;�iʼ�L=�
�<,B�<�� ���<��P���4=&�ջldQ��5>=ң�<����	��17�<�1��R(;Bc�y�j��ͭ�Oo< n=��<�A�;��< �B�fl����
=��)=�Ƽy]�<��l;E�B��2w�c;H�~<r��� ��tX8;kO=h�<�~9��<�����fU=�p���]M�ٵ�*�G=�F�N�A��6M�����QC�o�ü�+H��&Y;;p]<@%�;NHI<O|�<1�<���=��v=��<R���d`�=�AD�Uļ�zm=��b�s"*��0M=wԫ<28���:=K<����e6=�P5=���<��'=����A���x�<=1G=-B�;Ym�b�<Y�`=Q c=|=��
����F4< �7=O8D=\M�D�$�6��<~G4�Z�R; b���h�<�b�!�3��.�<��?=�~�4�=x?��ۼ3A^=2����e=��ּ�.�<�I"=��=�R8�hj�<_�=��T=g4=jKD�e���7q��)�=�e�E3���=-��F�b�&���%=+�O�0�3=��
=:f���>p=z��<c�<խ%=C-<�
�]�[������e���̼�搼a�V<��h=������<�s=��<���<��[<F3R�U�8��h�<�&=.�i�b�S^�<�t�=�-� +Y�1'�<��H��?��0=b
2=��&���l�<�1���Z=P�$=?�����<���0Ʈ����C =L�Q=��ϻ�x?="�:F\o�z*==�o�!q`=���;�bǼ�C+=(P=�]L="�:��r��B�����	0>���-�aC��>�<U�ۼJQ���x�t�=�<<���Oļ�S��E0�ݰ���*=}�;Lj�U�t=����=\�<��E;�� �β��XF(<�/=-%;<˥!=�Ar��O!�����;[ ��U��o�<Ĭ��m��<0뒻;&�;û��S�s='QV��~�`c�҈��{��/:=mG��,�z	<=�䅼в�<��R��i�Θj���i��<N�u<1s1���a=�R=��I=��|�
_�9tb���=�"�;KY�<~����Nͼ���<���,�C=�-=�h:�~{;=����:��9=�6�,3�<�<`|�;�I��=�S�l��<�|Q=1ja=g���Sxu=/{�j����=Bo���d�H쬼o���]&w���"��d=)>����;�$�<e��< ���=�<߬�<h��<��E=ξ�;*�Q���9;]�e=�Ѽ$Ϸ<�d=V���vS뼬Q�Wb�����ORO=m���댖;T�C�l)��˻�4��=+��A=q��=�w���~P=\-E�|���I��<9�"=2�ؼ)}$����k_C��6/<0�<�����:����}Q��G�=�t2�:b ���n=�+=+@�a�(<*��e�<��n1=sC����Ź�b�=��<P�<��;ⱨ<_�<'�P=l4����]=l<=lM�<�p-<$u8<ɾ���B�<��<�z<�8���.D��<5 S�I��;a��;5K�<VO=���=�G��)]�=z���Z�<���<r�%=�/=�<�c��9�R?���=́���;R�im�mڈ�����p<F<I�c=����=�#%�u�:�T��μemQ<�"�<�Fʼ����a�s��E=�d�<	�I��]e=�&�<��S=;� �_�K��l+���y��XX���y<.p�;gs=f ��x�<&���'P=ÿ���`�j�!�ü$�/;��:<{@����C.=�i,��/w=ς��ñ����
=��+����<�(+�&P��4� ���=SR:���`�=��8�Z=x=� z���N���>��6[=���<���<��y������TL���=�C=�&�<o�9���=�H��<|\»�t:@N=$�-;:-	=�<󋥻K�={�K�չ�<�Q�_�����[=e�V�I��<�s���=q�T��<[��w�<$=�n�����7��.��9<��\��=���Vr�;K��k�]��fn<ζ��Y�,��;���f��A��i�;{Cz=)u-=�|Ҽ:-<<Fs	��V�< q��e����FѼ,; =�x<���ͼw|�<�>�<��D=�:+=x\�?pf="v(;�]<?=R<N	�=H��	�0���R��!=�)2��#�<�ݕ����MƝ=�+*:�*�=��һ->9=�����n����<�>�<�_�<،�<�$��L��I7���<��<h�=p�g�=�T��f<~!=:��;�=&mE�70/��n�<@q=����?3������H��`[=9Q}=�E=�"�B�
�QE-�g��*C*=�<�'���o�t��<���;��;q�����h<x�`��'�<�4`�ˑ⼨��<������F#o��FC=zA�<!*5=�B4��+��NN�Aa�;q�;��0=b-Z���M=��<�ِ������_���E��!'�<�.d=��$�:�Y���C<&	<E���s���L��Qr:�%��zBK��R<煚;�	�<`/��r�C�+=�"�3���g��C
=����AɼjVK����$=釯�{n»*O�Ǜ<��R����<ԨU=��<��_�>� �;<�P�2;=��l��<)ϊ<���</�j<1B����:���;{V⼐�x�����<Bq�r�����
��=��d����lz<�����hv��0=_�1� Z=��;�<'��<,����ż�����#~=j�V=ȍo��?|�¿�������,=�Q��+�<��#���*����,�bS)��>=��0��d<01G��EF�t��y�;��<��k:@�Y��� ;��b=^7<\�;�.=,��߆6���L�ѣ�<��&�a=���u�x=��<�x�l��<τV��4�������)���W<ʉR=?`=��y=���<|
�W��<ԩ��q<�g���4=A��<Q{��6r<�qN���{�&��&nf=�n�;fHh=t���s����ۼ�!=��u��o�������odA=��N�N�c=��1=��l<���lka�Kp=���-����<Э^��(=���=h,,=,��p2�<��#�iջ��]�}��<M$V��/�<��W=\|=D��<[1|���=�be��y�:�3��4%:=�kg�yI�;�.����A<���<�Š�-t<�zf����<�[�;�+W���p��Q�eQ�<2�xzv�#�����"g=���"T�<���y8�<x�w���E=`�4��Hw�j^ <�ܰ<jK0=�/��*���S�َ���Q=:3��)��zD��D��Ő�D<#�����2�Qe6���	��<;�ܱ�s�<s_=ϭ���+=R�*���<���YV<��z��o<^q�:��y�q�7��#t���`=�ջ$�d�'HL<y��<a�<��4<��H�j=R<O�=���fO=�y����9�Ѽa|V����B��;U@���##=�ș�,m���tɼ�=�=MP���<=�S�<ge׼�1����;���鼬揺�=��#<���j<�袼b��:���	.�<��<*�O�Xi���	=��D=OD�<�_&='��	�<���[q<3�+���<�_I=��	��<�	���:�<�0�<�����ռ�9=��ݼ����0��~==���^�YQ�<���O(9=��=��S�A*=f��<��ۼ!����'�9�+;,	�b+�<=J.<��h=&�2�z|�˒��B* �E����Z�{���Z]̼��ɼ��)��~�<�e�=��=�C=����J^�1.��H7м�~1=U=�_�%
�}kj�Ls��eR���=<�ʇ=��I��KA=B\�<@����<�UA��@<r�<o�)�hZ=:�J����t�@ ���A=G�=%L;)ݻ��_�x6�;}Ac=�C�<pK=g�=me}���c��?��8�#���uy<_Z=�X='{@=��$��vR����<�wL;(zY=�
���M<�Q"����<v'�=;�;f8��� ���%�9=���<�ڂ<�G=�i�;����Y=�Ə<�6�<��6=��ؼD)*�53M�
���;����>����*=�긻���&��rm%��hN�7P=�8=_��<ľ�<�9;=�AѼ���a��9ߺ�)L�y�=�5Z=
C�<%n�ٕ������C�W*Ǽ^���M~$��
��|{�q6Ժ��?��ʼ,�4=����Ϊ�����M �%'��e�S<i�&�������a�b�ʼ�U��Δ8=���<\�;<U�jtԻO�D�!F �	f��.J���/=�)D=�E<�n ��3��� �m�<0���PC���1���K	=C�=,N=G�=�<����G<�R��=�Vh��}��c�=�v�<	�9�=r=���<c��<�'=g�F�Y�=;}"���;&)���oT=G��<Upn�#%S���S�&�*���	��?o<����� ��% G���<���<�����5>���0�q3�����tL<��/�QD�<���<k��<Ju����<��N���f%@�%?=A�����ż�T�<��;�;��A�X6�;3g�����z��%M�<���<�	:�ʼ�n���ۼ�G:�?���o�:=��h��u��u≻y@D�{�A�]�����<x��<Nxv��JG=N�H���.�UnX=��}=r�g={��8t��=��<��|<�1(=��<}��לd��I<Yq�=T��-�Y=�L����<�(_=�H=�d�<�1=|l="f��B�� @�������G��ӻ-X�<�U��{M=���*9N=�I0��bU��ǔ;�<8)�<n�yDڼ>��<3�� 1߼Ћ�1�+�A��C�L�bd6��C&��
"=ȕ�<E��8E�#�W=.�<�-�<� N�sE��@�<\h =$��<���<�Xt;dw�<��W􏼾�d=KWZ=u޼{Hx=P=�+|���ɼ�+���&л��=q��<@� �:�>��B=,Ⲽ�o���7���;��f�"�j=
�t��:��/>�����I;6=��L����;�&��a=9ze<b̠�~��;�ʼ�t$�S&�:�#�� p��0d�㷈=@;2�	��ᶼ4	z��<t�;0-�;�A=�+�<f��;᱉<�d+=�/l<��Y=т;Nj�<e�z=�u�<oƼ�˼̏����r���t=��?�iW!����)M$��vf=-(���)��U�)2< H:�uYX�f����ϼP�ټ2�?=y�F=,>�<��ܼ�O�WV��gч�YzQ<���<
p=�?=Ǎ��T��<��N=;-���$=�ZL="+�:���Y�?�o0��m<e=a�,��`�;�O0���,��y%=]+s<H>߼�����5�<���;65�ڇ@<��/���g=��˼�H.��J�<����S�=��<�І=]���<����K�=���^�< �'=.%n��	�:�?=;� =�T��L�V�JH=my�<��"��>廴E&����<�c�(/o��6*�-�7=֢�	�e��z�cdo��H�:��#�3nE<�'7��V������SS=(���(W����[=>�	�;�n�+����@�����yJ=ԍ=�@���-=r���#U������@5<�e3=1��<a&���v�;=�6��M=�ܫ.<}B�֠�}y{<�I'=�N�<�����cB�a��ia��8�u�źʩy=��<*!���8�<,�c=)\��ǜ;�N6='�U���H���M=��<�<��=�y����<�5�=�V=�{T=UD9�Zd �����<h�U�@�<�	= Y��md��Ю�I�<���-A=�����'�^8=��<�#[�y4��� :=W=�4=-M]�q��ӓ�ն���;-����(��-3�e�����e�=�Wa=ɺ�<>,=C���6�-�B�YPR��
=����(^=�}.=1�?��A��Ou<����<gH1��~ʼw<TQ���к�%$=Pβ<�	�<��'��[�:���;C�ؼ9o<=��e�������<���U=ˑ<�"N�E�f=�1��WH1�y�ʼ��=�0��=A����<gh�-�x=$QC=^��<�y<=D�V���<���=D;��< ���Ӻٜ+=���3�Y�ɺ���Bz�U����?��

��=�i���_c=kˆ:O;<%��<r��<��/��=@�~�f'��4�Z	A�\�<�y����$��u=����=�p���:=�����: e=Q|�;U��?��<*��<��`�@GX;��J=���<�8�Q�w<���<�_=���1=�w��*k=e;��L8��E�=�14=Y�-�"N��䇼�E,=��˼���;M�= ި���<������]F���z�a�Y����2���<��Z�=Ma]�-���9���<�56�s�=��=c�%��tq=��弰��<��<�i=��P<�g�;�AF�9Z�C�]�{1=PN=��9�y���;���v=����^�\S����>�<�=B=D�=K�-�a��<+�#���A��-=��_�y������9��� ��,��fU<��<�4�<m��<�����<� 6=~lͼ�[ �-g=�Q˻�P����<m=`�=<Ki=|	�<��V�����F��(�=A����WN���[��bm��,�'<Q=bā��6F=0?=}���:��<-Ӫ<����Ⱥ��w=���<�	<�NI������l���\<^<���,��pc;�kG����<AJ
�� 
=NY�<Kv�lAD��<�#] ��ߤ��R{=�;6P�;�@<�ƃ=
Q���xؼ����,������fE�G3=V�����R��]y=%�t=,��<D���v�<�b�<��}hv<��S���=�˫�g�=[�J��(�=�h�<��N噽��������~X�>c=�ư��}�<�{f�u�7��-<�4#=-��$��<#��Z��2h=Gg�d��;�;Z���"�RcH��w�<��<��%=eܺ<f��<H��<�@@��,���̼�����^�<&��ZP=���<@2�<6�=s0;q�<���<~N�<�ɼػ1=�W�<v�b��F=��:n)�<��^=N��<v:4����^�=:�6$��f^�g0<l��Gj��-��3��Q <~c�<<X�<�k��=y<;�@�=�
=ҪY:﷼Fa3�6�%�1״�Z�k=6;=�6B<��/=�v��4�<�����7��Ai���=�}$=ɢ��S�<�t=��*�:��́�mO�<�E�:���<��B��I��1=��V�$�� �=���<5�a�I83��8���<k�ɼ�QN��;=�#<�,����<�Q#�Ԣ��h=���<��	<a�������'�WS=�J4=k$��������<�I�<��;��<��<�d>=���<�fǼ6� �-J=��@=�n����J�G��8���l#��Ø�����3F<E�f��;?������A��$�<�	Լ�Ψ��?��=��\=hP�<S�]�zD=�{"=���<�"4�6,%=�7=0>���	=��	��N9<����!��\�_=C�<����(Q�<�x�=��<zQ��L��e�<HOJ�(��=�qL=�,0=Yc=r^�������L�u==b�=�����<u��s:=���:�^=��<�V=�`�<;��<��k=z�L���<�v�<��P��_,=��ļ�9?!�=ED���m伏�<s|E����;���<��Vg�;r�V=�|�s��F=��=�g<�@�<>ѥ�������A=Lc�|�9<���5��<x𣼓܇;��b��=|�p#6I��8k;Q=�����/=�"��<O�e�ݰ��H��:�.������><�2g���y�.G;#b�;�ϲ��<<=�|��s�^r����e����<8N.�7
n�@�7�������;"b<�4����<����u��P=}�/��,C=��$�ꓚ<I��j=����8�<W=� L����ū�<E�;�J�<<|��3!�<�R�!<��n=��/;���o=-Ҕ<�WL�G�B�2N�<Lr���2��p'�5�k<��v-�o@.=���<V,�<���-q=�6<�h~�8��D���f};>���.W=�ox;�K=$pH=��<u��'=Hu�ڷ�<Az���L=�=@�^�<=\���<9�=�Z��C�:��ڤ���a<���R�	=���<���;��%=�^;��v<�c8=�%�<�} =�k<�Ŭ<~�r��+=��=�~4=��;��2��s�=p~#�گF��Έ<8�O�"uv<�i�<�Y�<�3�|�м٨���!=`�N��==lnQ<-Q�<��*=�=�<1Ľ;L5<��'=��8�nO�;D�h=��:=���<�b��l=����uE�;[�;��A���N��Ts<l�<2	��I��>P=�j�<��c<8D<w������6����!<fZ�<�#�;�M�;C<���<��Z=��<�=ȥ'�vp��'���l��m	�+?i=$oB���=��<J�_����vs<����_�j=�!J<�!��W�5�h1=�hF��x9��P�$`��n
=��x���<�_�;e�\� &m=��)=�_=0�g�����=�N�T;B<��y�;n&Q=i=�d�=��<db;�V�<2s�<��!=�"=@K;=��h�c�<�D=@�e�/����*n=�|X=�둼���;���<���S3<�N=�ɿ�qs��� �ON!=Jx�٣�=���.=NJ�<����,\�t�J�p����H�}Tm<�b`�m|���=𙢼�m�<?�ϼ'��;�E�<՚�:����o:����~-�X,�=�Q=��8�`���0�;�Fl��l���ܮ<��~<�PM=�9�w|�kX��;9��s�(>����-��L�<7�#=P�ؼl:#޼R �<8'�<f�};S�<�&��=��=�V2�bջ�e�<R�w=��f=(�"=�u�;�|���/����J;	Xi<�9<�o�̼Jd��i<��):~�9�i;��=J?=���<���<{z!��.1�n�=�x�2��w<҂n<
z,��~`<aε�f��;��;'�s<6�w<�bs=��=Dki<��¼{�4����<1��a�<d ,��y� ��<��_��<>�!<��<��9=��f=��=���<�q��� �g<Y�f�C�S�W#>�r�]��ry==M<V��<�6=v�<x��������N�e=F>�<3/r=��8�L»����#��=�=��k�r�M�M��W���J�eJ�<?�"=i�\=I9H��}-�}�<#J��jJ���N��	{���&=~��x��j��<��F=����� �<��;���u��t�;���/�dт<-��<^y=�s�W�<�~ۺQq��~F�Ht�;E�<��b��*X���U�H7,��^;���<Ƒm���
<e����.��c��f�%<�T=���<fPP�+��P�<6���|(ܼc��.p���ټ7y <Yfa�H0��:��;�}�<`�Q<*3�<�1f=V~�<t(���Q=�Z�<r������GM�<
�G��d :.�2=4�;*hu��F�<L$`=e���|��=���𼇔�<(��	�(���^G��<j��n[��� =��:;8���= .�]����)�dџ<k��8���WB;�y%=
u�=n�)�|r�<�n�;\Y=6�~���]�~�;����<�1�<!>ļ�Tټ3�F��/�<��.;�����K�`&���!d���Xd���_��5=e���}���Լg�8=�H=�hj=�_ȼ��R߆<C�Ǽ�!�<�=��@y,=���<.-~�@��<��˼X�\�����.�s�c=�P�)	G��YC<V�A��$����<o��<@�S=�
����}��K�Y!>�=G=~_<޳��&ɋ�J�=�b<>g=�ʍ�qP�a����9<�9X��Y�:��e��jB��<j�ʹ1;�;�<�(�<���<(��;D���D<��<��r=�΄������m_=��引�yA�Yni=�� ���:��f�;Ӧ�8��?te�����?����<ln�<.�<2;�<�m@=Jah<�J=�C=+.�Q�4��E1���ݼo�n<-`Z�i�D<C�=E���K�<�S=f�<|�f=��Z===@<�z��<~{��5�������Ó�$5�1�o�"�	��=�}�7��:U�:�=�z��O+=㬑�, ���y<s=��c}T<�=�� 
S���< H&� �Z<E��<���[Q��0�Ǽ�ּD;�<�>8��GL=��޼ob�=��G�"}�=��B=yb��f=�Ѕ��g=kV"�ڬ1��;=	�ȼfR��z)=#߭<[V<l"��:�<�=���P7����=0Ԓ:}뿻���;���I�<��	<��[=覎;Vg�<�8��|�&����N�=&��aT����<�Q=���҂?=�Ov�:*�;��<zq׻ƣ=��n�-�2<��u=D�o=J�s�����$+=�R�<�����Y=�w=�	ɼ��D=�F5���g�뤕=�༘cB=����3��Љ��+=6�2��A�<T��<�� �a���$�<��=贐<iO<���G�=����p��YZ<��߻�Gi=��X��ɂ�ϥ=A�����<���S�7=#���T��<YD�<<�%F=�_��Vi� Y켜�F<��k�MP�ច�jTr�k�:6�Wkv��+<��N=nkR��c��*���uH�k�[�4�����A<4�j��}���g=��r<��U=�|�h�i�1�B��<>�6���$<CkҼv$�<=9=�sj��,�m���}�����\��(����a��7��k4����<��X��ͦ��m=�#,���޼������?=Y{0<�#I=H���5�;��=TYA=��5<��<�4=��� ���y��<*�����L���y<�XX=*��<]|��UT=s�j=��l<T�0;f�=eN��-�Ҽ�:=�P�R(&;Z�S;i��;f.�����<k_F<$������;2�<��ݻt$�N&��=A�N�)�=�=9���"g�`<Z��6����%�W[B�o��<2G={a�fD�;b�f<�+~=�~�;M������C4�~k�<�w<���mw�<cQ�Cҁ���"�Xb�<���x���#���;�|F��ût�<y�L� <R=��U��?=����=@�<�����0=$����i��$E�A~�~��<5�*=�(=Z�K<��k���s=Nca=#�;���F<Z.���=��=���f����� ���=J�!=z[�<ㄅ=5"F��G=�o��#Ż>_-=}�O�<~D�>��:�<�y�<;�<��7��
��ͨ�|&�<�<���L D<GK���-/=A=��τ�<�<�<�X�<e'<P�=�v*����<�e����=g�[=�׃��5<��/�>�b=��0��Y�<N���<K��ą��$<�/{<���<Uap<(�=ׂ@�� <��=X�μ���<]G�<��<�:*���������q5�;�%����<*����?�J�*�9@=fԡ�~����<=��O���=��<�G�<yG��o��O+S���<[B�<-/�<V���E��<^"='�<tA��7 �<���<��<�ǼA�ٞq<t���';C�?=i�=̼��<�wB=��ͼ�F�i#��gk���N����<���<����N�Cb=������"���c<�|�<g~|�*��^e=��9� �,=�!4=��e=��<��<RT����<�|�<6ZY=��6�N�<j=0�3��<UXs:`ı;w=�f=W�)�Ύ��i8�F���<��_=µt<NO�:hռUc˼���Z=�sm=Iһ�k�#=�{L����,ڕ<���<\I\�z��<�~�<����0=�0�iIX��~�:���<� ����_6Ѽ�μ�0�;Dr�<P�0=��'��;r�ˠD<�.�~�f��X��Z<"μ����kü�Bn=���;�3�;w==G�u<2�¼s"*�U=���9��P<��D�'zs�5�*��`�:�)�;NZ����;c=�H <�$=9$��*=N�;���:m&=������M���B�6���8M�<��<(��<��=�(A�;S
<=�2�<ּ��p��AD��;[��<F<C9�;h��$�<|����V ��;=P(=L��<��<U�j��=;�.	�%w<Gf4�Ƕ,=8��k�͘C=�]=��^<�	c<ob�<h�=�!���C�����<��
�1,����-����<@�![=��Y�ۺ1L =D@��6g=�n�;�d6<<�=!cm=1X�����=)M�<FI�B��<��:<�~}=�/=�μ�����*=�f'=�Oػ�z`<�>�<�	��A�f��,s�<�6�<���<gR<��t=�v�iGa<Z	��i���ź�����O~#������-�����Y�^�#rq<�.ݼȎC�eѿ����<��׼���;v�,�#=L�<Ɩ�<�Ƽ@���	|��?=�5<*���D�1;i�=&��;	�X<�߼Kp�<�=@p=�?,���f=�{=��[=��=�pi<��F=������sP�;�f���f�;��=Q���n =��<wU<<<�<k�I���=w�(=7z��
��2=�XS=�����ꇻ���<%��H�;lS%=�V���D���d����k�<= o��|�;4K��q=�ȇ�2-G=�żd�+=C�<�/�<�ç���<�����?=���H}�F'R=��2�!J��"P��a���*��]�R��bS=/�=<��<v[��1<��Q=������6=��w��xּ�n4��Y�;��<�N������VA.=Z���0&�T�S=�8�<�0�;�o�pn�����?A=;﷼����l��fP�;�D%;��̻�=5��=��?��&����R< N�;�<�.=��j��/�;bb���R�Yqp���M�;ă���<h/=�ֹ a/��rp��Z���ἂ����jh=�="I8=W=�y;�#��(e=.��<k�;��pZ�;8�m�R�V=�^T�C|�<��=���37=�0[=����5ܕ�1����#�Æ�寽�$�(=�NE=V=��<9�d=4�S��2�<��<�dJ�]I�</=`x=\HR=��1�i�	=��o�mD�<ixD<�w��K=�_@=�kI�P_d��TC��I�<TOs=�?>=�ɡ�XET=F!<�7���>����VI���<�
=n|�z&w<q��<nXD=u�<65F��*�|� ;z�=T0���W?�_��iGa�,=��m�<���&2��ݮ<�rϼ������;D%=� ��TW=f� <�4��.^��Ғp��a<�Y���
�<b�5=�Z���F!�7f=�&Ἂ/ ��-=7҇��MM=�F߼�L=�Wk=��<c:5�9�&��;�0; r�<%�T<�	�<�ʼ?䆻񳨼qM��q�<�1��͑��H=�:�<�\���<z���[�]��=b���S�=b���f���ɼv���$0=њs��ü/:�;�:ռ��<{���Xa=LUƼ��<�!E��I=
�==�(���^��pq=C�*=�J=��[�4�1� 2�:�7���rv��9��|�T=��<����&=p�?��mf��<ĘD<T�W�T�R�=T-̼�nq=��;��=V p���n=�+�:+&e<�P���j<,�<0����|=���<��<a��Ծ＀~�B�	=�H�<���uRлL̖<Rn=x�s=;�<�l	<V�;X�=��	=Ac���ؼ	��<.��< \�V�z=�-��V\.��=��=����m0=���=��6�)�P=;��<Cl�ӹ�<�;���#̼tb�Z�F�u;�bA�w]��X6�I��=�\���=P9�3��Μ���<�p�<Zm<�<�����=�܌���;�5�üx�ѻ���<ʥ\=�vB=�7��ɼ]��t���?A��}<�P��d5<��1=���)��;&���xc�;!$P<_F�<b =ɸ�<�I��h�W���f<��`<P=m<q,'�O}�����;Ez<Z��B<�T�<�A;��;Z��9#�<�(߼y;>�k�t<�/��2鼋̷<ȉ<e�<�<���8=�}&=k5�AA��0��w"=�� ��Qf��=LB=ߵ��.��büö��Q~v=!GĻ�4����>pʼ��J=P"8�,��<�w�<����^=�E9�7�c����b=>ü��4=��=cju=K{=��/=��X�益����T$W=C���=���F=�!���<�$X5;�A��
�<�L�<��P=�ł�{$T=�F<�g<���<
�׎ݼctz����<˅��@�0�T�k/��ʵ<�ݼ<�(��s8=�ص7(j�OB����o�
��6�$��:���<?�+=R�=5������<�@]<��C��;=� 9=qzE=x�o=�{�;y࠼5�=�uo=:3K=�ܪ���H��F=�?A=��ἚT���k��g��!a� �B=�r�@|U=��ƻ�S���&<�ޙ<7|<�3�<��N��i߼QD�J��/�>�` ��lD=���<��d���Ի��J�[qd���ϻÚ,�|e,��D��_��F�p��Q�<o�����g=���;1!��6�<�)�5�g=c����]�I�hO=�r�<���;��R�S�	<��K<�rX=�#ֻ@�4=�z=��"=�]<,A��ȗ<��� �<{�R<��;���;)�<9;K��cp�Wl�<Nz<Nĳ<|��<�?=e���x<)%=wCһ�<��g�I=.�a�D�<	�N=�r���#=/3U=�Z.=9�ּ�ه<���)��ƍ�<@y��p�wk�<y��<l���A^�����<�{#<)�=s�<s���#=�U���<��<�|��H�_�8�:=��O=4��;t>�b:�<�=;�;k�r=E(=F�ۼ;=��n<�C��m<\M��3�\=o�8�����m�H���Q��Ľ<��C���F��V&�iE�~�	=};N2�F�:p�(��N��wz(=Eu�<xit=�`���qn�y�8�Ȱ �Jj/=�����; �<�"A�V=	=��*�b<��PH)=���<�\�;<����}=�M�=����O�<�~i=̺���(��0:�,�s��==�<6P=�g&������<�z��J�;^�A��.N��*_�p =�<B�=Mû�$,��� �ɈO�{=��_=?���#Q���i�V/D=>%;�6���;�T�=��;9l⼖
=�1^=��_:-YB=�7����Ի;cY=��&<M)����� B=���GY�,K*��N=ϭ�<�N=�@Q�E	�<}p=ee=�B�۹��3��3�����<�B=u���l��
f�ͫ.��[<`���I߻1�;ю�<�޻%<,7�;������;�M ��+\;�q��� =��޼�l=U�)�b7���9T�=�"�<7(;=2� =���5�<��=���&�<�.�D�`�0��W����c=-�D��=@�ǼV=	���}<GCҼ�t��ǩ����ܻ&,G=�㵼b� ����>S�<��Ⓜ<LP=��2�Ee��[�=�f�;*�u�=�x�<t�=bKm=��ؼ���;p��;ـ�=�T=}�L�$����Q<�[b���e�wû1��<I"S:ۻ��}OZ=��ڼ=�4�=q|��	���<��g=��<�����7��;[�t=�Y=�/g=�p-�\4I�m����$�9X�<޾h��/M�[q�<�.��Gx�$�= �O��g!�Ĩ*�]+ڼ�A\�`�"�V����滻�L��S�}6X���|;��M�|��;��<�yͼ�~�T~k= H/�?x=݅4�F��<�����;Sx;��<���9���<����3h�ד	=��M�������s�W��Q=w8!; W�<�K�=�eY�(�c=�C�<�W�!=�<��źۙ;��<E�&;�~���<�%�c��ͩL��Ǽw9����<Eû<N=!"s����<���<�
ܼ��g�#U��=���<{�2=����=p�x<F�!=46{=�������N���=x�]���R=K4�;C��<�+�<~���8Y=YFT����;(\=d>�@��;���;	�<�s����;c�}=/��<+S�<�W=�3G�����*=�S"=�4X�[_:\�΍�;�N=�� ��<��bԼ�bȼ�����߼"�<4 J�$�`<4po<����λÁ�<����\� �W�3�k=^Ʒ��v�<�ܥ<z��;A��<�C=�,R���+��c}���</��N=:�`��@=�n0�cļ��E���d=��<n�	��r?�Z�N�5��<m��iû<�G;��&����I�_�&8$<���������,=���<M�5=�h= d�<U�O<��>�n�&P�<�Ъ=�����<�^<�@�<0�.;v=�0�+=<�<�PH<��;d��:�X��,;�<.�!�������<Z*�<��d<`��<�<I��5���ɝ=���<f\=�� =��'�i==�����;=w�̼�L:��a��8�;�F�<�^u��T�T�L=��J��5�<�G=H;=*�P9�X.<�`=
�3��=����xY�س�����U?��@<��������M��Ђ��T�:�f�;^i=�l=���;C��iym<��
�8�üֻ�;mG�;x���==6�2��� =Cȉ�02E=e=.�7=���SW=�e�4�,�6=�1<�n_<m5�<Q<=��z�j<N'ɼ���d<f�1<g��<=мga�9T��`1��+.=��g=t �Mj<	MW;sU�;#�ټ�� <��<��Z��"���[�<��*=[H[��z"����s�"=��Ǽ�RP��B=x�w�lm<ǥ?�m���j<7mX=�8�7�9� 	�ma<������<q=��&�~<}�G��E<��R�F=�X�;ص�;/R7=��=���=O�\�sإ�c�-����<� ��hZ";]�Z=��<�a����u<��=�B�0�L�M�<�1�{�@<��k��<�!:�0I=$Q����w��<ĸD��I�<� r�;a��.YO�5�����r�!��r����=�J�;lK<u�;�e=��Ļ9��<|k�<p=��==��=��'='�C���=';��&�<{&v��|;U'���d;=���:՘���N4��[�����aU�ei��쌲;8`�<p^l=N���n<�m5�)��<�W�3)�<�f2�N��<T�<\b9=�k�eB�<8=�Q�R>=�6�[�+���<9j���+�f�7=�u=�e�P�8=�f�;B�<�� �U��|��;�N<0�=�3=�B�<q-i<�r�y>��_�3�����<� =�8����۹(�< .B;��g<��>�939��H�*�#= `�<�S����#�/7���P��Et�,q=�O=X�5���;���<3u[=�;��eݼ85�:���+<�y�}�o���,#��#?=oK�&*!=��#=��=���W=ua��{=�4 ��s��'bH���<{<�d=)���_�<`x1�!�R=��;5����ׁ=؜=5>\<-T=L�!���O=޷*�H9�l�< ���=x��;�;=�7<��W=�<6,���A�OsH=�>B���y=�ژ<`�.�I��;�d���C�*0g����+=@Eg�]-�<X !���ؼ�K�<Ƌ�;F�]����L�q��<�G%=e���~�Z���4��C0���K��4L�vNr��lw=��B;xU��+�O�/%<	�	��;��d���I=�� ����7>=^;�;�՚��=r�<B&z<��^Z\<��h=	}�<'�U���D<U֚<���;�&��N�<7�R�0�：��z+E��w�<�#=��<���<ϔ<���[-=�|*�o#�<]�<0���u=�˼z<L�]n���<����E�;��缃YN���<<2]=/�=t��<2��iO�4�f;'-��X2�,�7��=X@1<v�<���<�H�<�=� +<x�����7��ؼD+=�S=L=�v��������<�N��#�\�<�.;��kP��}��:�c�6��i����</��<ޢ��f++��nF=��ջth8��.3��,~�a�=���[�m;��7=�)7��E�C��.�=TM@�υ?��?�<r�L<�J=�j�=K��m�O=y���o=�9%=��<Őc=o�=D�ڼ}+O�D6�*?�<R��(^��V�	t<G�7=�#1=�|3=��=&VL��4:�H=�^����x�Jx�<��<�O���E=o4�yC�<�_�;s�<�]�j�<=n�*���<�i���(�;}����\�<B@л?�<�|ɻ�ۼ�YL���K��ģ;��<�L�~i�;�����I�<��<a��f#��h�:ޛ<��2=�Y����<��M��4X�v�k<dc^��O=�ٌ�P-������<c�'��fμ���<�c<��(`<{�#��<��=�W�f�<�O� B= ��!<&�`=k!�:�Y#=H5�Bn�P�W�j�<T S�R�G�JB=�[��u��<��J�����=��!�Lf�<=��:y\<�		�_���L<C�ѻ?9Q�J�3��aѺ�'��&X��Ӟ�$�꼘B|=��<��;>�޻����NJ=O�-�A���pͼ��ּ^�=i�(=�k&��J!��<�w�<��=�P=uE�p7o�3�����}G�kDK��2=�.��eM��P��z��<�L�<]5=�o2�_1=1��:�&�Xy�<bc�DP�c*��ӹ��?�<�X~;7(=X�S=5���I��<�<h.�:���;(�P��˻�շ��� =ۋ��-0���3=:{�/�=�A ���`=%G޼]=I=�˲�V%{����R�#����<��<}]z=>����<���;n>�=����5;�!����d=G�=k-k=%���f=�D<�%;���]�)�==9��� <2�E��<�⼙^=HG�<鳌<c|=�}�(��<l��WҸ<fId�:*/������#=9�6=��}=8��<9���Uj�L<>�!;��L���(ݼ�~�;1�,=$��ˋ	�ƥG=b!M=+�v�u�,=z9<��<�++���5��(m��g�����W�<��?=E{\����<7tԼm=�Q�;$]�<�������9��;M&���Ƽ�� �=d<Cnk<!���S='�P��=��=�$=��T��C9��% =�l=�J<�����^����Q�8 =iئ�Lٻ<]��<��<��=�B�CJ=���ż��=N|N<Q:_='vB<c1=�����˨;�x[�-�8=E�=��]�.ؘ<��<(O���w~�r�=*F=&I�;U
��򍽃0�<��<�;=m֯�_~�<@[w<�0=FM;�LJ��j�o��<�5���l\=���</�ּ�Kѻ���<�[��H����� ��;�<.����K�������<�s=.eJ��g<$7�ۇ*=�Ś�Ha��lt<�{C=d��*�RFջ����،��cR=T�.��+0�/=�/;��[�:F=��k=�k2�3�q;�x>=gt�<�v"��8A=~�+�2��R}����9�����_pa��u=E�<�9W=3��<������:qͼ�K���W�R#<���<�0������1���ܢ����<�U<�<�'%�L_���J�=�Co�MOu=v���G�:�_=�V��v\��zN=�BX=o��<��p��>	<P=ڹf;G�G�?�=��<�������0�`�a����<>=H�[�@�X=yw=;��c�G��0==d)=�I��L��^t=��1�	�k=R�<=��C=%�ټ�R'�a������<p=Oj=jC=��ռ����qF<���<S�ɼ]��<�Fc<�=@�/=�۝��=�1������'J=H�R�a�ѼJ눺M�=H�4=S�>�n�<@>���4�kt��Uڔ<I-˼#$=�}Ƽ��'=ߙ������6B<[�P<�=�7����Żi���aϼ�Ѽ��Z�)�;=6=�0��>:�F�P=z� �m�㼙��:��R���E<@����l=�
=B�1��<y�u<�x �v�ʼ2�Y=e�;���=j�ɼ��4=��<�ӎ<�Լ��V���.��R2�k^����=��;��	���;~i<�|�;D�;#�gs켝g��)O<��9��,_<�(�������)�<p=P �:>V=�sV=5؆<�x����)<�r<d�n=���;t��;����?=Rp��;L6=���<�p�ځ7��&���4��Od=ZE5��֠;b�8��J�<˻?� �}�C��<5k�|�b��ߟ�v�*<(t;x��<�qB=�j��+��;�~�<{�k����|{�t�
=D��E�ڟ���π<��H�T,��8r���p�;W�;2�J���/���;�zr��d=쩀=o�Y�<h�;Y���2 :����SI=����l�<��3��Ｑ�==/9S�i<d�<u�8=V9�;K�9=�f���%=�tn��(=W��:�I=�8y=�E̼P=�A)=�9��6=��/�`9漗+=��<���BI=�jú�/.�\�	�}�F=t���b/���K��4==E��8���>A�<��3=v���	iA=�!=�F�<ǿA=�3l�A�s�B2+��*=�Ю<fFn��ZF���e=e�=�\=]�)��x*=	=��6=��;Ox9�582�i�Y=5g����H�}� 9^�@<���1�.�.ռ�S9:�M,<p���R�x���o�ڼ�|H�-�����6=F�>�[�V7��`��Cf���I=���.=p�8;�.=#΀����#j��- =��<�%,=K�2Ka���<��Ǽh�����<��7=q,Z< T�<�|R=�H�<�i,<��1�4v�:��V���<R�=�4��@����;p+=kVO�-�Z�;l=z?=�9ۼ�E$��9=r]C=�T�|��([=��ɼ��=B���#��q�L=�����	���Ѭ<s躳�c;ez)��z5��d¼ �_=`�4=�A=; J=�p�@�h��J;��i����;?{�<-]�<�M�<1&=��;��I�<2�?=�٤��ݼ|녽��ͼ͟4����<���<�.$�,�l���3���<�=��ȼ؝'�������M�����n�C<lڼ��1=�")��$���*=�R�<��<*�<L�=`P+��?�< V� F� j�\7��n��<}��1��<|#%���J=��<��7���M�@)B<`l����&<�R�i^�<�U=9@��<2�<"�6=�g1�z�<�=��`=d����0=��m���[�zp =��a=ώ��~=B�B�R�[�ƑR<����Cq=Bü�a����I���,=�A��U�";�;c��<��0=�'������=ih�<�w�Y"C=p�ܼ��E/��Uj<�lU=:�ἌB����3=���<���>=S<G�ʍ��W<�����=^t$<4M.��$�<B�W:��`�v�;μ�0���<yF.=Ph1�6�<)X�;��<o�U�Y�{�_�;=�&B�B��<��<Cc��Č�+��; �+�Z�I=Y�<��P���:X�$��H"��v<��T=0��<�Q=J��;I��f�O��r;*�6���MXI<|�Z=����] ;�z=z1�<6$+�]1 =2C��ޒռ�D<��o@<=�9��G=p�<4ރ��<=�d`�\��Ia�<�-!�y,�<�����D*�Nk!=^}b��sŻ"�o��ˉ;=����\�<(�1=S�c����D�=�ӥ��M=�ҫ<��;��*<ȡ�<�R7��1(�"�i���<I�K=�V�����<y��<��<ߔu=�Ɛ��);��]�k0Y��$>��ւ=����U�u<�@@���=S"����:>��x=��J�����,H���;!�$<H���u�<��;xxD�qoY<��>=T�;=�+=�==@c<�.�=0�&�V�6=9�'�F`����<��/�_�����=~'=�=��k[�=;?��3�?W�n=�?W=]$:=m<�[I=~ȁ<e:�<����<	<O�`�&)=��^=�<~ Z<1��;�%���!=*u=�Bh<"���f(�+>S��������G����;�R�;s2;<���(W_��������k<��m��:���A<�	�;1��fI=��k<�u�.�6<������~�Ӽ_�<��<�C��a�,�ל��X �;�9���'��W=�s==ԞX��<�;2+=I_�h�,<��'��")=�_p=m������L�=�i������.껊��<�P�<�H0:��;�j�<b�=(�@�d'`;37@��jF<W=��߼���)q:݂�Q�ڴ7=L�9=S@��g�<��t=Ac0=��v�L[O=:�=�j�;�=�<gZ=�ס<al�������7=z�M=v==�A��e�;F�����=AM������"(��O�`t7��v=� =��<��9�����p�;;�#�<T"�	�R�Ƽ��
����6^�<�Ӻ[:��JW���]��<�<�/���=ɷ�o�49#���<`=m���%<�C�R�'������T=��Z��U&;d�%�� 0=n��h?�ZD���<��^�#�M=����3g��(E��C�<��7�8ą��J꼁ܼ��@��2�<�VR=t����E<�����*ü4����
=2���}$=���<]м��="o=��;�>��R��ϻ}f==����%�l}��9"����<�.z<�TC=���h[�<�d�8�=,k=T%�<=-g�6���70=�U��2伤T�>N�<���<�T=��y<�	�F��͵ӹ�]���}���<�R)�[]}={�����b�rM���N�/�d;�(c�2iy�?�O<��v=�)�H�g��Ԉ<>�<A���%�<���<�3=y� ���ż88���=��<�v&�5�6<��<<�ֺ~Y�jD��t�Q�����7a�)ߛ���;X�μ��I�(q� �ּc������tR�
��<6K=0�<��ڼ)�(=�--<�d�<y�==�(�;ͺ	�k=7ӻ6l�����1��5���NX=���d���V��+oh��g���g��;[F����|�Q��o=|r:���Y�i�����;�hF�7E��l�K�=�N
��T��������<b�R=?�=������K~���Q=�=��c]<��Y��$�r�H�i���L=�z����?��=��"�B~C�/+�v�6<KӰ�m�-=V�������{.=�z=��<�)�<���;$<�q=H�ԼT�H���:y)�<u}3�}��tܴ��Ҽ��<�T;�w�"�(6O=�Y��ۀ�y��N���n�j=ۅl:�A=���:��=��$=i �:��n�]��0|�<�`�AW�<C����U;Kk;����=��;=`��m=b��X���T��<�X#<n_�?�p=c��<��!=Oq�ɢ�`�u<Q=<c4��߯F=RL;o�ͼK�=P�q<6�9�;�s;H�&�a�D�r�X=[�����Ӽ��������炽]�2={��u��=���<n�=�j���,=,Y�<62���.<�T5=R忻��b��U9����I��<��<}���:�e��>L��叼���M���<�։�a��#/�Y�s=Lkټb���#ZU=����q� �׼���Y�5=�_m�9,�)�[�*���<�x���Y�<OһV�t?ȼ�=�T�����^y���	=�C)=�����~{�3�M�ǣ =J���{5��4=��L;*�@��0=7=�v���<�މ�6�#��|:���#<��޼EX`���r���#I�<Q��_���9��|�e<g�<m�;	���e*T�uF=�%a���1=�ە=�F <g`���W����<ը�<N���n��"��9l=3g��<D����0=��=Rb�<kG��u_#��ؠ��+8<�9�<?M����X<��;,�:�h,a=J�n�����6n�����YY�1!0��GM; �	=��<>Ca�:-��);d�=����#/=�b��� ��)Ow�S��.N<��`�~v�n�*=�r)�J	�P�C~��\e�=D!F=
U�8�=1�ߌ�I�^��\� �9�BX�;B{��PU=���;�8=wJ?�ף=�ɑ�,�n<kMy�,��<��PH�;�gc=�z=B%v�ླྀ<ѩ0�[��<  .�q�s�:���9���;H=Bȼ���=��?�(���c�TPB<�?ļ��<Yo
;$�=�v��mȼ�/˼�?���<�=�w:�1}=��,=3Z0=�=�B��N�p�V=���:e�)=���fr������)����:g4\��m��-8=O�x<g��<���<Lwy��q�;UЋ9��=��a<&w<`���]��<ꂞ<HQ=�ݼC#=<�=nc%���b�-��<��mx"<bc�����2C��$���ļ��<�BE=H8=��<��(�ڻ!�4���<�a<|�<q?ļ4b=#�Tn=��+=�-=�7�<�ۼP��<�p�;y�<�g=��Z=n0��{�O�2�����ٛ�� �dѯ���p�8G=)�e�����t=���=	�<>{�<�Ɓ=���H(=�&���:�,�U�$�H���ݼ+#=��E�9=@�2�|��F����:�蚼*��]S&<��i<gX��(c=:$�<�ӏ�a�8��0=Х�<��d<D��PU�<Q�<��?<�ʁ���]�٪��jļ�ǡ��g�;�
j=	;�Z���P���D�j�<�	=
��B�P����k�@�t)�t�g��ļ��8�ͧF�}_I=�1J��')=���F��!�����p���\4==�dz�n��#��oc�<u�<��H���B��`8=����䔂=Sn�.b=u좼�uB=�$=���[��W�;^�=��;��<1�Q�s=�`=q
�F��=�һ�j�<��N;���<�-�9.� ��~��\=l�	=�w�<�Q��^�<@�<�����8=��'M�<l1���+�W+=�i��O4�6H��L�<���<�(~=3����C��ڕ;�~���sL�ȇ=Ή����(���$=��V=�iS��0�M�=Y߄���Y�Ǚ���`P��BG=�U��H�&�P��o%��y�=�*��Nǻ���)�2�w=���J=�^�Ms5=�K,��e��N�w�<Z ̼#���|.�<��w�S�|���<�v�:AŮ���"=g��<�g&=tq=�����m��A<�˼��*�Q��
�<�#d�����e �c���
V;HB'��B�<M�'�z9?��c=��B�ệr����<F4*�_:Q�
�*�Y�O�?�=��)�Ѭ=���9��6=g=�+<�I�(.J=�^��rF=5�;叩�%�=�Um=�e\=<=֘<=F������;4,=����S�3���S==�<k��<�I��=�Nk�^D��L��[�<�8<��w�˕!�|�v�	��r�;��=:�����U��:�@��/�Tj�0�-�Y�d�f�<���<|TY��;�	/;���G����<>�.��_�<Z=�]�<z� =&�]��+�X$�K�k��;�V=�4�<n��'s%��B���<��&��~���û����nN��μX��;��+�� �<�h�9	�:�W:]=�R��a3�Q�9���;<��<Sy=~Ť���(��̡�T�!�oU;�{+��^<!G��l��<���ܼ��L=�z=�����Q�O,7=��o=��t=�8���2�C�$��!�=�G���T�[ak=�/���?�;ׁ�<A�c�[�:��7<<܍P<tE�C=�����<�=�e=*wh<�H�W��m� <�9����ɼ��ƻ4(�<S�M�x�^��Uk<�#!��5,=!5��d�c=�?4�z�(�� ׼[�e=K��U7=�>�6��n��}9M<���<%�=��2<�|%=d���>�=�I=��)����6��ǿ����\��g����_�F�c�=?]#<�t#���;M�=����������H�z=�<�C��<)u��J�޹L����=:��;�o���qV=���
�\�B4O=QlU:)	���X=����S�*������J_<k�h�� m<j�=��=�^�<u=����ڛR�XVd<�IC<�~��]=�wt=�8=�7�<� �<�&=�= ��zW������S����kʼ���%�Ώ�J�0=#X.��=>=rϩ����5��=f�=��{��� 6���LQ=p��<+�Q��5���U=Jo5���(��_`<:�h=��N��H7<�/M<#<��@��~��o����=�A���3�h�\�[�=�3[�:T9��t�G�ڻiȻ��H=����@J��ѥ<�c�h�O��ۙ<��;H���G���<�9�;0�=��t�$�Y�<��߼'I�8G=I	5��3=��X=	i=�M����c��<@��h{�;�X�t�F���<�=�&�<Ѕ
=S�==����}�)=���<+��<0�E�(w-=���O�P��jy<��d=&�P=T��2N�Ғ���:�'C=�f;<{j<=�H=���<��}<5�}��f~��>=�<�U�=@�<\������<0�f<!��:$b<W��<�v�=ϩ�w�=�"#��L!�ʹ�<�%=�i;��C=jd�8��g�<��ʼ��S����<b3�;r?=��=��Y�A��<�t>=�-=����j=��d=�e,�IŻ��*�Ķ`<DB�E8=6	���H=�� =����#����� <� �IN=��O=����@|���(��M��<=m�<NA���?=M����r@�MM(���*<*`<ۏ:��k�k=��;;� ��B ���G�Cy���r�������5�d<�j<!v�;�V�v�Ѽ"4ļv	3<���u}��s����<!�*; �h=B[)=���N�:<�n8=�m=V����x�Wf�:!2���0=կ<�G�i�=�J�<����:$=Q�$����<�g�V�=�y�<:q;^l=�X�<ɬ����;�#q<�7��E�q����<�3C�P큽7�<��~=	��>�u� <$�d���<�c:��=���mD��)?=�"�wSS=�~�<�6���dG�#����T&<2d���3��bL=v�X>=��׼il,���:��=�һV=w�=m�l;QZ�<5�мq�<ss��x=��<Yg�<k�L��T�;�'����<:t�JU�֐�<]�;(q��+=���<N`Ǽ�K=�NB�[������;����<�0=�ZH��=X����<�9=A c<��
=�v+�x�#�jp+����<Ñ�;%|=i�<2y�����:��Q_����<`�L�%�@��!��c'j� ��D�=)����'���;�/�<,�u=tƯ:� ��=BB=!��� =,��<�逽O�<&�G�/��1$���?�l*;�#=#>��%w=�q&=^�8=:=J�)�g}Y���=�yA=�70=Le!=_.�)߳�<�
��\���e�I%3;.5�<�����1��<��g=��<`�S���C�5d����;���:1��;+���ȵ�@wU�/W;�^a��&R=Z�\�,��kz⼪��=y!(�hq:���<M:U��	�%�W��!�����x<0�<�Y=4�+=���W��=���:��=N�$����6�}=G�
��L�</_J=�� ��p9=�3����;'�"=�������=�:	�9�����ʫ!=V�<�4
=?|�<��o=(@<�n�;�W�:5y�����<�h���c:c5=7Xy��3���;E d�Q����[�nX"��6���=.<!�%=f�=���R�S�=D �Av<�X![<�J0��_E�� ��kF=�ܼ�P�<ʤ�<r�=����Q=5l�8�T�NS=4{=و.=�ܴ�t����H<���-�Ǽ#<��=ǉH�Q9�;:��W�<!����@=�O==��@4;,��+q= ��8՝��_=�K�<K2j=�+�;���{��<�)[=|?�<ˏk=�/�<5��<��g���u<3�U��1�<��x��~��(%<ȣO����Q�$=ER\=��=�_��y�m�}<�΂=�&V�-TO��j�(y=��;�N�v���3�׺�h��<V��5�<0�s��#=/����g=��t�Y<�-=fh�<��<�@<�D`��H=v�k<����)�DK��<<,�<�\=����6����8���<�V|���<��b< ��<*�<O�-=��켵 �;@�<l꯼]�=�5�<���;/� =}�O�+�?=�d�<�V�<񚹼�ZQ�[�7=N^ż��`��pϻ+(<ߦ�=���<�X�!��<�<�񂽏��;w�N�5��qG��VN����= A�<D�+<�^+���_;�,�8{=T=a
ȼc U��SX�?�=ԇμs>=?�4�,и� �i�cBO��@*=�O)�%e;OGq�' =�@,��id�R�����;�*���?�e=�j=����:0=I7���8��ӕ�l�����<o8��@󟻂��&ȡ;O�	=7P����Ue�=�1=of;��:s
a<II�Sv9=G|�;�<%�<�"=�;G=�:��SG�A�e��=�]/=��}��NS�z���-�uLG�/8[=`����<~a=&�Һ7oF��-
�#,���A����:º=퀾�gs_<N�5��a};y��;��:X֢��eݼ$
�<��1�/q=~^�����;Y;,5.���D��oo�/v�{�u;I{�|�w<�K=&m������
�heP��c[=����}<�E�0�X���b���;�ؼ������=00�U�;=TBx�.Ϙ��i�4�Ѽ���<j�.=���1<�:0=�m���`c��(�:��"���к���E\��=7L#���=F�)=gC:=�糼eB=�^;�C���ͼ=-�<����<�k���켉�0=n��:�<<�6�O�X��7���$s��V<�_E���Y�5�3�lq�<��P�`A.�Gd�;�����1)��aj=�=g�Z:5��fC�A�˼6�`=�gp�%L�<�Q�����r��h������;73=��<��H�3�)=� U<���$Vo���;U�=�/=0��;�1�w�#=�i�;�lS<_�6��6O�Bw<�]w=Y�=V��;�7�z ;�י=�CƼ�Q>=A/,� I�<��˼uS<i���mh�����b�������u��rK=~r;r=�U��5$=R>�\�;���Mn�<cZ���ռ��M���՘z��M=Z�4=X����<ng��'�f<�`5�0=A<�GU�oD=��=;�=6RU��b=F�l��H�<bo�2�=`�ּ�r� `<o�J=��=�8>����M</�U=B�*��ޤ<�C����<��༟K�<����wX6�pM缾�ػ�45�3y=+V⼌�6�/��R��<�C�< �Q=�������<��3����<����C����H=tvƼ�D����<�<�9;w`h=��;�&�����<��j˔�,�=�k�"�7�~Ki=�^=S�<��`��G�<&�	<�;=(@<�7��+�^�\���w<�vؼ�E==2ἤ�<�4?���e��{-������E��kJ�st=�3=}p���<mx=�Q[=���<�tw��a.=�='/<T~�	���,E=�*�hb�<�=Н0�U�A��KX<"�&==RL=��.��1��8�9=[4	��1�|s��I��::���G��?iH=��.��
"=RZB�k�=�:���:�`"/�F�(=X%�<8>P��`3�=a���
=������C=B�4=B\!=N}�<a�<�>��,��a=�V�QN��f޼?�-=M��~��ȼ�G�<@y=���%��u; ���I=����v�-�ߦ����*=\<���h�<��L��)i�)B=�ύ;w�;0��;=/�2��<I'�/H=��S�i�@�g�~:L�<�j<�O<�X�<X!=�2=ɤ<��=�}�#=��T���\�|=�=��d=��O;�H_���ػQ�;A
���:��
��,�;�l��3<�$�F�|=��%;cO��)�����G=��<�)�<�B=�B��]=�n�<�!��b�X���yf��G�;� ��Am�O�<H2���W0=u��paC�('�<[�9��=�d��d_q=!�^=f9ݼ{==����|�</	2��)��t=��]*9b�<���<�}
<�h=��=�^�����kD�<i�)�"���?<�Ԫ<7m+���H=�m=��g<;�e�Y���1<�/<O��O4��H�=K�<F�к�"����m=y�<\ˣ<�7=L�=�E���?Ｎ�X<C=���<C�5=�p<���@"�<���uC=Ln]�u�!�6�< |�<c���wW=Ѿ�<�9L���>=�����nE=6��'�q�}~5�(�=v� �D>�=;�Y����<\sP=6���q���O=��W=ew���4��&=��.=8Ƽ]�0�����p<=��<Ӯk=ڃv=���{�=���<��= �@:��o�رF=
%�<�]=+�k�Ü�МѻY�;��-�560�8���53=G� ��Q�+q����;��ֻ�?=������<��=���<�w⼹:=z��k��<�.=ȓ��2W<�r���2"=W=W�f�:��i��g�g컼D�k�����⧺0vN�����]=�p�=�y��ْ�G���TA��'s<��Rj2�D�^=i�=�bu=����Nջ�����E+=
�Y=T��<}�?=�h��B�<1V�����Լy�<Ӷ=�;��9��~/;��=!�����(=��=>n�<в輤b���� =7�-�����vf��$k���<�ވ;\\M�AaG=j_?�U�t�S\�Zm=I|g��������~c=�գ���6=�ʻ�0=�u�<��%�<�D���]�*ͤ���ן�<�E�<���>=�KmI=�B=N�<	�<��C�$������r�pi�<xvn;j=�uC=9����]P��IԼ</)���;��3=������7=!=�-�=��C=�jn���R<'���v�<E�<�yw=54X��剼s�@:.��y�}���m<�y:�J��iM�O�K��T�<��8��*�=�r����
;Z�@��<���d�<��һD�i<zd<W芼D��:�X��N�D=Ox�;bzU=�1�ɛ�!=��^1�F���h�l6���c=��q=}l�<��p�`q�G��}���wf�k�H�B����e�\)=K��<rh=oN=��3S�<�Ӽ
.2=`� ;ճϼ���W�Ѽ.�<����"S��Qi�@�=�i=Rxz<\2t=�V�<n��<�����vy�d�Z=�h=��
����;�'h;38;xD-;�$<��2⼒���ʐT��Ʋ<:�"��#&�s!��G����@=�,󼊧<M9���0��y<F����o�@�8�M=�w^�d���C����<	���y�;!��<�;�<o޼�(-=W�<�z�^/��-Y�F��<?�< ���N��x�<�%ؼSkA<�#U�e^3=f�^=������+=�&;;���M<'���W;B�viF�?���d�����8<�,��w�;H��,=w�ȼo/(���J=VO�=����1㼗�%�P�+=ߨ�<lɭ��H�;�+=��;�3!�d�X�B�-�H���ы���R=�:��92�6��m=��;P2�<#F <Q�
�9� =bf�Th��P�<A�u�zu��1=�;���������T��r���_]=yd�
䮼1�5<j;@<�9�=X�|<�M|<��t<�G�;.�!�D	=�S=BƜ�����J����0<�s;�-?<Nq���<+�6<���<�J�~�I(ݼ��</�<5��<rF�<=Vq�<-<[=�i=���֗<�?�<~k{�h��d<l=e��;�����0����<�o�<
/=�
�{I�\=߰0=�ϵ:�q>=��n=A��<��k�<):�y^O�O��{~<��Ǽ7�ƻ�� ����<q��<�=��@h�đa�(u�<�»���W8㼰Bj�9g���\/��e=�n�<���<G�Y=�0�;�$<��ͺ��¼��<w��<I�=T�J�-<�<��<�R�2r'���=К=�q0��,�=��v=�h+��������Z߻$�#���!�=�5�_qE�ng�{���=�6�<�z��ew����;��<��<���=�B�����V;e���<��=c<�?>=n�\�a�_���<+SI<n�\O���<�\����
c|� �=F�^�H@D=�n4=7�F=�9=�mG�?0.=Qш<"#��>4��,h=Ɲ�;�ZB�.���<��#=Ri�<�M�	xa��b���;H�:�^��:d2��<�C�<P�<$�<:��<�[�KWr�ٴ<;�=�bڼ��<�b�i���<�=/�ˌ��8C����<~�=����Y��<q�u�Ý<tGg�MjT=T��<�nA��U¼�`=:�R��M=�oK;И�<�Y�;������<���L5��M�<Ch@=5o���mB=BQ��i+)<��=�'/���=s=���<�e=�j�<���<�=��f=�gE��\������Cm��D>=��#�y�"=F���%�Yc�<p�ڻ�S�<�y'��X-<��B;KTx��`�٪��mT6=!+�GQ�q�m=4��:�9��M<��<2/<�4�yV���BO�	e<e���&�\��<�s2=�%��Tf�;�_ =��#�OD���=�\�'3*=�y���Y:g��<=�*�EN/<����U��<��
=�32����+%<I�$��t=��X=��7=��?��Q����V��ﴋ�s=���<{=�_,�t��<x�=
�=#o������?; <�T����M�t	�[�b=��=|���q�)=𢬼�=z��=���]�j<�7N������7G=v~x=�{D�[��<��<��k���&�b�7=[������熪�"(V=H�X;( ��s><B=�<�[9<�c@=)U5�Pn==i�q���{=��P��ۆ<*^�<�z <t+���Lq<XL��T3��t���|�
Ϸ���=��l�1��<��<55�<��Y��O_�!�<����H=��H=�:����S���{�;NR��ϰF�G<����Eϼ��w���;�x=.K�-q�@=�u��պ���yֻ:��<�>=�}=��N�"y�20!��K=�$=%����
�&v0����;��#=hGt��+:S^��KN=�9��3��`ּ��=����Z���a[=�U�<�φ:��-��C��S+=�R
=57�<���<yg�[���牞; �=n��;��E�R�<�$=������< �Q<x�ݺ�A=%�;���;�����6�[Va���S=�$3���<}vټ#L���<,�$�4=��i�	�@=�U=�#<X(<r_=�6=��:���}���; �{=6�)��h=$�</�K�
d8<s}�;��i=m4='γ;P��g������T,��%;�X�B=���<+Ca=򽁼_r�0"�����<�����i9=~�(�x�=�j~���m=���3=�����;Y�^��<f3��h=�=Gn\=�Z�vvq��E�W�<9�^�� �<T	~��hǼKz.=L�r<_+�<����=��@�; ����v<�0
����<�&�<���<��!=ac�����<�XN�m��<v^��1��:=׺[=kkB=�J�G<?���<��x�����P�d��4=�=6� ��^S�G���0��
R�����̼o�J�}L�<$�
��Z�<6Zʼ*tB���A=��\&Ի.߻������<���<��x�������G<i�;�]<�H/��q)��[����<KL��~\=�I���h�I[���<Kx���%�<����=t<i�X�M���C�į=����P�<�'J=�/x=ۋ=??�<`=�4hh�"f2=n{i����<�"y�V�B<���<>�D=d��G+!��YQ�k�D�^�=�Q@��=����<j@���5$=Y�����uu���<�Yļ/~{=@q���{4=<;�<�
���,�<�����.$=��N=�5���J�{<w*H��0� u<���<�s�<n�G=|<�h>��\���X���c�g�u��P@����<�	=cE���3=��\;7�<�O<�����Q����N�
�K֍=���<��=�Jr=�I�h��;�H=И�U<z�;�PH=KЧ���=�qR�yrd�G���=y*e���;7D��G==x<�Z�Jh�<;�ex��5=�p�<��<��<��{'^=�ۘ<�A���;�9�<ľd�����^�#�/��<6��\=<ZD�:�B=\���c���μ[�]=�1<��^=��t�����8��;���<N�R=&t��fSA�MԒ;x����;G��u�;c\<�<C�W�ü�g�~6=ሼ��[��Y�w����+��,q���;�b����=<�h=u��<��R=��=��;5�P=M�Q�kn(=\�#<y��<u⼯	�:�!=PA^�������ӼH�<�q��\�ı�<�9�<9�<��U�<p_���T2��;���Z��);b=�x�<�p=�)H��o*=�2���N�����?=�2�<U��< �=����E�Ŕ/=J �:ߙZ<[��68Ѽ��<��'=�¿�m����Z<!w=��C���E��m-=G(<��=���;��0���)=�	#�r�e=�9�<��=�eE=7J=wѺ�Z=p����������:��<�-J=��2�t/)=��<�J��S��F�.���>;�a=�7d���<BfJ��a���1=Չ=<À¼;}=��B���a=,�[=lNY=M�9=g�K=x�&;-��� <�<v��y,�u=\7�8��6=�������:�K<��B<)<��x=��O=	 =̪X�
[=��Z�!�(��.��l�����Y�<�}��f��<��V=�=�<J�b�%=s��?��z�-=�&�BB(=����^<5���o�<���<C��<���;�����-=��b�1��;�'�RK=RF��=�;����<��:�\�ʼ��'�Tg���$�</���.�<Gy&=������<yJ"�~�>�����x �T*�s��<�i ��Zo���<�JD�s�N�trY���.�$"{��=E �<Y)<.ݣ�	'=M�H�X�c���s<9��w�B=�������+(���m�th���H5=;��<q+���d=��K�!�_<9[R=~�;%��L@=��<9�=>���-M=O�b;�jG=$�[!���=<�yg��n�
�м�\���1<O6�<0Q=:0<���<��+�P��;{��d�&���<�S>=RP2�P���:=:��<���=6s=�m�<C6<�ۍ;�.����ټ?�`�I�mH;y��9�C==V?��@^�c�n;LB��F6<+�#��pu=��4��l�<�{X=3#\�J��r���?V<z\��l͹���W�^�U=�������-�=�j=3㾼��K<�h�<�џ��L�P=~�O<4�'=w�ռ�hV=�+���`f����=����M�<1��<���9Ԗr<#���]�<�v=�@��;8�<��㼦-=�y<9 !=�<l���f�R<kC���rU;�q��׎�%�<��}��1�<CZ==�j�<Ȯݼ�=(W����=X��<&q=��<�J�{�H=�
���/=�uA�<��<2="<ڼ ���< PN�"� =E!G��۩;7US<��
�9�a���� �$=|b=:=?b<Qu.�"l(=������);�廣�'=< �I��<Y+�A��^QH�WPb=ٌ<o�L=��6�`���Vl<�n��Z�2=��<�	��Aͼ�H��1=�e<����=�:�Al=�l�N =��9�tp<.<��οe;��<wü�y��|8�a�K=n��:�;sg���7;�S`=�G���4S��H���g���5=3C�(Ƶ��ş�\A<��7=�����<.��%F=���:���<u�Y�0����99=Wa=�?V=�AM=����.<&�_���0=<2=2=d�C=�X=�5�&���?�1=�_='0����<��J��x��b��'a˸�='P��P=�%6�#I�lI,=^�L��D,=c�:D�<�����_��V��m =�\�vv���M�#���GjZ=xv�;'&M�{Y�ř<��R=� ��t;�N;P�)�~.�<A�<0��<WY�:=�9;8J<Ї�:��;���1=�5&�w�?=*���
�ּ���<-�s=���k�>9&<PT���9�|5=_ =��;<2v�=i#=�'�<��3=2a	��0�μ=ci��=x�~<�;ϼ�̼z����n����W�;�W<6�缦Qa��D�<�^=�Eۻ��u���3=о�j��Ǒ�=>/�<�Hܼ@�J�?m�&�)Bd=*dp<=����C<`����.�<��3<��.��Q��X W<C=`w=��J=�݋���B���&�Z�=GDT�8R^=��k�b��Ⰼ<!�����y�:�ȣ<F�;W�;Q��A΅;��=��<�\�<�\<�ʅ�q�(=*>=�ټJf=͗6�$l���x<�����z
��B��E�<(�<V, = �p��CǼY��q��<d �<�5�?G=��4=����pRF<�>��]70=
�S����#=�=<��<zi�=_ּ�'���ZӺ*}�=}�"��8���*;� ��H=,�����;��U�{	�=]���Ǻ*���:=��T=�������]�=�<�Du=.��<��;���<(ۦ�G�<��Lú�&\��:�@��9=f�'�tsU=�FP�$��<�<�P�ƣ6<0�Y, =?���� <��D<���C�f=tj<!�9<|%)=~8��3m�<m�<���=	�9=k/�n�9��q4�(�	=s2��x�<�l�9O�6=P/7=[���:�\�Z�ez=�D<�k=Ə_=а<�0v<���كr�&�9=��; 9c=f.5��A��={���3�Or�<��r�p�^�<�趼?\���K�u4���=e��<T�D=`�m�^=k���ڝ<n�
�?����x�@d�<�n�W���ݼ�Ǝ<-];=;�=\ه<ؚs���==N�����=�id=�x��^�m�@PE=Α;UKn�O'J=�6�<
�d��:���u�l<�	�%���O�`S�9F��<�开Fһ� �<RU�����<�=(Z�5-=յd�c�|���=Zp=F7ͼF�9=<��<4�t��<�C��==��:��K="����C���*Q�F)�<�ﳼR�=={���F=޳���[.��`�<�&=1I����9�\�%:F��L#�W�E�lig=̱�N�d<b�t=h�*���=��P�̈́g=�C="G�<�2��PDN�%`t��ռdy=P�=c���Z�S�P���6��a3=��Y���׻�Jļj*�|�7=�����+=����_uJ�C��9F;��<Ƈ�;�0�<S��<�J���z\=}t�<�fb��� =�,_:-���B���IX�a�r�}��e ��2���<���<��=2�=\�R=��=�	v�M���j�=�}�<�C
��W='ռ�;�A��<=�=��+<��
=܈g=r�	�е���@"=X�����B���� <��d�\M���L=�����~=	�	���O���<3�㻡�=�{���!<?N<�O0=e���uPI="9=E����Q=��r<�����}@�W=�=�<�Ty=�<^�B<}r(�Z� =��"��3@=ƕ�3�O=�B������M=�?4<+�=���<�椼�	��:<<�T�;�^6=�y=EKW��ʼ�"�����^=ֈ6=�z;�A|���
�b�պaV7= ��<�Kq=5�ʼ� �����5���=F��"�.׻�U9����6��{'�<!_r=|�6=`z� &�<���<�?�;L��#�<~�s������v�û��N7���)�|hY��^;�=��<R��<�Q���;;��;����5���  <��=Ƭ�<Y-`��Yn�E��������ֆ㼗�w<:���N7=�.?���.���P�G�O=�s"=�Y=~v<���ZҲ��1K=ۤ=�AJ���y=��uJ)<�B�<��;�л</I3:X�'g=���=��z����;Tw=|�H=^n<��=��(<��s� >R=`��=��C<i�<b+A�d��<a��}�5=�v*��"�a�[/�<��K<�����'����m�����>�=:"��6��`)>�����/҃���0<H-�<��O=M�'=��� (=�7
=h�E=#'�;K�%	�<�����G=k�
�: ��<.=�;q<&b=0=����<@�.�X;�����U�<!Yk<+Q�a{f:�-i=C�=��=�Q
�`G��+~V=�=aO�<���#J<�����K�I�:=�?
=�8m=td��5�l���P<0�B�"�=Pn�<�!@=9�H�`aS<�9��a��6���q2=YK]=���k�ch�;`[����=�i}=�c��9H<�5 <66=�9+���9=��(=W=��B�&}�;i5�=f��V���p��[q����޼?1¼��+���ܺp�4=9n��	3ļG�<�=7Ҷ�;�_=�?
�o�_�R�s�{%/��q;�6�r�U=2�=5 a=+漑�w�� ���d=E7꼭�����r��l5�S��<�Z��������,=WD:��"��/=��%���=<��x�!v�<B�׺��������K��O�/O�<L6�;�:�X�\����k�Y����C��M�<��м�nb=g�=S����4)=�p9=�C�Hh��a�=�=��޺��������#S�^=�6ż��<���������Z=lԎ���C�kW_��8&�2�B����<v�ʹo�+=2�Ի_�h=O0V=�n=RQ��	���B2�|v�+��<�y=�1�<_2!�7�=z-�G���H~��7���j=yV�<KIl�_� ���Z=��������
=�2/�q�7=`�=!f���g^����:�=��oW��c�<�KW�ڠ���J�� ��v�<�N=���<�h�t�"�祗<�I�"Y����)�֬-��A���<P=So0��s_�4!k�䫫<�/�;�/Z���O�U�@�I�<C}��=P�D�'qk=S�U���E���A~G��n����<1��Չ^�l�;	S���S<�(;:�;z"��E��ty=��?�bO�ydB���<�E��<���<����f��4�"�N;��;8��<	�������ͺ��wx��(�<I'�<_=�|���* �N���~�<���Q�L<�D<���<m*=D5=�|N�^a='=���`�μ��A<�(ʻ��g=�ʘ��#�<�[J;��v�z�̺m�^=�fO����<��=sX>=�P='D
=?6^=�I�;�������>�'w8:!���ˣ</�g����<mQ =�;��q��;=��'=�)�����OG<�`:�-�M=&�G=�o�=!.�x�V�J�^<Ut=�-��!μ�3�O�,���6�X<G%�Ɖ.=��=���<{`(=���S_�R��?Ӭ��p<�և��or;C&��ֺ=y���_��aϻf=&t"�ۉ=NGc=q�=%JA=x�� e���W=1@);�F��g�:g�<�c=�^=��r��P=Ayb�6zy�w8���=7��$�:�1�<ҽ��0���8�:U��<E��:CO#��4b�>�A��e�<�U=G�#�wD�ͽ<�WI<DP�:J���<����V�`��eI8=yxm�!%m<m�<~@3=�%߻�d!=W0.=�+�=�=fk=y"��9�;��/��F�=�A=����z���t=B�=,b�=�	S�Myh<<5������gy<>�Q=7@b��KּX]V=*�ڼ�i�(�/=0��pЦ<���
C=V���J<Y�=��<�|�<[�=𔪻�d#=2w3�ҶN�@�X�+�=��B�L*9=�N<�Hv���"=�:�<�	9=���<ZVo<X6=�fw���μc5.=�<X�m�p�=��K�"�< =��F=b3�hr��o�;�1<��}�K�}��0Լ��;�4�w�e<1���<}�;�v������sʻD��C�ϼ�/A��}b<P�Ӓʼ��S�b�)�U[T=�L!=_<=$��<��8)P<�߼���N=k+V���P=V�U��r8�B!��[ژ�a<�b��0=�-[��_0=�(�T2=G�+�G)�<,!=|2��N�;=G'=j�]=3�;=p�0�'K<a,����T���e;a���$���c�9�c��w	=*��-(��kg=�:ػT�A��>n=�⼲�-Y$;5�@��<�輔2=���>X���Q��Z=�?�B��<� V=�{��?��<���<߯<���)<5�v�~{��R����l$�1{{�A�c=W�y=��P=��G����;�L=U�{����<C4(=���=G��hs=�̋�?=���<GG'�Z}a�S�B=bD�%S漁�E7��C%=���<08�=�E�<��+��m�<�PJ�^<�<�z��	�<!(�<6j����;5�
��c�<h{���U|<'Z�f.=&����
.�!�|�9�V�X�p:r��U.�;y	=g�(=Ps%=�u�=5����qtD=�5�;�=ӏ�*~)��	=4p�<_o=#.*�l|X;�9�1-����<�좻��><?S#=�p;��V=���:q\���߼

p=H$�<�f��	<���U�l�ƼF=�x�Y�żۇ>=���<�=�d�� ɻ�!��<&��;2@�����<��<�,+<�?:=(i��y똼�S�<"Y<'�<,��	�x�P�R��'o�L�� �<�y׼�:9�^�����F�����:ϻ))��A�ۻ��S=!�<���<��Q��<k�_=����@f=�>6=��"��s�<�,)��0|=�f%=����=���S�d�!�ļ���<�e�<�����ȼ��<�Y	�;�2�qt�;�E���=R<��<}7��D"��8H=�_;7h�p���]i;X�q��B=L)=��"���o=�Y�����T����ܼ�n��A�< �^�SP��QL����:�r3=w��<w�@=H,��|�
��B�a�4�|�Y��=�h=,}]���4� �<��j���Z�<�im<��<���<&/ �m�N�G�8�F��Jo<�x�<�
�=tr3<��!�p���$�y">=x�i���&�=��F�%<t|��^�<��%��"b=�>�=�m�1�}��<�<�N2=O�<�B=#�=�μ���<�i�<�|�?/F��r��i���uC=�^J<�h�;&f�!@=c�4��m=�ac���	��{�<����M�khۼ�H��r�K(Q���W=�5����ͼ���~,|=�eR<�FE=���2����G=jHH=�rS=��G=1ƅ�O	=��5���<q
X��a[=�`��&.='�<L�P<n�%��c<S�;�8e����<w�R�f�=<d�L^y��+�@_=qV���[ڼ�(-=�u�g'=�?-��I��-uQ�G�׻��.=�1'������j�����<51=��N<5�߻�D+=IS$=��=+�X�us�<��6=Om3<ϑ;�k���.��[�Y^*=e$�/p<�e��;����?�;���]\�<\j�{\]���
�)�1<�G׼��=��9>�DҼ�>'��Cw��o=.De<N)V�TҼ�3��l����⥼���E$�6�<��3=�R=�9=}���2�F=<#��	=���<��<ԀA�0�<^�;��ػ��<�08=L,v=�l��=���;�B���n;��r���P=Y���TZ=�#�;uR��b���l�<n=��=<-�<ɥB���껀NA=�|{=@�J�Kz<n��;��K�+_s��)?=;�R=i��<�h��F�U=��S=��=�eX��� =p��= ����=f��<>0�<��=����s�ܼ9ą;��=Z�+�u��+ii=���<����IQ=��<��@=�VT=;�D<�D�=�h�;�;̰<Y鈽p%���+�s;�������<�[R�y#�<
�L��g�=hcq=vS�s��<�~+=T���ܺ���q=	у=�W�<�� �T�<=*+�O���LA��_r;�I=''P�$P�lф��?W=\�x;G��9���R,��B����=H�2<�/�<o�T<�p��3=V�H��4<'��<��Y=�(�<���;C�Y<�c��I����< ��<�,���nV:,������	W=��*�<��R�43��+���Ҽ�$�<|=N�k����<�����s�;�=����݆��J��/;�:����,�<5��%@���^�g�;�A[=>�4=i@=a�>=$�6=U =�Ù�S\�G�=2���Ħ<�����<%��c��;k�8<e����8=E�Q���1��6Q��UO<u�����==6zd��M���;�<�o�υ�<�S���AI=dqd��:�	�</�=��(=qN�;�$��(���"0��Wƺ�¼R��=V\:�.�:�3�\�=11�;`�ɻF�<0tu:�u�$,�ho���ͼ�{O���;�f�<m �<�$*�%t]��/3;*S<9VL=V�<':={�9�v<��q=u�B9�i=W�����W�<Q��<#�[�)��;`�=��2�fർ;7�</c�f���C�U�Ǽ]-=I޽<�eL�G<<X	3��0����<�4�����@�T��<u��<�C���Y�xf=��>�Ui�v[�;_z��-��;�d:��V�>�5<�g��;=<�b0<�I��^r�<�H���z�4����b�>o=��$=�J|=wb=�G�<(8=`�<�a����J=CU����H�O7�輔�J���4�3���<��!=�J�;���<@��<㱟<����+7#=zlX;f\G;������<[��h]��Ȕ�<�᡼�����B=�!���=/$�`�B=�|�<��=x�#��:�=��a��[e�i�,��MK<
��-�:�1�:=�hb<�)�;����v=H�Q=��`<]f=Ux�<g+�J��$�
�»l��/��{��<kA=M��<�E�;/e����4���F�9gs<��}��� ���<Qz��)���&�<kU�<��μz`;,����K=cM<�.c=K�R<�t=aJl��π<Ӈ��@j<<Kx<x 5=N�n=x<�J�{<cn�;{tX������<A�7��[\��`����s�==�i=����ļ�+��'D=/&&�s��:OK<)|��U!��LF%�NW�Cf�<y,�<�;�Lrs��j={l=�#9��p����<N�����?=�Q=��ʼ©=��<�����=��򼯶��T�o�-��.�lK=d�J�4��<!���张<�G)<�0��^�<��<6�#=�M�ƶ0=��-=� ��&�;�5�<N���|z*<�����7=���<q�+��.��M;�;D��<�.�;$�Oe��OV������<�:������(=���6=�Id�Ϸ�s��<��#=��=[M�=Q+ȼt�ͼ��<w .�� <�u==UJ<����
���<g����d��ss=/��H9���D="05��6��pp�������S��F�є��2�<B =�q=Z2��N�˼-�k�����}����;��<�;]	=~G�<��(���=s䥼��<�ռ>]�;�H#�"�=b�+�X�U�tZC�]�<�_3=пT=��M<؝i<������=\$���W=��<u���d	�=#|�<.�B=��=�2ڼU�¼\��<�[=H�h,=�w�<��J=(e3�'��<�%T<80��<���<c�d=�<T=d� �\�<,�ļ��<�3��MP=*�'�	�����<��< r�ȩ�=��;<ǡ%<D	�:�E;P�;��������=;v.�+l(�ñ<[���[=z����<Z�=�,=��9<�ZI�Hi��E�2��=yU%��üF�˼�&=�]�2�ӌ߼E�b=k�;�s#=�48=�D�O�b<�|b=浼�C=;�	�AeǼ��J=ְ.=�_3�1����T�ٔ�<M �w��;��<=B�I�YiY=nAh����<�=�M�<�k$� �B�e=!�<���<��<�z� qF��͏�/��<����v[V�|%�<ݤ_=�[��N�C���;�$=�Th<�����}���ؼ0�=eB��k;ժB=dK�<�`�a�����<h4�F�<\&��$=���qI�<� =�"1<�_��rk�g�>����m�~!=ǂJ<=s����=]Y=d�����~<�%?��׼	#��p=b�[�5{�<uu��o ��+"�iZ�;���J���=�L~;�l(=2�;q[8�C�;g�/=M�o<
k�;���<'�'����9h�C=��^=Ar���<M1,=��5��qW���y�l]��&��<���H���J��)= dO�M��<��=��U�������?��񏽄k<Xu������0�!<x�=8;l����<P�L���!<62<��c<Coo=!T��'&=S����ɼd��<w�X��==�s�]��<k�1�@�K�!�R=��=�;�z�D<�-��ۮH=�=�$�<
�C<H��<��<��<=OC�<>�=�[B=��g<E�B=��6<�;���<�2�'(<��<�ü�0Z;b�=H�s<R�t<�=����n=��{<l�� &0��ৼƜj�=�<)�<�[������<k��<v��:Y�7<��^���S���7=����x4[��@Y�[�<=���<�UJ��b\���=����<�d~=�<+=����L�R��a�{��8B=�+�SI-������ʻ!$�<K����;�=�<��<S㯼����a=	����<5����޵<'�1=ŉ��&yd���8��=�ؿO�䮴<y�8=;(#���<��<{O=+�v<�cn<��u<ܪ����A=�<.<z��;ڈR�缼��<�F�<��c�n"���Z@="�=���n���:���:�=���ׅ<Ǻ��;O\�ө9=ݕּ^�C<)o�<�$Q=��)=�."�Í�=��V���<�q#�2N�<�S��V��9�e��μ��M�<��H���r<��\�,���=2� ��"J=*�L��u>���K����!����7�"���Nr<2ԉ:�(��3���<��=���ta=_ I=M���L
��A=�]J=c���j�?��_�7�;����\&��\t�{t�<q�<BN<�7�<�wi������E�i�;D\=�O�)z
��ł�4%�=gd?=o:d=��X;�<��u�	6+=<]a:PwƼ��8<�v���E<��<�FP�c~]=AR�<��o=�Q9=�Ӄ��Y>��/<�U��kH=~�t�c�~��u�E a������/)=��C�tk=p� �:��л)SJ<�{����̼N���Xb<����a�;w�;��������A���}��1u���<�Xg���=-sü�=��=�6\=�3�<��<m �;�$�<�:�M==V=�[+��)ռ٢��3=��;����+=:R;s{�U@�/����[��ڹ���<�q��)���X�IM</�t����<:��=�h
=�,��Y#�Mw�+I�;�iu=+!컫VH�7KԼ́=�Q,=�-j��Z�l���9<����.<�*��QT�xy�:�?=;y����}�< �,��*+<�`~< $�C�m<Ɂ��</y����w�A�3r]<�<=��^�^������-�e��*5=�j<[8��>kv=��[=�r�cF�;�	=[hG�I�ȻC	�<��V��l$=A�3;���<��S=j��;���<��@��ޠ��8=�<
<�q<���<��<�����ļ(J=�	���k������<��S=֝=�H�����{���#{Z=���<�e��� <q��VX�=`"3���*����<��껠̀=��^=�=�<�=Eт��Mܻ~�h;^��<�z}=[����Ѱ<�A漀�M=/+=z��������<���(����<��=,W�#�6�u.;�Ѓ=N�)�G�9�!U�S���x?�<�M�<M��FY=��Q�󆾺���=4�9=�K��v)=ÙH�E�Ӽ���koi=d�<��	<�o=GN=��;��@�܆�<,B�d�h�ʌ�<�Ȟ���=�#�<y�J=�Dz�4�=��=�8��Xe<����*˼�����,<4PG<H����Yb<�K��K�:H�X�Z�*<qi��[=�A�;��b�i��y<�y��I=U��6�R<�w���,=��B��Љ =<DW��r&=.;y=�0&��͂=�=��4��vV=�I>�%�h��E����=��=u%<x�=�9��=w>���:��1�P}< �O�SlP;��\�kU�<kR9�Y�W<�����tܺ)�$=��<��=G��<���<��i����7P�<��"�k\�n~�;�c�<!z;���<�3a=�=������;��=EU�<��ʼQ[L=��;=�]=n<=ƺ��7&<~�����/=��<��A�|�7�^�����A<�����'=�7�</���h�J��z�y-=$�S�xSV=�z��Rr��
<nf��b"�h;��x��:���ѵ�7�<�5fq������� ;vЙ;�!=�{ʻ�0s<��a�)Z�O�C=W0�<`)a�'�C=w�=(t���"𼞦�:�f=�%%=�8"=�Rl<�;<
����W<"�=';?�G��Y�<v�<RLE<5�1���u�nI�<	� =' ��4ݼ�z�<�1����_�;��a=�)�2==v��<�h��l8�ʺh=��p��V�<��#=��D���<>�2=b�9=]�f�s�g;��O=�b�D�t
���g<�}u<J�<Ĳg�I7�;��=�=�-�<@R{<x�����Vu���F�d�A=�-<�3=�]=�pż���=�e�;θ<�炽��p�'u�V�$�>����\�|�:=��:=v��<78�::�=�|=������z�7�Y=�i�<a=�=� �@=n��o=�i��#=)�:g���.G��{�;��\=��'=��1�~�^�N�9)̼y����`=ݳ,�`-<� �<����z��4�<%�C<��-�!�<:�<���<��P�ɼg���6<���<����G��]�χ�<�6=�/J�q9�;;��'�_=&<j=�U��i-�=���h�J�ǩ�@�0��[�`�,�>5�c��<X�Լ�^[�g�u��vE��d�H�Q�<>�T=��k;t��>2,��Z����,=�#��Sq0=���<"\_=�A=ȃd;U��<B�=�y=�=�"�¡9=(��C����9)9={s���ك�5��;X;=�Џ<�K=���:a�T�ָs;���5û�q�<�'e�1t$�X�:�ź���,:/=!���'�Q<�&X<ș�<�[���=��\=��";�h���Rϼ���=DeU=��.���$=�%�<�_���Z�<��)�|�W=��d�( 켄D<\��<��(=Ht,���?<
nk=a�=�d=^e)=ح�M λ7�i<�K\=UC�(����h3����{٭8��������)I=�X�<S�=��<��ϼMG�ۣi<Hȸ�n6�<-i&=��<��?/=D��<�]<O4�Θ�����dZ/<����;��D��<n�S����[9;��;�{�RI�;LG=�ț�c�:aI=F���}���.��ԗ�<�=�Q*�b��<�R-�#7��Gk� Z��.�<��2��O�������<���<i�ռ�)��终������<]�)=T������<�k!;�v)�`�Ǽ������jj=��=ߜ=����s��{/<H��;Z�(=L��<�-�����I��<��s$M=�-:��T����6=p*�K����!R�J�^��ۊ��l=������C���<� ̼�����dc���=�M��\O\=�ǫ<�:=k=Ì8�_s8=\;=ݥb;�3����=� =���;�=�]�<�.=)��<��=��R�<v0�h�V���n���ἷ���BS=��~��]N��e(�щ��\=�Lg=�!=�kv;6E���e=
e�U� =撪��g�'9�<=@�0�0<�j8=!O=�J)=�F=���<@���\���/	=4YC<�z�<�Ќ���%�)k�<�B=.���z<��T����:���<�����ƻ�����<�S=A�����%=�y<w7�<~k?�"Uu�]1=�ڈ��1�<'wE���:�H4�z6=,==[�<�z����<�j�t���;�(�����<1�
���;Ѕ(<�'8�{�<���0���IO9��p�����'=?�p+=�[�5y-=߄?=-�=��$=5>Ƽ���Ҽ�I���.!=\.&<��Q�s��<jc��R` �v�׉<=_f�<v��<�\7�))��m~;�O�<=��<��=z�A���D�d?���B<�=2�I��;O}=��=5���v==��"r�!V�==5<����'=0ՙ9 �8=�V_=��>=P�,��r�&� ��i�;��2=
��<��=~� =z�J�s��<z.�=�W3=����0�8=&�=�x���Y:=�z�;$�;�r=[���گ �^X2���=�V�� �BT=:�w=�Z�<bA<�v=с�iE���f��mM��L<�=�ΰ���<+��e�;��<+m�oC=�|'=�Bb=8.�<�ƪ�q�<�� ��L<�0\$=�Uq��e�'���9֡��G�ޭ�=��=�%��D=k��������L���J��H#�f�T=QH=�㖼D;B<��Q=T�=��z=f`�<:μ2��<p��<C�<g��n=�r�<g�#�P���"y��X�c��X��D�-={�i�:���Z���=8�4=�+��߳�<��=i@������㼎b�<�6f�׾F���<C����C?=졍:����y	��=�镼����H={�Z��S%�����fQ�<*�4�B���;Fd,�y����i�����u.=�,;=+=��Z�;G����@��\=e�'=��|<��T�y��<Z�����/AI<�&=��Z=�^��$�;/��;Yjv<��=����#%F��U=~ =��8���v�$<̐�=a��<�<uhq=��5�4�;6fW�iyؼ�ކ��ݖ=zP��Ͳ�� �k�f��<�*F�LU=�0���s#=	H���=�;a2=�<���I�Q�ٻt߮<R1E���h=�׆�d3��M׼���<��z���$���C/�������X=�l�;=/9=n���=��.��K�LX=�j6�Gj�<�ۻ56/<>H�<�b<]�8=�;�=�O��;��м��ռU1޼e�=<��)�n&��_EC�8�<�8<�!y��蒼���<8���;�0=�q+�xR�;"��Rp:�����iP�颼�<ɻk�^�����/�F�#$�b/���t� ,="�4=��M<�f�L!=�52=���:e��=��;=O����<TsD���-<g��,�G=�Ft�6O��zM�<~���g�%��3�<z�#�O�0�hd�9���L�;�7P<��<d�;=7�<��[̼��/=F
d<U�D=F�f�]="�<S��&p����<�+=B��ļA�$=�6����<�=�t=��=dܮ<�/�<H4�0优<���<O<q�<�Ɇ<w% <��6�!�<�<21��MZż�4=ۂ;쳵<�J�;��=HZ(�����2Q=����Ϣ1��;`2ͼ���<
�B��_o=p�<Ś�T�6�D�\��y�:x�M���E�=�;�<K�S�<=�=��'�3���A纳��<_��k�i�,�2�5���s�q@�<n0c=Ψ�<h=ݼ�=�ӆ=���<1,I������1����;��<�<:�f�C�6�7cT�J��:K�=)�/<�*��М�7�:=��L�j0==i��<���>�A�CB��z��F�>=�/=���j�S�Z(ּm�ü�����'�;�hs<�~4�=�z�N,�</��t5�<e�K=��<�=�)*=��
��Mh��b<=ͦ�<E2���=�2��X:$���/=l?�⼹�n5\<��<���;<v�����=��(�Ф=���<�L<R�/�R>��	�k������B=�>��J��FBM�w����<A�o=Q?"�4X`=G�j���E=�RV��ߦ��M=�&h<�*��C
=*��<n����<A啼�u��=�_+=�����i��);�0=��G��?��@|�����ߺrfW=��B<����a�G��%u��J=��W=��k�g�C=o�<aX=łE<|,�<Ǚ<����`<�P�b<q��<��; ����<��Q=hx���<(=�O�<?c=C�q<���-��:���<��<�gT<����$c�7D= Q�<9����4:=�� =:��T��<{A����<���}�;�^8�\<B�I=�6L='�E=�29=+�	�rJ��@��<���߹�<�~������<�h#=��Z2=�m�<�"t;��+��݃<�qd<��<��K=-�N���"=��=@����3=�&e���A<1�$���@���찃������)^�ܵ\���'���7[9=Nh��H�w=�q=A���~k<겖�᳼0&5�T}^�e?=�r2�Oj�����\Gk=HQ=FP��y�Լ��4@�ǯ�<���<y�Y<�O�<�������T<���N����͟<:X;�,�;-/l=���}��<~C����<�l�N*=��g��b,�)5�e���E�U��(���'=�5���=�=IB���W=}d ��'c����<�<�ȼ�S�2�_���'��M��r�0�o��u����;;��J=0:?�{�f= 4�<���W�<g!��b =3Q�<�?��<=�1.=�2��$��<��I�8y=�31�>ּ��<�ǃ<��<��W=B��<q�=��r[��Mr�� �������'t;24;^�������<�>J="n�;Ԍ�����:�-������c>=	w�:>9��/�y�%�l=}Nu8�h��ړ<Qd�� ��f$=�XѼ�T����k�&�=B̵�s�
��8==�@;1��)�"�P%R�4J =���<��'<PP���R=��=�z��gL@��,��Z��� =P�=�E͠<��4=���=��F���?=L�<k�<��=�����F�<JU����.��<>�f<��c=�m���o��E`�z�<Q@\�+���O��<2.`=��i��c��ih���p=�>�d����8�Z<G=�`�<�~H=�@+��{5���0��	�:�ں (=ѓ(=3'=��K=+����L�q<t���ͻ�O=<Qw�����=.y
����<5F�<dŨ��5�|��<z��-�غ�0�;WCӼ&μ �<�Z���	��<ͻl#׼�3I=��=��N���N�@T=4��;Mu�M?�;����j�h�)�!2;m��|���ϸ��z]=Z))=,�%=�z.�{�.=�,%�_V��ЍT�%�j��n?=]��� ��̮Y�yӜ�Vށ=:�q=���n��<�64�k�=s�E����!7��nL��5�<	ᐽ�v�<��p<O�T=�} �m�Z<�j��LH�<}��;�R@=�%�<�����v��l��QȻ�pP=���d�m�K�=��:t�y<�=C����.�=����e�;e�4��V=�v<���; �ۼ���<��ʼu�l��zd<���<Fʎ=-�<h[ȼ	i=��2=:9^=���P߸�����K=�m�W�O��:X=�9��<�V��1��^N=; ����+=�N=��%�D�P���5@��0���O;=<㌼��ѺL�=_�<7�k���R���R<�����<��;��=1���-�=�L`=����.�����^��=�i��bu=�z�98����&���d=���<:=�2��x䁽vW<��4=�e�D�Ǽ�����:�����8=�r&�����k$9<��,=G$=�㦺73^���6=�;<�pJ=�Dn�1� :�,�<�zZ��w�`��If�=�n����==��d��Y���o�;%�(=�0$�-���W6ǻm�=����
��<_�C�Z=,��Xؼ��E=�;�˖=��n<y�<�Էg���i�<����Y�=��Y�wz7<�+=��H=�h:���<�1$=4dZ�6ó;)X=D3Y�:=>4{=/��s�����=M�<�7��w#�-�鼗I�Q�V�4A��z��<+���/�<�,==�t����<Q~�<�Q�/�<��B�pJ0=�0'=���x=S�w�Xҹ�cfļ���<E�/=�`3��֋�G�\�)��T��<U�R���:=2!'�X��A�<#��s�=?��2uҼNS�*ݐ<� �<`�wx=1�8=�b�I&��X+M�f�=��~=����:Y��0�S=f5�g\��L�X�F;�q�;���<����y@׻���<����dd�6�ɼ�౼�|�;�`�<�}�<lcܼKи��삽b��%Un�:h��.Z��T0;�#�;�-c��C�;6Z�<�� mY��9�2޲�E1W�~;@��q0=0��k=W!�=�'��۲�L�#��J$�,_ºÀp<��{�Ǐ�<	a�;46<�DZ��l<T׻ǟ;�.�P�;φ��)J����<,˂=/0��:D=/�A�X�U=a�=ߋ���<�=��<�d!=�5�=e|: Lt;Q���μ��==I�A=���"�j=�/D�!�"��ұ��Q2<�/=d�f=(M�0k/��4=}�7=��m��P��L�Vx<~�;Y�<�R=��/�����<�lC<�
=�#=��p��9=�\�<����5d��З[<��j�bR�m�<P�<%"�� �<����ɛ�
����I(�kۗ<����e�t�D*r��?�0P�d�����!H=-���n%<��}<�p����:{�A=��)��S5=��J<�i1�i=H9P=��d<8����0���n�="[e�GP���n���$	?=ö;t�L��<5A=�w�<��3�m5��K=��=_�;�&����Q�b�)���;e&^�}�=��Ҽ#����l=i��<m^#��U=���<n��<�Ri�ϋ<�k�";�[��%�<P�򼡆�;��P��=k��=߼����U��<��Z�`����n���xn={$%=3=s�˻��.=\$=é#� ��<�����'�k�.\9���"�*����R^=0���U<�h0=�4�`)�<�S=X8%=�)#=F�X��n����$�~�n<�%=}�]=PjK=ˤX�#�2=Z�=t)��_N�;RR�n����9��Y=��[<��<.p��1l=�W����<U�U�m�3;h=
=@G5=��x=����&��y����D�s�O�Ij�<��<�8g=EEؼ��N��<]:B=�<��t=�:�~�<�\�<P�I���6:����U=�@�<��<xA�כ��)�����P���[=R{�`1<��l=Kׂ=��o�"��8����#<ߏ�<T]��Pn�@�A��I�<e(=�\м�4� ����ɼV�+=��<A.2=ꮌ�B�2=�o=pnW���o;�D=�M�[==)^<җu�kE�<T�,:���GD��=��U=���<�r3�Is	=��c=ʝ�<���_��8�<��c7���R�}�(='�<A��;���K�;�ր�$�;E�J=n֧<ݬH��.N�E��;�=p�4=>$=��0�K�q�=޲�� �;IJ�:3L;�/r��|:U=���<e#�<����sH���q;���n����X!=~�<������<�"P=����?;��?F<3H�;}?<k+�<]n�9��)�iO�4Ov�*M�-�;�S&=q܋=�"�\�y<����:=��I��'��l,=�?5<K�O;��*<?��
�!�;�������Z��;±|����<�����d=t�_=�=ެ����fj��Wʼ�(�=���dw<G�=�����'�e
l=��<�+�<V}	=QM�aH=�-ɼ��\�1��`���^���D.=�E;�k<:��<8I~;Η!=n��S	=4*=�q�2:��������¦c�M=��P=# ��~ռ�^��Nb��TN=�g�c�:�g?��cG=ݾ"=&rz����<u�!=s����wZ<��q�����-�<�3m=����T��V�<W+)<V8=6#<�?Q���Լd�+�x(��i�p=>ר�T��;x�<<5���<|1L=Z�ͼ��{��;�� �O�<H��<ϩʼ�V��r3<�S�;5=�������B=9wd�VJ��@��Ӽ�\E=`k���<��%�Ź���c������'=c=#X�"z�U�0=�O<;��<>	�t'=��< �<�|H=���8�̼�B;=G1���I��E���/+=_��;�>u<�*7=!h%=W���N;�ٙ:��R=�dL=�@B�
��<��k�U��;hXB�h�[��Q,���X��F =�C��Ѽ�`h=�} �N��;�X:=��D=���<�4;WXR=��5<�j'����<b�<�*d�L�_<��p=S�9�T��F��Ta��IF�����Bk�f�c='��{�<��ż��P���<����<�lO���I�~[p<��v�B�P��]���$�Ɵw<8��qO����$�_����Լ��<'�=�>+� �m��,��Ͷ���`<�ޥ���r<�j)��I��P��!!=n���o��b���W=�	���;�=6�<�y=q=%N=�7{�!���l<�'���B<=�!�<QSL���1Φ��6�<6W��H�\�fss=Nur=<�=��' w��X=�J�<7�8=U���3�N<H�<�,=/V\����<�J=���<�{p��i=�hH_<�d�8�*=�Ƿ<]: =O�I�3�5=�W��=ŭ=�z\�w�/=h��<�+;�es=5?8�(n'��2��U� ~&=E����N=;�Ӽ���<���<:�p�?U����0��|VG;�T��D=����%�#=Zt�;ޗu:8���8�ݻ5��bLB��Ot<n�[�o���<?�<	1,=I�=��oLh���;�x�0�-�� �����<K���7�<���a�.����;i[B=Z�O=B��=dx�c�Z<�6��W�><�I�=
㗻���<����=�q��R����X[��R"���<^�
�#R׼܍�;��<@���G�C��C�=Β���gM�DX~<�E=%�P=�}����0<��<��Z��_��<!R���T��z#�P?�;�7=E����Y=Y
�C߉=���;�_<=w��K:�o�=I�<�O<2�3=ˏ�J��=+�={��%�;�w2�#K�0���-�o��<��=6���b��i7�ƌ���,Z=&��<L�<���;M�ɻb�4�(�n<^z%=�F:i�=�B>������}_(��DF��+=�|R������<^nm=�RF�"�ռY݃;qC:��kϼ8��a�=od�7hI���ϼm�@=�y;�����=X�����*=.�7���<�;��<�=�	��}���:<��s=�x���RV=��<�UӼ�E;:��=+F'�_Tv�=8��V<P׃�[ɼ�<�8�<�����;�u;�E
F<�b����Y=�ϼ,�=ӫ�b�	=#��;� :�ϰ ����dB!�o+J��<=Vd==�����ܼM���+�<�k4<�My�}Ko<Q�ݻ}$'<�J|�%bܼ�~�B�a�#�M=���<��\=k6��K8�:7�@=�TG=2�?�1#;x�/=�Us���s �<�
`<���<��(�
1�<��<�a��)�d�Q+�Ê;��H�3>Q��e��K��;�P=��B��F���==�
�R�E��-��qe%=�s�<3ټ���;��{��e[=Z-��D��ꬼ�⃻/1�;�����A�M�S=5@��
��SP<bj=];�<������l��<D�`��`<ń	;K��9钮<���<֛
�y`U���H�F��4�Y��{?���;��8=�j��X�<�(���[��_9;_$;]�<<�;��(=�Ga��B�Q�V=�b<�MżäH=�t"=<<�� Ɇ=�ҙn�]F�<o�=�~�<��,��w=�����<��<���<�-��
�<g�<����G=`�g�/�n���<�y=��C=��l����;�lO����;���<M,9��餼'��=3��<ۣͼ�8=��<�vf�Di��O��<�=Ɓ#��֪����8h^�a�<>�z��+P=��i<�=��MB�[%��ϩ���<��<�yI=���<���<Tw�;yl~;�h=�h%=�R�<���ħ_=��=xC=8=�H=sy��s�;�3g;�`�W�o=�>���９ G�a=��ib��tx=�4B���L<�0��F�<-/=��=?=KT��u(;9���<���'�A���R���=(��<�T=��Q�D�=a9=�	z���`=���:�Wh���V���9=�����N����<X�f�R�6=�Y]��
l=�Y=�Ȍ�5�j��%��hм�~Z=���|�A<�(=m�(<r][=�*
�	�v[�:�_�;����F�=����r�<-��<s���	ڻ9�d= �i��!K;u?��j�A��ݎ<���: c�:�)��UO���%=I�<+�d<�Un<Ħ���=��=lT����輑�������'�;;@�.=>v߼-0����j��c�<��<��E=��Ƽ5�@��"�<�==�<��߻:$��Z=��2<�8<n�<\FS��Xü��<=����|�Z�N
�i6����Q�;C�/=-~��5�=�RQ��Vļ�38�;�]���y�a� �*���FP�����d�����+�ĉ"<�\��z����-=��+��6=6="G��T�0�2��=�/�V�W����B.��м��+=��$���<�=�,=Ј���VB=\�E=Ƴ^���h<��G��[�� U<�V<��|��KZ�N�=���<D�=�ڎ�^��;_H��AOh��C-�#���Y
=�7����;f�Q�,cT���<%��<��+=�%�����AX=P�L���<AX�$7�o _��3�<y�:�NU�$q��(g;���\�&W�q��ˉ(�&6��[r�<�1����:��=?����c+;�3J�JN=}�]<�I=g�A�x��:�$��aI=�h�9|g,�'/� ^d=�5='�/;q�����W����GƼ'�ʄ&<�iȼ<|����<
\<+[%=��B=aml���i�A��<$&I=�C?<���\��&=X�7�d��<2�_=���	�=���-Q�<��;�cN�91��V%=��p;`=�R�<��%=��輬�Y<�nؼ���<1�;)���Y@������Qa��nR�T��<ӷG=�n�%�5=�M6�!�G=z�s�g�<�#�<?N�5�%�2������x�:=.j=T=�:��z�<��>����E^D<¯W=��R��[���f{�Ǆ:`�{��i�pU(=�LD=4�E��k��HA�MdV=f�=(��<ԧ<��E���;��&��;k1��LK�u=��|�R��2����+�ԏQ=e��<M���8���(+=FZ��m����o<<�ͤ<z�i=d��Iߐ�z��<����L켮4ѼJ=u��<�q@=DD=,�f���=����&=�mֻ��T
�<ua�=*��t���:g:P=r�=�5=̈́T=1�=�'C:e�X�x��U���"%�3��(�8=�9~�m<�;�Ӎ9�����Ā���;�|E=�R���Y�;��`땼W�*=]w�<�e��Z/���=���<`��;9��<�O�;:y=Vt���i��
�T�B=�ۼ�����6���<^�=/����=��f��Hy����<�b>��V2��7߻q`�m�G;���s[���:h6<�����D��_�<�����y=ڧ=dY�<u{�F���h=�~���A�;%�F�����<qSټ*ܻw,=X<g����<�2�&3��?�c���$=:.�<��;����<�%=^m9=#h=��~<ml=|�s=�S0�zռ��9=�%=H$=(H༟`���<�6�;��=��N��$5=r�=&=�ɦ<��j<c�^=-ּ�w���=��A4<��`�g*����R��A�;���I�*�6P<0H�0�J\.���v<FEC=�S��~S=b'����=`�y=�&<��w��C��v<!D��n\���̰�l3�<�V=.	���H=��N=�N<1���t.3<��E����;���<T��#�м�xT�d.7<2�P=�_��V*<�Y#=t��<_�~�n�G=3��;���;�����;�'=zF=���;E����׼��/=<�:�ؼ������a==V�<�5=��K<	�(���.=?�r�7�=2��x�.��M�<�Ӆ:5�d;*�H����c:<O�<��ٟ��_=<Bo=쿄=�㐼��<��;�=P��N�<. h=튊;�������R��<8)=�ݷ<���=|�<�S�=�>������FN���(<iw�<��=,8�����9<�IK<0����#�<9���<���ǘ�;[�=VӼ�ob=��Լ�ϟ��Kl<a�$�g7ܼ,�=��c*��JR=�Ԍ<_��<��.=���:��8�{?�
�=�= ��"=2�!�]j=Dfлp"=͢�;��0��2F=� 5��CQ�G��;!kx�/g6�#�'=,��SI3���<.{F��c�;��P�C=��ټ�'ּB���}����X�"<;�k�dPU=}X4=�oD;���<�K��F��<����r3�V�
=)�<T�G<��<�̊��I<VM=~$F��O�<����===qм A	�	�=i �<	��;��Ļ�zZ=S�6=CrQ�qJ�=���L�e�V���I��ls=���!�h9�b��M��<F<B�o�=�{n=%��<��P���Լ�@%=��)=˃��-1c��Oh�Q�T=r�=�༐(�;	�$���;x+�S������9�D��=����m���
><���F=��ߧ���:�=��<:U�<�f@���7�B��g�������+=�kl��R;�$E=��+�l`=�$D�<�A����)���0�N���?<2�<@nV=�9=;V�<�7�;��=+�4=�FU=�N-=;�=��W���.<ȃܼZ��<�Ș��Q�A��{ڕ='9м6�;�:�?�<��<^��;��6�����_<_:���+=ʇM=>��SB=<UU�|ф�+�<��ԼY.��(a@=��F9�s-��93��{����.��<��<4^U��] ���<J�?<��=�c���^Y�(5�<�%��f���̛�t��<%��=��a=���<%�O=.
��n�^���u<Ĭ<��=�X=�<����%=�ZR�#�,=�i���0=�fF�뉈;���;@�=�V1��g�u��<�w~�x�<��x��5�gg=Ö�<�-c�Qsq<Tf?���=�&{��К<K$]=g�t=85��ǃ=!�7=C1==	 �E I=�#�c�8=��;;ga=���<��7�K��<�,��]f=�=�*����7�:��<0O<��;�h�<��m==)<�P`=9�[�F�d��!߼ \̻���<[��=n��;�p<?��;k�B;�d����=LR=�=h��=����l���<�,���O ��W2�Ջ���V��A�<ǹN=^N=6#���<=�����=�+=���)�l�pC��@R����x=$���I=��<�噼:M'=3�弯�c=��
��}}=^�/�(�@<��E=��<?.=l�<X6E<�hB����<�/S=��=	"=b*=��!�9��;|\�P ü�`�<<M=�LA�++�<Q�$�:T$���S=󑶼Yr��_4��jռ����˼[��^� �����X�<^F<.X�;����w�<�S��}K�����luK��L=��k<���oI<�x��];}c.�����T�?=���<�;�<�1Y=�<(�9=X�<�ƱI�W��<uz=~Y��oH��R�7=,RF=�v��K����^�<����G伔2<=j�a=��=��(��R�ϼ��<�	���K�j�<�r��Ni�:@��;��l���zIټ�̬<��9���=�����d�={��<�?�bY|��Y=�!I=\֥<��;�p�<5������<�W=��:����?=l��n$=F��<5�;�'��<����F�C�~X�<zzm<�^T=ŕ]<M\=	IM=��:��=�-Ǽb|;�E=N�;I��<Y��<g�<���An1�ay�<0�O�֍d<�i��SG�<fdw���1=������=2�;`'�< 4�<թ#��B��uU�Wn�a{l�3���e��tK��� ���H�B=W=��(=9v=VzQ�BM��**=2-�:�C�<׵X=�.�<�:�r>=�i��i{����R��ϟ��5!���<�C�<������D��\u=*Y>;X�.=%f)���<*�ּ" =p�Q�@Z� *p=Y�g�#ɻ��
=@P=xCe=�BQ=�̻�ӻ��f�<������<yj��<wV����BvR=^�tS컽3���m����<=�hN�7���L<�=�M��[
=�͍���;=�Ҽ�@�b`S���>=�嶼�6�0=�t4=�;�,���?�<6���=F�v�b?7=����L3=S̝<��<=<�_}�&=>+�{&(=�<��!���G=yL�<�7���7���?��N=�:8��E=���<4�=�:�jD�s3Ǽ��N�߶<_��<�,m��0	9؎�<$m0<+O�<��=QH4�Z��<Õ��m+�\	ϼ�}�<ߚ�<��=k9`���;�#%=�}`�2d�<�;��0$���<H��<i�<Zjx=x�-�i���<U��/�˼#9���=@�a��J����G=�<$�e�=��༙X�<�;{:zI,�<�k<���?=4& =@[$��V=���^�.����<Y��<��6�^;=���<f��ǔ=�b
=��=��,<d�:=�qV=��:,P�;y��</�t�9��<�:廵u�<��<;h�ȼ�=��)=~�g=�8=��L:N�1=��j�\�$<Ό<=tm�/"��=�1���=�w*=`��l�� 0���g��:=��i�&Z�ȯ��^G<����P��>��;�
�=�1��E��'���ZL=��;d��������9� =�{<���v*=1�p=D3=rt缉�<z`��i����;��f=��@�������0��u�=�3���En��ҧ����<��Ѽ3f=U=<��@=���,7���=q;8��_�D�G<?=�c�������Z(�<,&S=7E�<mg=�،=��g=���+iK��N�<�����B= T
=�'／N��Sr�<&*=�C���&=�Ի�<�<0]�<Ÿ�;u�s���):dE:���=*P~���;T�L<%�4=��W5�p|w={�*��Mc�,��<Y� �l�����=(cV�%`9=j=S����;ō�<�p.��r@�H�,=��O��n=j�r���<��D���Ȼ����A.=�(a=\�J��ف��?=:逽���G�=�,�2/�=Zh�q�==u�(=��1<��Y�)�f=hd��A�r<;���P"�<N&��H��e�2t$=e�<㌣�@��<TP���=�����x=qwI�Dj�<Bo@�R��8=Ú�<���?=�RV�uz+=�w�<T� ��C ��z=cU�<���+=���<}$��E��	�8<��d�;��<��6��yQ�h�t���f�<�s�<~�G�-Gd�N x�ژ,�J���W�/{���=��<�/�<�R���2<* ='*;��W=�M���D=:,�<F;�<�8R���$=%����<K�==�L�2p4=�7#=:�����Ｚ�<\�>��h��6�M�=��ۼ�Vk<E|�;�z�:�5L=�b=ʪ<ٛV����>9�<
�<Y܃�z/b=�1N=�	<3�I<����[z<I˻&2���m<ba����>=Y�6��Do���b�=D
�<#2��l�<���;&
�<+n���G��^I��o�<�I`�����v�r^���S;��X= �Ҽ=��r���7��%���OA<3�;�	��)�<\��uܼg�n��9�<��:O�<����:�򲻵|�<X��(��<h}6�J9�<6w��|����;�E=gו��-�a?=��0=�8���E �P�l=�^<=�[Z�T:~=[-�;V�g:�y_=�=�I'=�!����<~=��伫�Y�ڬ��@G�j��5"�;i=O~��FH�n�X=��ռ��=I���߰!=�ֻ٬<3�B=I`Q����<�=l�Y��V=�E1=�4n<^kV�x��<�~ڼ��<햼F�<�.<:�==��(=NM�]���=��5��K=mW{;Yr���Db;���<5=��<���<�$%=��,�&8`<XH�<�$�|!��B
�X'=ߞp�}|�<Z�W���0�Z�@�Ȫ`<�ۚ�@�=�RQ=Q���H��<��R� Z�C6 =,,=L�]=�5�3_�����F缠6�<�����m=�&	����6�%�<�)=Kq��w�XJ�`�:[U��iw=[�G��m���d$;����<�* �Q�V=��c�F�LgԼ��&�X~_�udY�C1���滰�8=�-_=��=;��<��@� �i��s��.���Iq�b@Ǽ��=���=Ш�]Β�� �<?y�����<j%=�8�XP�6���~t����^<R�,=b��<3�=�<�샼�(7�6#<|!��S��iY`���U<+d=l�,���>����<��<:P==4��<��<A<� W߼1mA=�щ��Ì��^o=�Z���B��Qr�y�
�V�Լ~�1�:oY<N��N=	�=&<�ds=��3�4�.���<�Ľ:kp�<��=�$�<� T=��+=���<8NR=5a�<Q5�<q�i��!�<ڈ�;��g��/�=���\��Q�=��<|N\=O��<;J=6���=�9ۻ��K�@�/���S�A2�mp�9���B�=�OE;�Z���X=�?�<�S=���;���;Yv�����[=������<Yd\���V��r��� ����߻�z=��J�_�,F�9�¼%�"<r�?=h<t=�O޼�u'���;�<|XO<��*=���<D�ϼCG=�ںM�<��I<��&=�%��|�<t��<!@���=qb�<����1x<���=�6;d���������<��>�6! =��0�8	f�D
$���;��<�5�<#�����<e�<��}<%ޑ����;z�<ٹ�<( ׼�y�9=�V�ꦅ;H�5=������M����u��V�<K��;���M!=�w��G�=��i�qf�[�B��_�; �=eR,=?�;H���O��0!=�-.=�R.=�|<!jM����<CP=<i)4=qy��`F=g� ��ἆfJ=>��<���<V�<�0c���'9|!#�� K=
q0=0��<���<���<�Ҵ<�y2=.5<�l~�A�m=�2=K31�
0����&�K�`�<Bѳ�{�C�Z�9=6Y��$7=�-=��y=�Q���8����<�zd<��I�-I��"<��#�7_o���;���9=d@:�t��=b�
V�=N�=�Kܼ���<���Ĺ%��B=��=���.�P
�<�|��<h�<r�m=���A张�Z��<�v<~=��Z=���<�k����=v@S����='��x<�� ���E�!(=5�Y�=�;{"=�3e��-7<Vaټ��[=�;v��c�E�\�@6=v����~�8/�$_׻;�K�V=���<��N=8�M=r"��%}=�F��)=~e���
=�0���>�\�<L�¼"�@=�FG=�3.�G�u<`\Z��*�0=8V<Xڻc5.=nKW�%�����=�=Pf�<ONb<|k=�9==�t=]4���|M��d��������S8�n~;VH=��<�+[�
5�;�-J<�jJ�y�*����=k�=��C�r�:���:�v�<��:!!�<*3�<>z�<�K'=��:��~��)=u�Z�3�X�.���-�<������<In���S=��J<�wk=5	�<k
-=��~�̄�<�O��L��<ƸF��N����,=���:)��<�Yӻx=�Z/3��Q��|7=8�4='E���*��<��@��м�$"���N:F�A���O�~R�I��+*����;�~��J������Ea=0o�V�!=��"�39}<�3=+�|��ߟ�TH=v,<<D-=D�<)B=o[j�J]Q=_~���=k|�;C#H����<��K�\��<Of�<�,=:u�=\��<Hj���<[;X<¦G�hw�=:y��B0�<��D�!�<E��#;�g:$��(
=�𙽆�H<�Eh�u =�m��h	/=�L��)�J=��%=x�=�@�:�)�L�:�R=1Y�<��	�0��.��+
����<+�ڻ�Fn=��c=��w=p <����$��u@���z<�7�\�D=���)�1(������v�<D:�<J��<���#�C=&=nh<� v<�Y/���s��#���O=�o=-d��iф�[�_=g�G����<���*�~�5=$GF�����d<6�?���d���l;��?=�u�x4��8��/�G7����Y������
��&c2;D�<>+�;����~/���U�S�;=� G=��<_��;�a<6��b�<�g��
=��r��0����9�U'0��,�z=���<^7��V//�Ŝ=]��<�#ټI�y=��`��q�<�T}��5漽�o�{Z=*����.=�_W=�1=%,=q�n<�t�<��=��G<�: =sy�=]�h���=>���#���=�-��Ԅ<�wQ=��=�I(=�6@���s���-���r<;҉;������<��P��aSt=�k0��8�;�[D=J�ż�9N<�o��d�A�ܸM=_/e�7�Y����<��Q=�I�(w<�����٩;�RW<��<���<V����C�K6��`P=6kw=;=#��=p1��x�X}��i-��N�����pZ=I�5=BW=)�:fH=���:���<���q;2;�k����Hv̹W�M��<�Ys)=&«<�o�=!�K=EW���p2=�5ڼx/`;x�E�w��<E. =T׺��\�� U=;��<t��~5����*�x)�<�&{�
�����<�!=Vo�4Y=��X�<+@��2��Z��<Nv����<�q̼�k7�a�w���T����� ���I=���<m�q���!�g�<��߼{�9<f[����F=evm�G?8<N&�����E���Jj����<�;�<B�)Q3=��j=(<���*t.�ڮ-��C=�)�<�憻;�<gE<��U=��ǹTeڼp�<�<��i��uF�w�ź��𔩼����<+='�<�"`��P��=�>=-�R<���Q?�<@g��r=�o�<W=�z<��R<^��� =`G3�8��;�偼�b2������Sl��H<�ǡ��BL=4,��q^E��6����=�P-=�G�VJ�;�[<!�3;�ƫ<g�<�2E�'�-=4_L��x���8�~�}����=%��d��?*=Ne�s��W��,I=Є
�e\=R(����<����{Ż������;�$^=
W=��R=}폼u<�R���;=�		<�#*=}>t=�@q=B�:�
=*z=+�����<y��|�0=u��G��������]�r�< ��<�=}��`��"��p���@��(�f=������I�J�X=��;�"j��ǼT
x<��,=���<��+��,<�@`�.Un=F$o<-��]����;��=��K�; �v�}�=�b�;Ra��3�=�~?=�Sʼ�	�:>����G`<7y���<��q�S���V�P7=#�7���i=ȉڼ�.=��)�y�׼Sf�<U���=��=�c��̰�<<�K=�A1�2l�@Y�<Ϙ=뛊��F	=�#;ۋ��B!�w�<AX�<*�<�b���0ʼjk�j�`�'z*��y���};�u3= u5�5%��q
V<�j=�C=R�&;����7ɼ�rN�%��<�!�����<3[�U9R�9hI���#=����C�'�	D��]��drU�!y��!�<3�<]-;K�=��r�.;_VԼс6:�0��;*=���<��<�#=�1��s��:���;p`�VE=���<��cOB��=���s���B=��;�k�.�Z��F;��r�;�漮j�<�ф�6.2�7Od�jZ%=�RT=���;�A3=,Y$=��[="�<�
����<"� =��0��@߼���<=��<}��f6p��5��KG����<��ؼɊ=����pӁ��b=@��<婆�?}�<:��<9A=�Ї�厬��=��5�=eǃ�uּ݀�<K�@=zW<8���qfy���<���=��n=�8M=��f=�/;ߧ�<�[������|G<W
==�� ;6f�>�m�C���6=n�=#<s���ř;�/ؼq�=a�<��/�Ұ9<�b=�~=.܄�>Q��`r;ʽ=-d�-L+=M'L���<�68��Qj=Y�<^=���E%�<�=��=��+�;��:�`}��xW<7}!�tT�<y���&��[1=��*=x�;ئ;=\8l�BF����(��T�=�Z��D��f>&�=t��<T쏼�1�8)=:,���������ȼVU�;}�o����~�u� ���r=iR9=�$t=��{<����0�
��NѼ�x�<��M=ΈG��4��Z-�ه�;��[=�Mh�M��<,!=��R�v�3;Х^=�U����<g�<�օ��\T=q�D=�qȼ���;M�q��8�;����Lg޼m>�7D��z�<�2*=�g�<�.��x�=l�<$��7$��0��� �Y)X<�B=�x��S=3����!<��&�@!�Ɇ4<�ru=�ü�u=�<��d=h� �f��󼥯<H�=�:q6�<��=�bJ���.8Q�x���]<D��<��;�,��|���1=颌���=�`�<&��<z�59�^(��=p�(�8�a�m��ņ�0Q��1�P�=ٵ���)==��q)j���;=1V�<�N����0��|z=��~�yX@=ʀ�9�Iu=��+�{���-�м�����B����;�&�<�/%<R�k�D�<4e5����<p..=
"=�F��B<��i��B;=�@=0/�<�Y<�!�-���p�;�X���bC<��	=.�A��Q?���t�
s�������x<m��=(:=�Sn��ӌ<��f=�;ɚ*=x�>=�x��*��a[|=�D�6bK=��p�!h��
@�<��%�w�0<��E;>J�Z�n�<��<Jʈ�5�?���/wE�m�0=�N�=������=���<V:=+_�<��0=��Ѽ�C���1<�Q<�A=�%�<��%=��?��&<K�<��*��<�<x<[�`=~��<����<G�v<)R=�r�<ݸ_���<#����J���8=�'���=
;|>�<;{N���o�3��;"�D�X���0��O?��v;u�/�^#����k=�v�\�X�����Ι�7�t=8�<�>p=�	��K�| e;RU�<m=�����׼�#G=���;���<�A��#=q^���QE���)=*�9�IV��MQ!<X_|=j!!�᝻�<�Dؼ���H�H�=�Z���= E=��<�弖~c��Ӽ �< ��g<e�:�N(���물Q�^�n�=�W=oP;��~���ϼ����l9d���f=7x
=\e��c=�5=��V<��T��;/������m=�Ⓕ���;]P�<i�Ȼ��<�����
��a'� ��<%�G=l�=ja�7����r���$=w@�U�u=�,���%'��5k<J	=�:(<�W���=��=Q�]��X�<ǐ=~c<z-;<\9�м�;��=�H��'=/+3�^6�������żi�����U��u�<!L<	NQ=�
鸜�<��`��_8�}�"hE�%�9=	 �Z�1=mW���^=I��<���+�߼-Y9��5.��Õ�ڜ��(u�<Ԝ(<� �;Z�c<�|3�υ����t�:G� ��᯼�IF��C��ރ<�x��`����F�"%8���<"@��ֶ<�wؼ��k�YԼXZ9=�-9���*=$�<A������=�)z=��J=0A�<Ln�+�
�=�ϼ�N�<6��cY=Ro���ܼ��d�X���K�<��\�\�<����,ϼ��ü�>~<�ܼG���2�@��q��<린<>D�<+�=�n��-$�0�=j�A=��ּ!4n=}m�<	�=	��<�툽��R��QлW�y��D=��b<��[<%l<�d(<>���2��I=��<F���w�}�D=���;i,��O���l�L�M���D�kWD�s �װ�<�Uf<���;_���(�W�/�_a�<����$t;Q�<��z=A�A<���<y��ó ���ݻ��޼Nk���>�=Z����'5�I�R�6q����O='�C����;K^*<GH�<�[8<
=3��$���=t�R<��-<(�<���S3!����<A��<5,�8�f���<W�m<�(.��ȕ�fee<Ԓ\����<v�.=t���	A=���W��<>�=���<���<��=��=��)���L��J=#=,�==a�.�|�>��W�!%伭`l��A ��n�<�I=M-�zf�<d����FH���d�ß�;a��<�!u�c������=IW�di�9k{5=��F=:�_�\�
=��=#�;���;ud���<��Q����<MC�� �z��}�=�= �<�������<�X
=�|�����<w?��Kq< j��=<=?��<)��;��纛�C=І����t�
�����7���F�L=B
/���3=]y˼�]C�y/��O�*�w�#�W="_*�M�q=�e�`�S=���<�(�<�����R=m=>=M�<�I��=��<��kuǻ�?=<��N<�u�D����T={/7=mB�<0�P=
���<�L<ms��+�1�5��<��(��़�[-=^�;4�=�i�<:����"�P�<$��[��L[=Z�<�5*��?3����.�}X��7��F=���<�s�֕]�i#l�-�����<��i�4-�+/= ��<�`��ߒ<9�n�?V=�ɻ}�X=J#@=�;N��?=�u���b=pt��C�����,�ļ�mN�%Đ��D������<��=��=� �:h����S=����lP=�ّ<���<B=l3��|wl�*j��@�	=���<��ƾ�ؑ�:���<�L�<��0�,�	=�W��%�;�����<Y���@���J���r<Xl�;e��<��<1j[=Z�&�u�0=N�3=��<k�9=+��`���<=���<(K�<v�<ؙ�;��1�<��=�h�< i�<�3P������YU�y�{�ᤙ���Z�Y=��Y=���<�?<�F���s�=��<��f���o<�fE���3=~�<�!��!Ứ�.<�9k=x�v�]&�}�;
�U=^�'���g=�<<�+=�`==��f�Q��;Q�<���ţ<��� +.��@�<H�a��
;��qv��Rs=L`(�81i�Ca�<*�H=#�=�Dx;#���/�;��O�j�=p뛼�RZ�ef�������"�yS!=N<�<t"<��<�:h=~�Y�aR�G���D8<�E*���$=Zm�;�G�=9#�;T�<�}���qL��?7=ӳt=�Hc=�G �n�ƻ�E�[[���\��N-� &�v�w�=��<[�};��"��\=>=�:��<�಻6�i<�.=�xU��2v�D�=|�/=�Ҽ���B��<$�w<�!J=��o=��S<7��< ����3�:�S�<]��<��N=o(��j$=-�c<g�<���s�۽�<[@�;� *����+��0�(���-���:#�E=�	u=�<���;=��;6P=���� =��<V~��\H=�~S��{缱����5��,I������p�;%7=�
�<.5,=�U�<.6�<w�����;�=Bu�2��<y�S�;W���!��>c=r)���2=>8=pUּ����W=6�4<�W=5~*�^�2�	\<VG��s� =��.<�A$��;���<!M�;4�6=xL��
q��F:;��~<D�'=jy<�.%=y<�ټ��m�}��<;��<�@C=C�U���ѼI*=�R[�f(����xO��7�=X���
:a��x1a�F=�m;{u���T=Ma@;8p����n=��;g�=7u�<�&���<F�`<�#;�iwS=�μ��;s�jx =�k9=�����`�<�L=�d�;�>;�/"����;���ZP1=��X��7�WJ-=_\a=f�$=ĭ�"�'=![^=%�]=�t=�׻G%7=nH=s0<<��<�?=��i:U�J=ɧ6;e>����=��O4=f��<�����1H=��i���6����BV��A(�;�ۻp�<UΦ<�)����1=��:�%%=#�=|��<4��< ���.�[��U��\z=P����#��H��o�d=f�<
���Dۼ�<���'�J��}Y��N*;@稼�.<�"5��u<w���f���r�3�G��D=�Nȼ�˼��=��=�w����;�wk=�S_<�x��M
�j����6 �|#m=���<�4<#P�<|T/;�ƺ{�=
�v;Z_���]=�
R=��$�Aﯼ�+����ټ��<O&ؼ� �;^I=9��hZ��w��CY��1>��+4=<����<�qJ�Ú;6.-�d�6=~cE=��[��z��U�<(��T�A�YTV={ֿ;��<��=:F�(B=er�<q�C�Y</�'=�ۧ<*O+="�@=4oP=;��;��6=[I�ڗؼ�N=Wtc��=(��(7��+='�}�6=��=v�ּ]h�;���;,�m;��?<���<6<�?6�}��<�^g='�>=]Z�<���<�s<�����_C=]�q<R[ݼ�X���$=9��V�<�������=D�J���N��=�=�1�<�{R��@f=#==��[�d9�<^R<�o=���� ����T�O=˂��a+��_�<�,Ƽ�K�ʺ�
zd�X���<�U�$=YF;@�q�X=H�c=��<*=ۼ��	��N=u��@�	)'=:)</��<�}S�����$������"�KMI� «���:�
����>0;=%;<���<��!���;�M��h]9����g|�9ݑ<�N=��.�?�8=�2c�0�-=�͠�o�=\�<��V=[[@< #s�.�b��N�<�ۃ;�t'�>=/`m���`���=1t=�W/=����f��"=�?���;v�=��4<:��;vx��h�<�Z��w�]�=�C=Ff�����Qv�K�0��h#=�v<�^�<��(��Y켍���*�x:~���VV={׼��Y{F=�#�*��<o� =�VI=ι[�7 ��@��pS�<�~)=tY=�o�q�p���߼�=7Ey�{D�E�(�p�ݼ��1�:=b;��F7;��}<�΃<�&O�M�K=^�Y�u^˼5:<^V��W箼c:ռ4Nw����>~��ƼG�%=��=z96<��|=�����i��
��)=7D=��<�(�<F,�<ٔ���u;0E#<���<
��<�)�<m����S�8��<-|<)�=�o꼢��;�<[6�<�X�<���<U�;-x�<bq'��G(=9j��K$=����һ�{�<W��a:=�lK��:ʼ싪<��Q=��:�#_�;��ʼU��<\�(���I=�|�<��;��H=�Y)��o�N����\�0=n%=K��<Q@L=�.)=j`-�"閼�.i��n�<�ƈ��UU=<=s�i��DƼd���������)E��͑;�罼��<E�=��]��I�<�R�;Vw;W��<�[;��j=�����G=sD<\�6��3S<���|ܼ���<ҕ�<�q�<I���9��j�����:aI=+¼)�J="p2��gѼ��!�Ws�<�`b������h%=�(=���;]8����8R��v
���g=7&��m�;ԯG=i
����:ma=���S�<��Q<��=XZL=6�$<���<;=�	߼������)�J�;���<�V���5��!�;�L�<�)���<��u�������X�u=��<,Zʻ���<(&k=C��<�����-
=�8=&�Q=~�O=�f�<�z`<E�=��"��M߼t\Z=��w�c
9=�N�;�����M���(;��#��GF<M�:�a����<��:�x<3]�;��0����������]������IE��jh=��s�O�<��8<p $��;Ѽ ���d����%��<=�Z�<"�d�8w���"=)��<_�M=dQ,�8ӈ�bw�< v=HB�}B<!�e:��|�e�^=�"�Oܧ<�"�<z�>��^=-�a�<^[
<�e=L�=�p���V���λܡѼ��B����;Je1<yA_=���Յ�`#��i<��T�T#�˞�~,9<�H ��
!��~���|w=r�e=��=��[�,=�T��$!��P>����9�=:��<>Pp=u��:�[�[ُ�sM�Ǧ �ҁ传�b=)�r<�B�<o�Y<���;��=�(�<�<��e==�U��'�<[	=O�=��ׄ<��;R�+=��<?:u�r�Z=��^����<~[�<x�V=$,�e��;Ș��7�:̉�<(��B�5=��e<�F=[G<Mt��3b�<�0+��� ��%�8��(e<6�h��:�<�뙼E��ž��=p��<0C<���ٳE��{A=�K<Ƞ������c<\��u8�<,jU�ϣ����p�����)8=��:jS�<K�(��e%��)�����<e�[8��,���I=��;� ��=�>=a2A=e�s<H���~��<�0Y��f�<>�=J�Ӽxd=c����]K��L ��?�;f�;I���,����<�1�=�$�<Gc�|�(<|�P��==�9<y�;��������M� �D>�Ʌ�<\Z�;~<�e�;�i�<=:��eB���͡<_��;\�f�-Z:�ܚ< I=)��<�qȼ݌�<�VJ����\7&<Z�<�]f��~>��;ܶ^���÷<'=s~��zV<Rj=8���U���<���:��<|��[I4=Ը=��<(��<S�T�U�8�U�F�	=y�]��n<n'��X��S=�&=VL�"!��Q���Z=�xȼi;S=��!����~�<}
#=�_�=���<[���4D=そ��ܼP�f=�<�5c<l�=�=�-=#[;�#=���Lq<?8=M_<<���=�*�<X��<��B���I=�8���Լ8�;^b�
q�8%=�<�I�b���L��V�<kp���A��$=��!�{J<1S��G�~e3�0�$��j���ŻнH�Sl�����=a����;��b�;H�<�	�投<^ud�3�*=F�Q����<��E=�q��e3=�Ec�3y)=a�����P��!ټ��I�d�K<��p��Bx;��W<����O��6�μ�� =�UV;g}$=`�=a��o<�}!=(�<Xc��0=6�ȼv�-�����＂�?=�7.=c�R=�
�
�<Lگ<2�7=�i=Zϼ��黱}�Sー�����<�:F=M�{<���<�+=�c1�L(=�^ݻ�o==��n�	�&�2����<����5%��o=��l����f��;S�=iB=��=��8�zB��KC=_u)�a�]�M�g<�g\�J�<dp"=��t=�S��{��-�J;��=��;�.e�:�E="�1=�OT<��K=J
���:=�n=���<O:�y%f�K�o=��=6�<�n�<���<G1=��;��mv�K��<qN=z�=��#�������S=~ԗ��(o����!H_����<����	.�<D��Y*�6�b=~z��<r��fg ���==��<������<���#=�I��Ӏ��p��*=�=�T��Yj��nT����<\;����<3�}�C�<�bA�� �;��1�P��<�����M�V��/�X��ꩼ��p�&L@��U@<�c�<��v�t=W��y��<ƤB=T!S�"�>=e��L�<�f�H�Q�$�<��<\%=��̼=���� <��1<��&<3T<�`=��;5i@�M�f�Q�M<�؇=s=U&d=�c=��/=і���������1�=���)�h��Nj���<��<&��J�<c��<8�(;��<����o<;�I6��`���R
=ֶB��
�<�м���e��=[r<m���J�<_d�<��<I��<��M�׌H=��޼�׼��f=R��6��Y��3�-�4}���o�<�,�:�@=��	=�6=��z<�:�q��;挘<���3=��8䂼�n����Ѽ�a��F�;��==_D���E��h�<^`ڻ�O�<f�/=��d�#�Ƕ�;ED�[��<�@�<ӛ����N=��+<#��Y���c�&=w�=��<�n����=�x���-=��;m�'��s=;�ڼ�pg=�S-�t11��A|<^#ֻ��/�^ZH��%̼jC�<��>��w���Z����/}<��)=���$T��ݍ<�u�<���=�6=�'���7�����=��]=B �:��Y�tZ�:��<����U=̖1�L�<�~����=������m���<7@s=��e<AѼ��9=�ǥ���j�e����=S�-��s�,�*��;�3`=��<��4=uػ<n�Y���(��=��U=j��<�6=%�J;��=n�;�b��vּ�LƻA7=�x=��<u����M���3��,J=��C�,}A�_�h��Q= �/�h�=��,��)r�X�O= &�=)@��1=��=�$N=�	��6��<�I�4?]�?�A<�L$=L^c�]�,<��J=��]��8=�V�ĕN��A���J<Kb������ �Æ�~=7�n���=�Y����&=I@�<*\�G��)�;w�=��ûo	A���<��"<lJY=cg�XYԼʦ�ǀ�<��"=��+��0��I�<��<�$���p��I�<6��<����_����#��P;?�S�[��;m��<!�J=��,=����$A��,估-�=�=���-�7n=W�<0�9�V���t��Wm���t�c�=�8p=�e$=G7;2�	=���:q<�3X=�a��!L?=�i�;\�#�:ח=��A�����-[-=��<N�Y= ݪ:�޼bڔ<�Kۼ�e=���#=��<��1<�I��:='���?W���<�`o;s�)�k*w���t���ў��'I�E���=�-��
���藼	5A=�i����<�!��"N��P�:h��<���ٖ����F������˼O0��-GL�it��2>=Fn�-�<9�!�I��;����7=���-�=�
9��"@=B
��}"=)�;����,�`=�1��˻��=����,ϻ��'�O�)<��ʼ<}D=����l�JU���԰��i�Gia=v�N=�%�L�<�vO=��q�n����b<����w튼5)
=L�<��L��r"=T;��6=�с�'�=��$<�t�A=��=� �<t/=&bi=�1@���k�WZ���6�\�<�7D<�iu���&=�!�;3������v=�xɼ��p�H�N�SN<fu�<x�F=U<Y��jH"�<��:�O�i�<X�7=�m�<�m���]@��o�[���!�O=i��uА=@5>=2V��+�2;tg8�����~$=��<fB�)�<��?=��P��=�-�kRԼ��^�%u<��=��#����.�<č�<(/�>8��j(=���tw��?�<���G�h�_=(H
=����ǻoX��I=zp=����n��?Sϻ��;�㠼E��<҅)�(E���::�����4��%�;��<���?�M=Y�ǻ�Ǯ<�DL��~������I0��U=}�>='�e<�U��(�<�ؼ�|�;Zߩ��H;<��;󞞼�c�Ý�=*�*=�t��L� ��м�FF�;	'�y��-8[=����X=)u<:?�=%?3=�{�<�#�<��<�Kּ;�{��E���-Լ3휼LP{=����dj�׿_�hB��}pF��L2=��B�@[=�$o=3��<_Ϥ�u缧;=�.��>6��z��D\�d,s=�)/<g��;d����1<�᷼���<�am�9%<B�_=�D.=ҷ�<�)��g��lҼG<�<!�4=�s�<�1=W��E�A�J����<��#= �ɼ�q3=��=>�߻��U=ĭ��}�V7�<���<�U�b��<Td<6N�;x?<��;��0<3B=/&μb�
�B=��5��퟼��<`h�������<��0�HB�<�?=�E=�4���0���<�ߵ;OUW����/�<����v���]�6+m����;~[=�����D=�9�<mS$�:�=7`B;;i<}�0=��F�t�s�Yߧ<��M=@�=�X�;%�a(��(ܼ2?��;��<��=�<�A�,�%��<ס>�ӀF�?��]�@��+=b�F��HC��w#����:���<��ټ8�S��l����Y���`� �'�B=��	=f�=����v�5<��
<����:C;�.���M4��n�+7<�t����q~=�9�=�K7���ü�!=c�3=��@���k�kcͻ��d������{;}+R���<|�`=�2A<i��KMN��M�=O�<o���X�;�<gp���C=YG�=a|ļ�uż�=�O^<=3��<�y�<I�����Y<O�&=��<�%�Nu�n����<�`=!��<8}C��h"=x�+�Q�m��;bsٻ�}S�r���<�k�z1�X�<�=�ҧ�<�9=��=$���|�)�K�4=wOl<�tY=f@,�Ez#�PC��a�<�}�<�D"�Y�=/6�7��<`]F<L�0=>Y�<>�>=41~=5�;k��m-���o�m!:b�J�V��"(=�>��Qͼ"|�<��7=���{�<)F	70r���|<ȃ�ÛҼ����E8��=��f�ɼV��5`S��R�4
�<�QM�����Z�����b��<$��2�E�v����tdf;@f#;h	��-�[>��[�R+��7�<���}�	/��n+�:����!��ۭ����<S�S���k7=,���`��Y��!<��/��>=bz4���]����<�<��`=�݉<�g6����;5��(M�<���<D��;�낼<��;!�/=�k���gW��17�֕w����U��$� ;�x��;�;��0�9=����uu=�{i=�T�,NO<3s:K�/=^S��i�\��ώk��f=w��<���<�u�/��&��<��O��:V<hX���o�:�;�z =�Lt<�G=.B=�?�<�'�BL�<ɔS���u��]�5��.�C=��|�������<�ƌ���c<����<�XT:�(�f5����3.�˔�;努���<�CJ�no�<�+�L��Bżs�;�N"=��i=cET����<��8�������>�b_M�p$�=���cG=+�����=CN���T漹lC=|A=U>ܼ܈+;�p�<Qj���»����&���<�� �ˆA=��+=H�������.M=��ռ�$R<��^<��h��[��׽�<�E��@=�ܡ;����=�#��<��<��<E���;U�;��9�`f_=V�=i=$�N;c<�ș;��x��V�<�\k�T=U���w�=�Y�i�,���A��v!=W9=��<b��<Dz�<��<=i�X:y=F���,t�g
����;�h�M\W=b^�<�%�;���i���p�< ��Al���a�<�I�;Mw��tْ;��i=P5{�ӗY=�#뼲麼+%���R�2�M=�䃼V,<��a;iּ���<����-��(S=OE;�uS=�4�;�Ud�Q6�8�I� �C=��U���<�6�;A�.��C;�=�0;?&�*����t���l��< �L<�m�<���<ݣ<����@=��<@��gֽ��D=��=A�<)#��S==�lݻƓ::]D=�G=��	�(����<=��V಼O�X�2򳼓�<Kx=�v%���;p�6<�O:93l1=�Y<hc���!=��8=l�R=3d	=�u�	����F��-k]������������ȼʢt�1�oN�i�ȼ�=`4��	=�@z<s
<��6��x���?�z^<�^
=��=���O;�-����a��Q�=�-�x���H=":��bc��R%����<�D=*�3=��=�U����h���ȻO���:@�#��Z'<1�,��\r���E�Ш;O�<=�65�&n=��i�ĪZ��|�)C =Q���:�T=Ӣ>='4(�[��<�g��2b�x��=?�廷Ry:�.�=O�}e_�Cp'=2�K��Gw�]]��e,V�q�(=�����h\����sQY�P���88=hW˼�p <a��P�ź�X��s���{�d���JǼ��Z�F��8�<'�^��[=��<Ȉ>=���9h�<s�o<��.="�G=�	=����%t=/'<�R�<r?^��0,����;6�Ѽ��*�R��:�ƅ<���;=K6��1=&�%<��4�z=�Ȭ8=��;��<�2���Z=Ͱ=��=>�-��.���<s�l;M������*��i�F=��^=t�%��EQ�H�C<J<x��<a�]<���ƒZ=̿:�!��<��c=�(=M�=_�=c�<*���	�;=\��<�"=nl���b���曻��<G�<(&	��Ǽ<�r�%�g��9���U����[=,(
���.=��q��V�s����z��z�<�R�<��<=�'=h3�<(��/L�;k�-����;��=�����X�zb�;�W=U�0=`��<6��<��m������ds��=9'
=Y����ZD� :�<�N����g=�R�B�żP�1�ɇ�ut	;�A��c��AƮ��J��A���Y=9;���)q���м�^�<T�l;^��<��;��=���Z]���=j`=Íd=������8?��6����J;=.�!�����-��%�ɼ�Q�uZL<laּN����D�9�}��5=���<E��rY=��<��=�W'��#���J��� =��n=�I~�����T
�<��G=E�<�`�;�c=ʩ<22D�j�*<p��<���<�{&���'��/�ك���<�,p;k�D��\==�/<ڀe��0<�[����&� �+�R`�I�ͼѰX�|
���Ǫ��5[=b-y<~�&��+9�W=��=e��<�5�<<=�#5<�#�<��.�~μ��k�_B�:R�(=|�<T� <�MԼ�i*=�1����:���r%���4����;-����Ƽ�qB��7�-p"�Ea켉|=�sX���{����'J���o��z��p�;k9�|���m;qA<��!F,=�����m�<�����M=!p��Wɼ	HݻřT�WM�<�ǂ�r�:=~�W�]|�<���;���xY�k,���!�<x��<� ��|���6<�o�<��;��<�ҧ��<:q�<Q+��N� Yq=�<�
���W{����<�~����Dݼs�r��7���1J=	�.=7\��m����J��=@f ;����d=x�N<��W<KA0�sM�;���`�#�aN$=&EZ=J4D;�5�<��<<��<������<�F��8B=x�G���<?�3=$�0=b�;��=g�x:�7�����ʜ-����=#P�<�G�=�no=9���V<V�K�8��<a¼{į�f�L=~hA;������M/6=�J޼K^X<�lt=�ܽ<_�[��m�����y�m=���<�7�=��<��=��M=_�b=�==��<���ڬF=�Nļ�93=��T�>�=�������Ѽ�fr<]W7�c�.=CT��n=��;���C=X?��J�[h\=��ͼp�=m�H=s�3�DDu�����<�u=��J<��z=+��/�=�-W��~���{�`�0=��M�J�=��=����S���%=�%мO�c�"SK=E%r�9�<:�}=�Zb.� �.=�R�+��<��n�h=�n!;؁�<� X=��"���g=NF= ��l��<1�ֻ�
<v\�dӟ����ft��amW�獽�i�<<i|��WN<ɖ�<pV<�PG<+�<�dn�'��<D�Q��^�M<#�a=%c����;=F���B<�{=xv:�X&���Y�R4�<�?���<)�Y��2��k=�C�=Il�:��<�f�&���#伦|Ǽ5�]�/{�tC��GYg<r�@��Vb0�15v=�+���#=�P=�xμCE=�jw<i�#�4��^<M'���;s�ļY�'��ü:�(����<3k=��<q0���?F=�e��D�;"�-���=w��+X��g\=ٕ��-Z�$~F=x��<�r=7�Z;	�����������{j���A=��鼇���F]=����4f=U�"��H;Wz!=6�n;�6=VF����<���;�̨�����s�J=n[K;��<�k����~Ӽ�8�<�is=�<�(�мF�~��<"͙��0��$�������̼<�?=�d�]�<F�!��7�}���X�)��=5����C*=�؍���+��[ּ�,x��?Ӽ�@��&W=���H18������<�J-=���bi��W� ��(p�L�<�R;W/<���<��R=p��,�^</ׁ��
D=�� �ܥ���k	��-l<Jg�O^�DF=��<C�r�b��<����LY<��C=f۴=w����>=��������吱�?�/<,����]=H=;��c=z���p����<G�;��i��CJ<1����za�F�� _�<�L=/|;W�;�O=�J
�lq�<)�� Ȟ<��?<5��<Hl[=�}"��9��7�
�=E�<TYh��t���lS<Y O����6�C;�=�d�;Dܘ��C�6�<=��e��S=ΌO�w>��;�SC=$Ǽ��J�}�Q<�=3'\='l7��+�;H}���2'�$9�<���H=�>��T�d�r�Ւ;=T�D=���wA��3;$k�<�u=��M=��üT��<�qR�<<�EU�6�<׈��_�<蹫�>2�<y��s�i��?=>�Ma���W��IK�Jܸ<"	<_���~��8Y�<��e<挌<k�+�nm$=��;���<dR�=�H���Z�<��h<�=,�`���W�t�$=���t8ۤǼ��e=)�S�
��0E<��E��C�^�=�u/f��8�<�����<Y�;���<�	��! =E:/����y�"=��d<Z�{��Z�gB=�����p=Fh��*J	�0�)=ɞ��<IH;c"�< ����2���\?���V<���<�N= � =���;{;��S;qIY=�-!�d��;C���f��"��Zg<�2N<��=̩�;�g��O�#=`G��jƼ����~��˓��xx;�[=��μ|ٷ;���<6FV=�*=hb=�;����<X�t=8��<L1=%`\=_�ټe=��<�������<杭���0=B�X="3�<Pa���߼({G��[7=d��@��<�O��f�=@���<=��;y�X��HP=�-\�Q��;h�W���>��7Q������|=7V�=� 7��Ga=�H�<�Qx�:�
=�s�<��^�aP���K=6��:�/��F�<�L��=���<� \�ȕ.��ź���[��5�μm �;���<�!=U�<w�J:��:�_I=�t���<�C�<���<�gy<Y4;�)=1Dg�b�2�^=�6��p�ҧC���I�����gT=[E;��=���<��<��X=���;n}#�����G��D�;�u�%���4�ֻZh��5�Q:=�9����T�Y<D�@��Q6=΀:=���'S��K==�7�<o>��� ��>k���Z�rj=a<�&#;�KB�\8�;�t�<��m:�:4�m;��r���;�`	=ǔ<��8��D��T#=1���1�<��H<'�Լ#M*����~==�_�:H*�-�?�5�4=�)y=L��<�"V=P=<t�<�[?�azJ=)��=5����T�	�ݻ�6-=�����a)=A��<a�=hr= �/��&=�}=��F�����Z��<O�+=���*=���xr��b_��D�;��,��=n���=�5m�`>ɼɰ<IWݼ�_ּ,A=`QM�2D���B��2H��)�D�5=:�<oO�:��������W=�6O���T�)�:=�];�R����q'<�<��=ywN=�@=�����3=�.<���<���;��%���&�2�M=�0���h�����S=�l5������C���M<c��<-�<t���(=�ռ�n<<u�	=!J=V\�<��U<0�ܻ��HN"<��D=���y�W} =r�U��e��g�W=��D����o_ۼ�<0���h��$�==nYG=��n<���<��;�ԼcO�o��;;M��A�<D6�<�&<+�����$�*'�L�)���:��'�"�Z=:!=M����Z<�DD�}��<��;,�f��`����乼<�L�KZ<?���+��aQ���x<���<��	�ݓ!=8�n�3��<��;tdf=ْ#=�O=s�u=&"^���<�hJ���N=��5@���tr�� =�b=�yC��FX=���;�^��3����;��=��]�<_����?3�)B�?[<dTF�,p<=�<�ɯ��3��g����˻Ɇ�LI=�dI��T4<�<k<���<�4;=���<P=%�<ܿ���S�BL;#	��;����I���n��㼲f&=�T�&�=��,�h	(=�|X=/=9��<Ш[=��?�h���J�x)P�
�j�e�@8Q=�V�#r:��<�Y4� �t�1[=b6=�xw=\�a=MM��e�<���f'�
�c����7�>������-����<�$�<7�f='j0�ڿ2=���Dd��>����=۞j�5=0�`<�=ǟ0���Z<���<	�꼆kq��:��)
�=��?�,����ټȾ�.cR��D��I��<�z=����a!���k�;l� =���<;�)=�S��u�e=�X��2=�Ἴf=&�<�!=�<<[�<惍<_T�;ծ#�S։�
�H�ӄ<��Z;-�:��,:�}��lk;=]_=f�:^?�|�=�M=\;�Z�E�1��8�ѻ� =+�
=���+R=�������J<sQ���=���5��,:�IT;���9�y0<��=��	=��<C�с<\u�<k�/���<�r���0�I' ��E ��<�:�<�[��}~��h�s�x=D��<�[�<g�;�n&G;�<Yf��"=1x��m���P=lü</=�O�<K����=ʇR��$=��=j���T�=i�`</�A�mО��}�;��<��5�,�U���8���T=���%N�nKD�؝N��Ks��X���	�*��<^�Q=�=�g�<�NW=Uj�<Z�=NI=��=���ǼT=�<�e����9<m6<d���¹����Ҟ<��M���=(<�)�;"�<ָ!;��:''�X��<��S=�_�<(y�c�/=���<zЯ<ɣb=���<M�L�,�<O=�C"=�`�ח�<?$l�C�i=����갼�j=��;(�p�݅K=o�?=�G=����i���@�\�t��>�����S���;=�I�;�(�<�hB<��=c���<�:��s=u�ؼ�(A�2l�<v
-=)���Hi>�5bW=@J��a�;,��ߔ��j=ɪc=ҟ�8(���=;.�:�ꚾ<Y9�<�W==ԐD�;®����8�=�u$+=� ���q�<�lb=m5=`�������:$����Y��&���;c�;�����<�)�N�F�%�0=��<�V =���������L�T���1�<��
��N����%=�'л��-�f�y=*��r��<�"��[�?������`��͚;���eVE�I?9��q=�R=HF]=cA�6:Y;����ɼǅ1=�!�=Y�`=�=�^<<?=kw�4�a�� K?<a?l���$�c6���|=�G2=��<?��<m�$�����<����~�x��J�<���;������O��;5��f�<L|<���<'6��U�p}Y���O=e_f�)=��=��=��r=�<O� �_|I=�
=w͵�ѩ����pۼ��9���8�S��<w��<|ی:S�'=-y�`�8<�^=�\a=�8��S����j�7d->=Q�&=�<��j�y"ûP
=e�<K�Ƽ��4��蟻]������<W+�	��m%�<�'=�N�<H�=!m��;�<��p�2	=h2���<n6=ƙ>=�𪻒79<c��<!ZW�7W�<ON0<�b��=�;^qq��`�<-�f=SA����;���<�kd=���<ۓS=��Z=�%�<yDX��Ao���4<4x?� ���u�t=SW�::�A�T����y��U��P=��H�:��l]����,߻�=�p'="�����>��D:=��<(��l#�<>U�<��=�[����T:�~%<��S������i�Î���6=V�U=uڼ	m�<�[6��8i�f��U��;�Ґ<,��=1��;E���;a�2�<��=B�h��@��rB��̞<��E=#�R�c�!=��K�\=�ӆ8����;�;u�)WF�<|�N%��dA=o�;`5=�Y��k��6{=�̼����b��	U=ە�;�I6=IEr=qf�ls=T���>+���b,=�;V=4�C�5�Wz��<<B�-<a*L=�k�<�*�@���o�G=��������"n;�����(����l�&�<[s=���
���<��T=��B�Gʺ<��^=U4@�̍=g͔<0uo<u��	:��=Q�=�T=�Z=2�#�D��;P*f=�(���48�il=�/�<4�	�o"]=y$�<ȵ"�割;g�1<����N���ɼD�=0-��Ͷ�OH<�s�;1y�;�<,l뻂c�� =����Z���c����=�#����}=6a*��C=frC�m���0=�4S=L�%=3z)=vi���as<џ��TV=��=XH�<��g�~E��r���t=V�W�"�ļ��r=��<� �;��.�J�7=@��<{5\��~���8<��<��2�&G�<.�%=��u�W�,�J@N<�!�<0P�<��=����g+=)����<ڜ<p�L�^�q=��.=y���y����;�񲻎M˼IWC=����%�;4=�� �_�8=h^�_ܻ�S;=�Y�\�;�.=I�=�<h=��j=  :=I�d=#� <�,�<��ļ�nd:��<"<=�p�<�	�=�"�/���(�L�͠�؛A��A��p}�_<#;��[�y�
=���	>i=G�=\I�W\e=ȁ�<�)���4��e.;�����8=�;>e=���<���<{_��;F=!v����<�t�����g��q=���K�RJ�;�!�<� (=��;�Էa���<k;м�}*�֫w;e����ǻ��<���%fN��=!������n��NV=�$�<��C=	G�7�&�^Xa��(���䳼�=�����{����M��*F��G�<��J<�f�<�<~��p	�<�ۺ,�R��9@�}����yR�5�7�Ţ;�L=������+�v��<~�^�_c=�Vt��� =�$W�W�}=�=w�F=we��<�X�=HX�LXK��/=-�0=�������o�d�'P�<���<����L�ϻ#�����q=(=�<�D=�"<��V��[F=����6�<5.�K9 =��Jz7=��<A�5��@T�{9I=p�|���޼��;T����<f��=�S}<�?м���<|�<�Y���ɼ�mT�->U=$A=��0������}�@��N�w(}��A����:$�s<��]�^�	���|<F� pQ=�j�<pp_<����м��}�9��c.�;oS<;�S=yҫ��H�����IQ<� >�2	�����>���x���=5y�;+=�|��:�8C<�o]�[ߠ�M��<��=��<8��$���Q <9�9�-7=z�I(=p������z�<���<Ƚ?���H=�Ȼ���<���L=�?l�Te	��|5;���(P=H5<%q�<7���x�=���� l=UG��'�o=φڼ3�ļ�s =�(l=�2=-�M8꼡�4=��u�.=�¢��ck���g<���<�e��	^<Е��a�4=z|���껺ײ<ZL��=d��=O-R=���?M2=Վl<��=,��<��P<����*��@G=3�/=�n4=;�o=T����W<1�o�/�=@<�:.C�;�]e���=ꄧ�-޼��?=C��}�ü��a��5 =��I: <�����z=��<V�=���<~�ż�ot<*�R�'��9
P<=hK�;ﱼRiv�8��E��;�2�(B=�9<�����ü�[�a���P�%:�ǻ�7O�Q�ܼ_"y=Q�	���%�7�=X"=wDD�3��/��<&�M�<u=\ =^����,��>(=e=,C}<�$���I;�2�#�Ӽh0�� =9N���{�3㱻S=�<��=B�o=cA{�f=R�{������s-<`<�K�<��Y=����<b�=j#��C�ܺ��==���<��;lb!<�NȻ/���i�_󻁏n���u��z!�cV,=�=��)=��I����=H�p=��p=k<*��<9~Y���-;��h�f�;��<Zg�<;�b�ܰr=pJ�s�2�G�<��f<�][��^�<X�E�	;�<V��f��m�=H�[�O'�<0fv��-�Xx	���=�oL�I`B�,����$<Ǘt�6�:�P��<���R=��i�3.;`����B:=��=9;���c���p���i=�#�:��k�i<�#�c=ݭ�=�F�M�2;�<=���=�QK==OL=�(=�)K=Ë=�N��[���4a>=~�Z=Pb�;�H���Ԋ��Mx;!u"�_� �//�`�;��H�@J�2�����<sͿ��ꈼ��0��4=(7��&
��Z�<Ԟ�<C���ڤ<:��;:=6�!=2�E=I�T=4�j�m��<N�q=��!�����8y)=Qk�v�0����<�S= �<�W�<��X��!9�9:�r� =ɑ"=�9C=i���➼ �ԼF����L��:n<6����";�@��'�;7�D<Y���h�lc?=��漚Jh�E*=���)������<�Nw=�V'���2=�/����������;g��<|�K=zH�;t���V<=26��݃�<��<�Q��h�<��	=1�o<s�+=����O5=UJ�<"�=����5��-f��z����<)�=\n!=�yD=N	�;9Aѻ�W�<Vh;=��3=V1�� �<Ā����[��y���Y��Q?=:"`������'�D�q�6�'=К=��<�d=�=��m=�s�H8���7K=���<19=����6�<��^=�1]<Z��<^ļN�;=�9��e=(�
�2r����P=v�,�r<d�J�:�wB<@=�J)�$���~�<Jq�<�T�֋�;�J"�,J�E%I�� v�e|�<��@=�;ټ?/t;��<5��<Hʼ�6�	��<��&<3�C�����-���uc���=_�<���s$�U���p�;#������0 =ɶ�E�f=+�!�veQ�=��L��^��%<V�<����������z?��%_�Ċ[���W���<=I�O�d��\�&=n�2�at6<������<�=Z�;oWT=iT:����/=��(���"=��N=�M�9%�;�ՠ;<�K�E���_:]z�����v6���bc<�g�G�=;,C=H[=<TJ=��+�$$<;�\���z<m �<�B��`�=�*3=ݏ�;n߼L!N=1d=)����m'����<�V���4�<�l��xj<�9�:Mv=@-�;�&=x�o�?��� =�~�:�<#��<�C��Tz�ס=ڙ����=�:��n�<�ڼn�� ��<���<䵭<Ҫ���L-=#D�� =�8<�[�W�� ����Bh���k�C���U��V�;,�e��	O<�\<I�/��z=T��<$�&=�ř��< ���ͼʃ�-�B;q���V^]=G�����; �=�=��=n�*<Q��<�H��Jq�<թ<������<�#=ﵐ<m<�)�;�<�g@P��u� �O��Oj�?�-= 	T=�n+��x���H�<τּ#�=���<2���R�L�4-�=�g����<�J�[C�<�i����<T���=��<�2ݼ��S;I~2�H�=����o�j�~f���=5��s/<=n�O�X�)+��'�=9E��{l��R�kt��[3k�e|���!=��(��.<�"=���-Ы����<���x��H������r=��!��_h����8 =�9.=%�'=�r�<d�<�z�q��:�a��BB==�<=����i�f�J�1�;m�;�c6=�0=p���$���q�<G`<Y�`=�k�<��ܼڙB<H�=�=+�V=s*��To��pI<�PE�H�C��#����Q=e�P��n�;�C=�-��3'�L8=8��<|qE�&��<�Cl<����.;w�L�ZZs=��j='쁼�L7=��<΄Q�"��<�LP��"]��9R�B��N�E=�oӼ��*:4Ἣ��<4��6a�\�b���&�;�=�v�;c;�<��<��+�D}==�l;�#�A���b=��!=��<��T��(�<"&	=K��;	�<���<,#�<�@�;�s������r�w=��=����Oku���y=�iɼ�F�<p�=ӆX��|�8�bh;]�D=�<ӻ9���^�;j�gDX���9<"�o<�T�����`���8=��=-s�GL���uX��Ԗ��G�=d��k�;~kU������?<�$�I�9�Z*�JM��^
��c<��+�W~l;Lnp<��R:��u�I�>Dh<d��<��G=T�< ��;�x>���=M��������'�;��ݤ�<o*��;��O�;�D�Y�q=[޵��+��Ѻ��ޒ��!U��*�<o@=\<��Z=k�T�ӕ伐�ټځ��֞��$1_�N.�<��d�J�S
�#_��;��u�
=B^(=����p0����<�>e�]'����g=v�E=dw%�2�S�F{�9��;�Z?��)��k ���x�d\ϼze�6W��<%<�+��M=n]o���=�}�h�"T���ݷ�R�����#��G��=y�=b!�;2E'=�4��B9]�>�{b=s/#<:�s==�����{<.��l�	<�Î<������K*<{㻻���@�����s���=�� <�
�;�k�;��d	���G=y=��Ԝ�z(���Mt<�Ȍ<�����y� f==S7�N�o=��<�=��;�I���^�n�\=��(=�*�<Ӵ� ��;�;T���=��<>9=�}a<�$g<����=�`�"�q�7K=�|<g<���N=��/�� X=��<��A��+=!�<��h曼1k��o�;�P�<����/Xb=�ڷ<Ac=Z��<C���g�I<�'A=�� �v����"�<=9�<��2�D:��7�
<��=Sp��+/��T��Ԕ=�2=��=��4�0��Ϯ��È!=�P��dS����=Kr�<ݜ|=��<�iͼ:��<���=45�<��滾��<,�=��o;�ܡ�u�S��=� [�<�<z=6<��:��<���<-冼��S=�į<T�<�6=z��<x��<�k<~�=�K�Z3-<�
)<�K��o����<�ZX<'�T=��<�d=L=9�=��F�Z���p�<y�g=u����O�!�4=�V��Pg�����)��� ���>ǻ>���=@�X<?l��>K=4���U��p��Y$=t�<0м�Í<p����Y��QP/�ZeN=�9�9_�\�7�h���e���<�˫<_���=U�4�r�ϼ��3=�-h�酉�X�<��;��={G=c�;�=��<��.�<(�������̓<2��;齳<�z��FM=7i��uX�<E�����F=�����=� ؼNm�<�>l=A�k=�@�<�^K<>�<.�>��,F=�y.=Eü�fS��֦:; �����~��IN.=�Xr��� =�LҼ�We=��˻1a��5Y�=N�iP��)���|F���V���[<��4�_Z�Z¼�<˼��]=_�N;8���a����2�(��;+�C=%4+���#�L)�<C�4<�=(6<?u�<pH^=CmO��"=$BA=Q]�<�Y�<&��<�Lk�	�a��Ҁ<�;=+�=� =�'i���Y<�J�<�ߍ<��}<I�<�H����+=iU�;��;���<�2=��<�iR���c�+=�=��f�����VA�n�q<�[�<-<�<�ӄ��b��M9=y�����<Gj=$T� �<=A����΍��m��;=�p�,kz��g���A<B�f�'���L�z�Y��n(<�=W�
=��U���*=>?Z��+��b?ͻ�D><�f��A5X�G�w<���<0Ja��P=�)D�t�=P;�<,=����<��R���m=�h�<]l߼CvM=��^���<��<{d"=���<.t=������ �5=Pf�<;�P=X�;u�;�\�=��^�KI=�Z8<���:ZE�<�v�{N���ϼo�<T����J<�<G�d=�H�<Ѱ4���O=E�'�}��<+�%=X�.=H���m=��<8� ���=k@;��-��7�<	�2���:�l=���;f���BH=��ؼ����ާ=��J�c1�����;Z���8�_��9q��^=�<	~��4}:�{=�F�3�='P=���;]�U�v�T���J�	��$�=������=���;�?8��)c=�.�71	=`�c�;6��?<!<\R=@�c=
>��	��Ρ ��T:�Čn=��Ѽ0�H���^� j����P=N�<�{���z�<�;Pg;W��`�4�ކi<~�}<,#e��%�Sq����	=���R=ȪϻU��<��R��=�>;"-=���9Uu�.$ �|�=/�@=����+<f��<�%��uh����<~!�<q6������_�l?��M =�[r���<�g�z:%a�ꔍ=��W��}$��K=��:�RC�K]Ǽ��޼X��<�1����< V<�{,�i�$=J�:=>�_<�鄺nY��Bo�-��	�G=C>	�|�[<��(K<4/<߲<\Y��8g=�(�<��B=n�<'`.���38=-�>=�oG=]��)���'��<�N����������y��5�K�[<�TE=�5��1;A��6��<�te��&=N�F�4�c�W�=W�F��發dC=�u�=�fq=�s=��Z�<���>68�,߼�J�;W�����<'[A�N�b:>;S=8X#��vh�b2�<��<������==f�><wQ	<��CH�<�N��n=9�=����O�<�R�;�B'=���<��0������c=��6��45<� ����;3��<"��Y�༰%)���鷛Zm�㨹+�����}<?$��o�<'VX<��)n ��j=/Ő<Y0Q����b�W�,[e<��=�=���:;�`;Ȕ=wl�<�N=��=�3~<��:�4V=�%��Z=�2=�A�<u�=�����Z�<xN�	<�;�Q#��D=���L\=-���S<A���g6��q^��Pc=�8�=��Mü5$=<3�<�UѼ_鼊��=�7=\d���_�z�="6'=6X���=���+=�u����:�E{=�i=!Y�<�������D=c5�<�<��tk�����l=���P�<�a�=�I.=?�q<x\�<�"���Ǽ����*m=�żH=��=����ҼsG<�8=욹��F=+�^��I?���ŻC=�dO=�W;B�A<OV:=�r�9�=׆J����x�g;l����g��@9�<1w�<�PD<#�.���a=�T�͘�<N�;;r�;�z�˻�<�wO�}�<���;�a�<��s�-�ۼ�`����;z�<��j=ɯ�<1��5=0仼\�<��%����A==���<a�=Cp=�=�#0=�~=�=Ҙ<p<�@��e=4�K=�>t<$������v[<��|=IWi<h�<���Y<ռ�#���`L=}k%<�#�Z
���3C<��e�o����s<�E�<�c���MӼ�^��<�ǵ�U���@=ptN=��_��#I��矼���<b?s<�+�����-�F4��UP=*}�<x[���a����@�[Z�<�	�+�����<��=}�o=�Š���/<�2�	>=�:��S��=�=OG����L�=(�	=N��g���<.��7Q��<>GʼP���#=�D��(���z;)���h�Q�C�=;>]�ܝ=��=����W��B �5��<x�W��1<�"μ���;n���6��4na�B�<¬Z��r==��<�=��Լp�~��G<=�0<5���AR[����|kc=�;O��/��ٔA��t��8� ��<��N=J��<����W�*��yV��+=j��=Z���*G7�sc�=ơ�%��<n�<c氼	�<�X-=�<o_<<���$�����<o��;Z�5�G�����X=2b=*��\$�S��;��2�=+<���<���kj�<�=�#= (�<��缩�����g��p<EoB�-=�1�a=qR�< �tm����w<��s��r���OM<[0���Ѽ�%:�@�ۡ�<9�<W�Y��P��__=��'=;3<��w�L�X���޺$�F�SD��ך���<
FW=ʒ�<���i�<.M�<[P�<9!=#m�h�$=�"=�[=�cI�_���t =���=��z�K�B�� =)7A=��=����=O�~�;�w����#��n:��)�UmX<y��r��<=��<ȵ =6"k=����:�c���<
���iS=)�=�?-�I�F;Y<(=�T=�D=���">���=v�U�F׈�Ćd��:��f����'�RXW=JN��%v.=6�����F=����/��<�:=�1�=!���p��:�<�O���<h������<�v�6!-<�)c<��=�e<��<�v�<"�<M_4���V=��)���ȼx�V=�6�a�*��6�<�H.=���<'EC�i�;	��<�ҏ<q��< �l�N#/<=/<��꼷"h��_�:��<�H=K7�<
2��X�c=�kd���@9��<'$|��|=��[��O<���<���<�FP���=�2<Y;<�f=���<io�۶`=eۂ<61��^<��7=���1���j��{-=�=2��8��Y8��
���FZ��==C���XN%=��C=G��oR=E�����&=S�]=�4��>G�<"�(���3���]����<���<p^|�M���$E��&�@{��d}���<��x�aa&���P<vr,�s��ɑ#=�Q^={��=�G=��_����lr��ۓ���88��;9)���<�Ҩ<��T�{�<��2=��<f�1<i��,�v����<1=g�S�� ]G=b��<�����8�<�����:���;���<��/="wY����A�C<m�[<%"���i���C��/�<�=�qB={��<�oܼ �ؼꇦ��i`<��e;P=�������ρ=q�d���1�-O����<㒼Q��V�<*?r=���<�!���n=�mh=!�N<�e ;��b=���f��<�H?�m}f<�ۻa�L���=�.9=K�����;f"�<���<���<�#x�����S
<�ZU�	�z���<�Z<��]<�l�������a=�x��L�?Q?<F��<�$ǻ�R���P�@l��PU<
AG�Gry�f�1;ͺ���ż��P=��<���;x
O=����	��C?��UK�/A=���|:����U��y=~'�<�:=�5=3�<�R/<~g��g�U�=�����={uм;��x�O=����3>�<�y`��n�<�d�G�<D���T9%���&/�\���<����Zr;-e�;��<2��\��<�1�<8=�+=�~^��.=�� E�X�>�M/���x��f���=��G=�{���Ŧ���;�X�9����|<rO��ݍ#=���:3�x=Fm}=�2��?v:�:=�����;4C���Jv;�吽}-=@R=Ko���?r�{�<�!���=��#=e�:��&�<@����p~=�7�1<N��;��;��C=[�L�/yM�ƴP=���<|��<e��?�����'=��V��*��2=�Ʊ��4=+���`<wO[��R��T;=���"������;_ke=a�n��1�<��<��:�T��;���<��=�üs�L=��L��=oˤ;.�<D��<~3���=��"<��=��<jv��}l=��U�D��	V=9/����<(2T�vmD=WA�<�!�ݕ��@�*3�r�m��ۼ~���|�<���<(A�<I�L�?�ż�i��"�����:�4����)e�<0/���N��v�<|��!ֻ��==tH���̼��N=&1=�B7�LY�<���Ი�c�<��������6l�;�ɏ:)���;�<�<.��M=��8�M�����;�V;=mv�<$��;�c@�"�Q���<C�l<�5_<}��<^9�����=�1M=f[3=}�=�Y&��ė<	���~r<�hR=7�����.��F=��=U���KӼ�r;�Ni��K�<�n<֟B<��.�}-j�P�i=Nu�<	�?�I��s`�`Y.���E��N=�s+<��=�a=W=g�l=V�N<�]���j�S1弪Wc=�X+=��z����<�N�=�1�"L�%�=ſ��⮼�k0��=�$=]�=����N;�Y�<�^���㾼���юF=aр<�^��DU�<�2,�hbq��@w��:B���;��m=��o=rT��$��痮;�<C=���<��m�'Rp;e�ڼ�#=hE�<+^��1jX�7�d;�F
�zJ�;ӥV��BP=�=���4/L���<��+�h�=���<yG =�H�<\�R��d��K׼xMT=�<D=�T����&K=��:V�*�:ζ;�L�<<�$���ջh�<�q�=Ԫ<�k��� =��;�tu<��O�_;��c=�I=��;P�<�l��T�<�-a<�==� #�P� ��ƻ�z�C��K�<�}>=>�=���1�;;E}�G����$"�NjӼ�K#������<��K�U���?=�(�
ϓ<P=<�M��u^�<<�(=� �!tʼ��7��u�;/c=W�M=	�(��K˼�<�!��0�(aǼWC�<��4=fp�=��%��'�<����L��K���[�h?)��|+�r�c��!F���l<`�<���4�V�k��Z�<�
�<��<.N1�%+0���:�ͼcJ�B�<~�;,w =�	�;�n�;r�=>�|��FJ��F ;�e�<�J�1�z%�W m��Sx=te�<"��<i<��W���N����u�#=�~�<��m�>�=;ME<L�g<-@R<;��<�o<0�2��u/=�0=��-=~�:��ۼc�=����	%=� �Ɂ0��wW<J�;=�}�=.�I�ZX=;�����<�l�̏,��Pȼƒ��@(�R"=���<K�,=ч��]4v=�;f=g����\�]����.=�����n��TŻ<�%<s�G=�`;��̏;�(��KZ�<q�=�6=d�F=�}F�=�<�&���4��5=��ޟo<���:�q=�9;�Q�1k����<� m�cK'�v��<m�<C��.��<�ļ�O0=��d�����<y]�;K�<3F��� ���p�WtǼ���<Z��L�c��DI���߻��v��x�
����6�򻹻5=C�%�(�<���<$!�<�_�<�&�@�y��<�6=��=�>�;�p�<���<uڶ�ڃ_��a=����VF�:���;H��<:�Q=����t��<jx=)��2�=^�t��2F�.� <3���iW;(=�BO =J��&�/��ή;���<ޥ�4O�<����q�$�2��eʼ�S<��̼�<�<��;%�������K�������W<��p�kߡ��8=%q��Ύ_=*ȁ�R���zt=�,<���<����Yɷ;�=�ɼS_J=��s���<��c=_�;��9=�%)=|]J�=���x5��ˬ���x��h���7�<[���8h��>�8잼i�<+B&<p���?����=]{�F�I���S<��<��<'r�CnS=�1:=��<y�C��٬��s7=��r=__*��D���/Ҽ��e��?���y=�B�ձ=��P=ƥ����<Tx�<`i���1=��n=���;OB�<e=��*$<ye����=�J=4&&��<�;Y�<߼�"���q�w;8=�%Ѽv7�u�g<�ͼpG='w��*�=pΌ;�hD;r�8��!��R<�<��<�]�:��=6�3<�<=�����W�<����U=vx��N�<褆�'A!�A6̼ׅ�<�\��<K��o.�=�����@����<,C㼗T���OӇ<"޼�=���=����q�)'f=���~)=`;��#~��V=6����;!=�J8;�<ݼ[�S��=������e<x�b��JB�ڼd������<-v=�\���><]9�����<)<s=��<�[���$R<i��<m�
��Y<�
�<��6��aV=7C�<4�E=�T=���;ԳD�;����Z��ѼZ%$�q��ҙ`<�Uk=m��<��Z=��<^�<��;�'���Y=�� =X�R=Uۨ<��<��U�����������X=*��<Ϋ^=je$<��v����<�`%=aT����/= Z��͗�<U�=��5�&�<��~�9~L��.�<�n�sg=�D��|��9�<r�W="�N<�L�<ȅ軂�<^%0�����:��L=~�g�mZB�n���7�0�@���g5�:�<F�"�������<�~=���<W�ҼƖ=��(�7k��O{
���<b�Q���,�wۖ��(=�嘼�jQ����$4�`��;�֫���*���pC<P���*
=��=�?#��1�=�S�z�
����<t�=>d<�'�}�h;�C}9P��. ����=:��E	r=oOr�J��<�=�Ϻ}�=5<����O;�;���Fh<�9�;�S��4$x<%��<�@U�~����@F=�' �� �b'8<y��z[=�-�d��pR=(o7�9輖QY��j�<j%A;�����0�<1���y��<�!�E�0=<n�:_I��r)�����P���J�b�)=ʛN�z�D�sg�<����D<�<a�z���j=2�=d$���:t<��<>�K��,���"�;��r=��<9�=���_bq�	'�<��E=T\��e�=��=�rN���;�2\=�~F��5=�f@=�Wx<�C;%a�W�|= �<I\�fW�<�̺�n���(��<�����:<2�\;sD��{�C���S������3h<6"�<��;.��=��:�+	��T��>T��i�<@���5�8[��~�3���7=J��������;��ۼz#=8u�<�&���_���*=x��;ֺn<����P=x��<??}��Y�<|�*=0�W�Z�༙0}=��<�5��,���
�<��9��P)=&z�<@�<�4='����<�1��'�<��g��6�Q�;wτ<������*�r؁=ER=����8=:q=�0w�W�3<�{%�U~%=��=>�Yc'=T�=xN
���<O�;�sH=`V*=.Y*=-�r=zk��X<���զ�;��*=��0���<'���I�< <��Мj���m�һo���@�j�H=� Y����V�t�Gpb�����BF=���;f"=��k�r#V����*=݂=��^�S���5=�\�<�Gw;���<��՗5�W_;<�+q<��=��2�&}�������9�C�
ho=�i=���<�����Su;�i>�J�+=3	=Bp�=S�1��-=��B�1�V�^��[q}� ��:��ż�xZ�V�S�EI���;5�{��3MZ��-�u�<�$,;�쇽���<��A�Q<��;~��<��O�1���]��8=}Q:<$��7b@=���C�"=7���I��;�=]� �0C.��-	�
�;;�����z=CX<im�;�8\=��; DM=0��;��<	r<���<��d=�R)=��u[=��.;3)J��/�<7�=��\����:��<�3�;tL�<�q�<3�w��š<�v6<cd=V�<=R���VmE���ػ�<`�p��{_�hu<h%�<�}X�be:���;.���d�� �xQF<�	��s�S=�5=�{*�ܤ�<�;� ;;zI;�߂�/�s=�e
=t�Ѽ�J�c,мj��;�<���pA�����Q`��B�<)�y��By=y\<yGB=l��<Y�E�+�!��Ǎ��Q=㭙<��;o9=&S&��)=��=��.����<�<�l���ú�K=��W��&�<II�<�`����J��BütKL�U���,v=��5�M =��n� 7=pg�CQ}=��;A�D=KD��r9�9��C#<�21=ڒ�;��G�>�X����<�$`<@�_��b<U~c�
z��RJ�;�HR=��G_��r�|<���<@�9=n�˼�м<n�m<�<H6=r��R(��x����x���z�d�<Ӵ��e!���D�r)��&���J��w�`�#��@4�6�\=�rE<�w�<�켅U6���5�Pz��$�;8(<�f:�a<G�h3��a?�<�ȼc��\o=���U��O�<o(|=�V:=���Z��<��ĻL�S=Z�<n��Ri=ƫ<�����[=k_g�˞&��_-�M���ш	=��;S�Լ!��`�	=5ϖ<l�=gH�<���< ��<�&�<\)�b���"�Z�+�i�,�~E+��8=w �u5!���;D�d��R軝}m=N����E��j�C�Ҽv�=���<��t;�V=#�=�D�ȘX=��i���׻���<�u@�2���nռ��J=?�;]W=}�=�Ot�T��<|�R=D�$�B�v=W��<O� =X�|<~�7����
<��,���<fvȼ��<qk9�^gO;��<T�+=�D9=5Wż���]N�c�=�Ԙ<h&P=(+��F�-��K=͉y��<ي7�A:�=��;��S
��,k=�=A��:O25��H���<g=�=9�'��*�z���a����=�}��9�=�G��x�<,z= �6=��T�_�<b)�;�e�<�g�;�W�=��o=7B伪h�<;�=��;��n=v���T$��7�~/4���<%��<��<�"'�����UN�����	��<���;3)=�=� =���L�}��<ҎJ=[`=�7�r9�LG���Y�:3]<�ƹ<����e9�O���=[��{�<)�<�(3�И���B�����T(n<�x<P�Y��R�<S��<��=�_�;2��"ݺ�*�<�5�:�Y=��4=m/�����]���y=��a=j�*�m�|<�ZM=�+����;��g;�{�:E�N���@���=�<O���Y[=�Z=�����L�ŦK��l<h(n<뭗���,�<a��mC<^o=�j�<
6/=��A�Ǖ<կ��S鱼�o���Z�&_���=�/7;��]�Z�G=D����l�i��<E�һ1��<��=�f�4�RiP=l��<h�-=�q�:���X2N��j\�X�1�r�m�=�<���<�V�<4����:ּ��Ѽ��<����fH=&�+�3� =p��;Iq_�qsA=��7=����]�'=���o��נ<���;Su&���N�=Hٿ��*I�fn+�;�W=ە���i=�1�<��c=�\���k=�w�=���E����<��<�����<K�J<�J<F�=a��<튝<�1���K�<�|f��.��n��Q�)<:�a��G>�Q�9=
ą��0�;��T�Q��~�׼8��<��=3�ۻ��N��DO=k&7=����R%���U<�f»f&�<������=��0< �<gP!���<Rm��'q��u�����;��<_��;�� �;�f�D;�<b=85���<������������; �=�u�=�A�<��n�����=�u�=���Z��<��O|��˰�=�\w�BK��.:����׼C����[�[�
%�3�=$r�=�꼩!�<�A��=}��}�;��Bk�����܇���.��_�<���<�Y,�r	P�>�<�w=r�;�{�<s�=C����&��l*�%LO=��"=��N���l<�!5;��u= �w<�a;?�q�S�U��m�A|=)"���O�]�_��gP=���B<�{��X��~?d=���G
=��;m=��=�5-�jE=I�ͼ�����C=���u8�}C;=2_�<��=[�o�q��k�=�WA����yN<4������}��̂��]�<�Ǟ��<�V3=�58�k�C���S�LVA=Z�s��a<�]�⼩a�x�/=}��;w<�O;��r=�*�!4=�0���<�oX���3�b�u=k<Y�=�m�<eR�g]�<�}��>����ļr�k)���G=��;15H=�̻�V<�<�ἶx=�x�
[���<{��<����9a��'�<It�<��?=���<(�?�})g=Zt<p��P�;	��;W�)=���<㛼�����;�'�<�7=�_=���M��qļb#���[=�;!� |1�fH�>�s=)�=�G�<B�-�r۰�[wI��2{:��R=^̕���=�A=�ʼ�T=K-=��h��'B��$.�;T�<Pvx�!h	��m:=�'��tM=�2�<��<������=i��$N=7� �E�<�"�B��V�-��<��^<.�b���;�˻�m.<J�<s�<=HS)�:g%=w��<]G2=ʼB�Dͼ&��B�S�;==T\=)Q�9jt=u�<��.=0��9A��#n�<��(=p�6���<���;���<;�S�@��<�1=��i�P_~=��<E��;P�<�|��S��\K��m�8�=Ox/=�ӳ�W<��;e'd����������<~�2=(��<V-����<kF;!���ù���h��Q=6�����:���9�$�<ּ�$�<� �<��@<J��e$;q2���0=b?�<��=�5�;�&�#�j����<ȯ�<��>=)��<>�T=���:�S��<�=b�;5�<.��aڼ�ü@�;���=/=��w>�W/D�*m��:=�B(=c�=aM�?p��E��<]�<=�uۼGD=�a'�h�<=������f�n$��i=�
<��ҼN����.=ځ�P�(;�;$�X� 3�����;&�v�9�6<�3_�20���N�<�<�;�+=H�/�:�;)D��A&=�l�;��
������<�2���Zu<���=�<=pV�<5$
����<�_=���d��<Y�!=��<F�ϻ����.=�i<��;
$�:
U<t=�Q�;+�S<��.�L*=&=�����l���g="u�<,���T�<l5<O48���/=���v��<�
��w=X-.�vwQ�Z�Y���e=��	�.@�<+�?�5�*uӼ�CP=PhB����\|N�3�"���<C�O<�����x�=b5�<A����=�����e�o�|=�y;w����>=�=ʖ����:�m%���o%=8�<U��:xnļ1|=�\�<���;��1�bE}=� ����;�]=/��=�)m=t�<6p�<��B=��7����<�7?=l^�;����~��� +�j�e��&���R��t>=��;��=�D�<i_e��μ/�<�(;�Z��E=7�:e�⼭�=]鼻�uI��G=D3���A�%������J�b�ɂ=��V�:���G�W���E���<�*�9^	�V�5:`=H.6=A~-�~$,=c�`;��A=�[�������X ��֍<}z�^żfσ<cV�.�=��*;��r���|<6=�ŀ��D�<�����a<�
�}�4=|��"��<��,��\[��==�7=��_�; Ѽj f=L_;;4��!�Ƽ�w����z��!�g�� S��R��=	�j=? ������n��2���J�&MR�,<�T=�tg�<��:IA8=����O1�M��2G%��� ��j��O���~=	�輴a���=Y/ü���;�*a�N�뼆�q�IO=�<���a�����p6M��}��[�<�;�Ik=K�����=R�R9o�0�o^=�n�K�V=wd=(��?8;��!<��ˏ=U�D<׍���<Y�=��8����x;=~*��9��?H�;��2=�V��|��`<�8$��J0=7W�a�)��ͺU-����<�R�c�0=ޛ!����O	N=�=~�}�����S=�o~<#A���� ��<i��<	�<
:=np��7�<�:"<��:�#&��<��<Q���� =�e���;��֦������<�Z�C�,wؼhN`<�B�4�+��X/={!�*R=��
#�O]�=Y��Ƽm��<��s=��	�_��;� ���2��$z<U>a=�6μ��:tb�l�#�<^��<#gA�x�
��3K=m�Ż���;tm.<#�=C��3��<2o=~��_��: ʼL^=5&;v�	=���}{n=`[���=�g�\y<��X��v�< /F��ch=ʆ�<���<��P=~'�=4�!� !=��=|��:��=���<b�*�P�C�;;��< u^�'YL�xM <�'=��&qH��
ݼk�<�8;}���>�a=,�����X=Y�j���»��T�V��<7[�<;~~=-*���Qʼ�D����;�-�<��F�t�s�K<E*�<[�i�e����=T}C=�8�1�=��ǻጐ�D =��=�2���7i<��9=���9V=��;4�O=e"K��q���@<��!�p����l9�� ��<���;9�;���<��=7廟�/<��l,�|��<�~=��y<<�S����B�=R9]<2����=d�7��T �Za<��2���1�t=E�A�柗��y�M���!�<�c�d��<�*�yD�`'=_���\F=��=:����Ҽ Q:=���;��	���=�"#���üo{׼r'^<��/=*��"|�<��;�8�;�(u=���9�F=q��<�ζ<?�n�82׼�4�<�m9O\�����7.:d�|�EHV���R�!����=X�[<;�=\/����<�./=��c=ݣ+<=�2�Va��䘔<�Z^=~R���׼
�j{P����w=feC=��X=_d���T�D����<'�/�0����7�<^=nԛ��Ǽ��ǁm<�����=*�&=�/���%=�b����;['��t��f��;O�k��
�ӓ�;�e=aSM=��<!��.��<��2�"�V<r�<h�7��nh�<<N��8�=�������/=W�ûɄ0�)�=c�=<+)�pw��: ��\$=F�=o,	� 7�����;=<�=2!&�Y�=R�]�<��B��nS��7=��<Ǐ^;T#�p@=q����Ue=���<�Rb=&������6����|���㼢�.=6|D=_�{<�����;?����b����N'ʼl��wq�:��$��8=ܾ�<�[ =|򘻭�"<3L[�$VN�f�+<��.=U'4�#A��B���?�V?0�Od=�
�<�#(�a��&��N.=<xC=`2�<3����v�L� �H=������=��x�C�Y�Y)��un��7�^n�<c�껫.�<B*B=�!;3g6=as޻���<����]<��Eu=ev�<j7"=��ּ?����8�V��uy�<��L�ί�	����^���<�ީ���¼�J#���<��ȼV~�V�I;B�U��:�<4x�:.7���j�i�k=L���<�=~ُ=yP=�=呻��8=	�=k �<�Ӥ��0��ӭ<��	��c��I �LYn<�- ;n�E�ѫ@=.[���:���z6/=oq4�!�j���#�w8=7�	=W\;����t�<	㗼h=�[�<Ќ��_���̻�����{i;R�<RY����<�<��0=�X];��k<6��9�� =���ޕ��h#=���J=��|M���<��*��/%;`����ƽ�i7"�.�(���V���:�,��:@(����=D�M��:>1-�0Y<�Gj���<m*���Y ���d=x1ڼȸL������X��k
�Z� =�b�O3��=�<��P�%k�<l�&��T����"��<����ۅ���p;�O=�w=o�Q=C
2=W�=x����;!=�K��	=�q��`�����=wQO<��b=E�������<�=	7�<>[����B��	�_寻�[ ���=	T�q�j���K���(��	m=�OҼ�g�<��#[����»����:>����:�G�ޕd��}��-�=�yZ���L��)g=?�;H�弊q�<���'�B=6.��ty��Y�S=9v<=J�=�E�=?*̼��=�?�����<ɟ�<��=I~i;�2����/C�����<��=$e���fi;�A���;��K=_s�<N�<�(=ew�Öۼ��"�͗�<�,J=Y��I�=F`�<QN���;/�@<�<
m5=ǭL�Y��;,c�r�1=��5���;�xB=ͧD=Ȯ�<���wͯ����;�'r?<��;+̨;%�;�?*�Z�q��#�o�<��0�Tk<R�!��OI� � =���ť;\g�;��,�2:6�"=��;P�<1�q���E= �߻G��<]5=t��;�<����:���_*�<V�F=E�6=Fn <����2���^5��g_�'����e=v,b�+$*�6҆�0x+=_�<#g�<��+���i<b`6<���<|"��+�<�I�<?T=�i<?������3=:�ڼe=��f�+<�,�<+�<�RA=�{�<����
<��i<����@1����#J��|<_�$���/<<�j�l1b<�K=�
�w��<�-��懺�!J�N*l;� 8=���;>�<Z�����Z=I�
��g'<xZ=��<�g-��P�=I9==���5�5�
�x�hJ*�3d�d_�Uld�ߔ==�|;֢=�X�<��9�]Żr�=��Լ���:$}���/��������o�<-�<��;��!�6f���a�䤦<9�׼�V6:�B�<tI�;� !<j�F�!�@�1w\<"�d=x�.���<�O��;	�;�  =��t=eB��9=љD�h#r�˚B�^�A���;��B�w��<ʪ}<�ɼ�H=ڶ<$4�[Ck=�ʇ;4t=b�n��0�<���c?�!z�<��Y=u�Y=�=�=s�Q���2���7=亼���<mV=��:���;���<u��@ge=��<��J<�F�<����e;��U=T���n�<=�&f<B.�<�=ʜ<��ټ�P���ʼ_/k=�Q4<֚�<F-����S�N��<�Hp�PR�9.���$<F�D�񞺼���W����:B'<�x��<�O:�G� �j�э��R&=�š<�7��]=��G�:h��S��<��<���.�S=�A>=& ����=e�K=�9�g�\=��V&���=��<��ܻ�����J=xR<�o�<N��j��k>�� !<�&�<;�L;$�H�Ո�;����^o<� ȼ08 =tj������$=(?��m�;k�(4�<�ͥ<B��<Ru�<���<���:�ɼ�������;+	~���<�T����<�#=f���h��<*�;��J<<���cQ=�j��Nq�<@�.<�!�����������uj=�%�<K�:�����lּ�qL�?�@=b�"��`�;�!
�9l_�a=C��<�D��<9�e�f�=eGm<�]O��M�<
=Z�t=�=E)=M|<��<?b=�= �.��3Ө��=��_=��5=��w< S��l�&���P=J_������Uм�e�q�,�mƻ��={^=����$�=4q��-��� �oR=/�h��C ���t<hx�;�S
���,�moc��B=��=��Q��;����Q��<����1����qﹻ��I=��+<h^��_��
�� <ؤ)<8(<Q�����O<���<QĒ��~<z�k=c�'��<�<G=���S;%�=�1<�s=}�=@M�;�`=��N=C�<ޔ=���n
#=��=�I	�8�S��ɼ��$#��o�<!��4޼b�Z=������K=���<7��4&=�N=��N<�]�;��;=���j�;�"1��9��=�=�mü񭤼8���y�H�W�u=nғ���b�=�~�P<��<<��;qB���4=�jL��c?=_��I��<�}�0��;�nF��q]��I=�m�;VI�ۿ�<w��<f$���<��9=@Y=��=���0</�.=~�T�󧄼Z]�g�d=��<�;:=�b<�[ټ=D�<��<��;=�m��v��,=���=���<;�x<I3=8��44���<�\=�|<�lA<��"<�D=@�0;D|`����<�'y�)��������<��=Ydn=5=�1{�}o<{=֎=�:��<ID��K�/=�߼A�M��/R=�'��
'�z?G=V�=;�=α�;����H4U���ټ�{�(�A��'<V}��@�Ջ=C�H�b<��k�<�Ӄ����^�<���<,�!= 񥼴�Q��P1=��<�"L;�x�<���������h�)�1=��^��Ԋ<Ĕ�<���<�=h�f��@=l=ծ};'A�&j=���������<�Hj���m#=��b<���C-�����6�ǼB[?��}]=7Q&�V�<2��<q����E������s=�)޼��˼u�=� ���]o;�= I���{�;3%��ʿ<�ӑ�V�=�;��e�G_��3ߠ;�<�����^=��r=ó�Z��<V��9|���r<���;Uy��l3��lyb��[ȼ��7�NK:���3=dٴ<��ȼ̋N==�<䐼DW<F�����0=h�m=&�޼`m.��eO=nY=(4�βZ�TI=D{������U�֊q=T�<�L��#=��Ӽ�o�<�V=s�,���=5 �<�8��x���
=D+�<��"���ۼkY�<��<�(:��8�=�}�<��h��O[���;�!�w�=�=�%@�H��<=)=㖸����:BF�Ad�<�<t=�a)=xhu���Y�Z��<O�<�)��+<l�q=�E1=Y�(=1�L<��e=>�]�I��;6\<=5�@�,N��\�u���ə =�a���;�;�=op<Jp����1�%���&s��sK=%~<�{�;�X���W����<dH��W!�<'7��]=G7=\Q��rL��2a;)4=B��x�= ?мM�$�5ㇽ5�B=l��;"C|<#Vf<�'�ym �Z�K=�-�Wc�R���T�<�W��8��H(�[�;�Q��~b�<����-%��~<� �u�'=)={��<���������p�(�䯼���ɱ�<S"�������<Mv��	I=ʥL=l�;Ys�<�5:�64;��׻�MJ=��¼�(�e��<x��<���<�k��>� ��<�
����<�NH<N����i�<�-J���F=�7?�%?%=@��<B1��|�s�D=}Iv���<��M�GV��ԯ;U��!��ZAy�u5Y�-�ӻI�T�����;�%\�������Իt�u=�=_�C�5=k.��N��>�K�<��=>.*��=�k���y<0Xۼi��<hT�=|�.=��=5��Rx=�[N<�w,��yE'=:\�<||Q����<C�;��y=�NU=�U<��9=/ 漑�1����:<�d$=��|<�պg��<�ּ�q������~|��ʰ=g���$�<�1�.���7V=YfP<��,��M= C=�bl<�0=~#�;�v�<W�;���!ͻ����^ѱ<�j̼�<p��ϻf�.=Oֈ;d��<ɤ<�#�<��pC�<H2��Z
]=�w�<!3�<�gk=}3�<�8;&W]=��"��^=)�D=���<�Gj;��=�Up=�^j��#�w����<>��<��S<K�E����<�E=¤ܻ�������O�9�1��<Y�g��]�<�A���=�CǼs��<��	��a��
�|���<�=�ǼZ��{6⼳�=F�=�)=nZ1�9�x<�F�����`+�<|��;����$�μ�[���E:�#�	2Լ�<�D+�1}b=׽޻�B<&G���};V̗<�Dv��(^<	���V;�O�>O�: P=Fug�d��<�eP���=N�N=��,����;��p<\�R=%���B
=5�3��+k=7䌼���tNļ��L<A��<��=S:��P��K�=\)��7켫ψ;�l=��=��<�8�|�$=��=����(��6𻫕���uF��o'��mߺ̛T��7=hZ|���Y��D=#_����~���g�EI���_�;g}N=_Y/=Ɏ�<U��n`�;���<�@=o�`�d�<�#�����Or�7��
.C=�c,=A���X:;3�Q=����+d=���<��»lc�;--=.�"=6!��'@��
n���������,0r=�X=^���:���[��<
h=೽���o1=�XL�s*=�#3=i�<U�<����=�z2���n=�~!��=E�Q<&�'=�~��2�a�\=8�(6�v�YB���(�X�5�	h��	=h���9��<�!4=��]jͼ��+=�ꭼg��U=���;�'1<���;���<gN ��fv���;-3��j|�]�=��<�<�<�1=7�(�$kT<�&�9���=��W=�q�<`-�gT˼�xB�]�����<:j�<�G`<����(��_��/+�7�<��<k�2=1�*=�=	"�<_�<��b;�7=�F_=t@8<�5=�R�^�l�V��<��;=�ᔼ�FT��vV��꘼�����ߺv.(=��<�++��
���P�<+=��T<w�M�]n=�Z9=eW����
=md����Z�
=��<���C�����!�����P��a�:b�ջ��f�����5Vq�peR����<�F =P�H=���<��.=��=0T=�Oi<H%����;�[�:%:<2�[�8G<.W�<�T<F�(��A�U=�,�<GG=�<�7��L=��\=�ヽ��?<��F�}�=%r
=����(�<��.=���;��
=9Nļ%!:crZ��I���<=����S���=��<��%=/�=8=r�N%h=X�[=)Wa=	JI��>]<,�<�;=v���r=`�e��*�<�&=v|�<pܼ?v=?�G�'�V=d�i�)��-=��ļ�=Q| =�I|=A����!=���z��<VG<&�u�x;|=��Y���<=.�M<e�S=�)A=�G��o�=���p���[�;CU.���W��s �M�Z=�&5=i1�<䶶<l�=�p�<G{�<缿<�a��,�n�'�{<�v =��׀���}(�M4S��ʅ=��=�1�<� �<�L=N�=�[�<+�k=�p� 71=w���/=<~=�?	=F�O��LH�:�!=�F=�_<g=�)=f�=Y��<T L=�ȟ;{K=����}�q�<��p<���<��r� �Y����<�7=hEU=R ��=�%s<V�<��2��;!;��.���g=%<s�0A����޼F�=LX=�e0=��y=��~�&��rk2�;[� $*� p�<@h�<J���-=ԍO���m=��=ϻP=�.=��.;��:KR7;��]����<�5<j =���<<���r(<7K=Q��k�=��t���=�3�<7�O�|��P�<,������9���(=�g[��&5<|��<��S=����l o��:~V7���<濽;����/=��<%.=z@=h܄;�0=��"��膽�8�;y��<�:��]S�����)�ȼ,���z������ ;[�D=Hw)=�?D�`t=H=����%�=MT(=/��<�P��ҋ�<o=�gϼy���/=:�<R�?��;p=y�<�"߼���ý�<C`=c��<��2:��*��dL��H=�ó�B

=��D=�h���s<&F=�e=����1���<��L��� �	=;9��R�<��8<��E=�H�h-;ғ����E�R9�"�����o���N��9:_����X�x֖=*�&=���<��L�m�<=꼤�=[7ƻ��'<M׼�,=��u<�h�<]#+�P�Z�r	<R�#=Q?=��@=�:&=����;�z���,�ٌe����m=	%�;>yY�#�����0�+�Љ�=�4=M�;0gZ����<��:�)��9���ݼ��Q�ǉ;NS3<�L����v<�%�;�(�<�%�<�g�;y,�'�n��zc�����X�[�}��� .�@T�Y=tm�<�r���Y��˻�Zi��v2=]%�0e=8g"�+Ǎ</HA=�"ۼ�!�͔E�F��;"sH=X΀��{����=\�<��j�lSR9��.�|���	
���ػ7�==@lQ�5�=�ë<{�Y:|D�=�w6<8�K��ě=3W���j+�__������,2P=Y�<T�J�
#�<_0�<7�:=F!�<hO�<��D<�p�:D�M�7�<�K��qq<2�Z�-~a<0�U��9���(����N��[Q=dp����&=HAݼ�h�Y�=�S�<�xb=%O�<q�"=�\;�;��Q�f�=�Ҝ<�|< ����<��\:_<^!���L=��K���N=�D;="�4��8�;�=o�ở
�<�ɫ�u�=�A��%����W��d� ��w�>=�7(=�%";DV=uy�<p��="�]=�yB�ܹ�<�)���w;e�<s�����<n�k@�<�Q<T0@<IF�b�H�|t߼j�o<{D=�-ּ��ۼ���;��M=Qt�������L&=HL;x-ѻTJ��)G����Z�$}0��J�<�s�; ~��|"=��#=E��=/;���<�d^<g�=v���Q=�FJ�!�==�H4��xb=oH=�E=e=hj�< �=��9=t�=�L�<D@�;�t���nH=�\�=U��<(���μ��s����=f� =�]l<��O=��X�[�:,~�����漗�;c�=�^���Ƽ᭘<ha=���<9�`=ӳ�c�0�:�s�<M�1�)�=4�м����F�<�Q9:��C<9H������ô���$=�R.={K�<��==ݣ�<�����x�=ץ��b�<��N��w =�}�:7�C�p!�l}���@��i���&;/E=��$����E�;_�:=�)�<΅�_g;"�a|U�H����!�x�n<׆D=s=�=h�R��#��;�2'<�
=����[� ���נ�<�T!����<_{��-�<�b4=A�5<i���Z=<W���<�1T�p>�.
D<T@ļ�*���E=8��:
�<:'U�?����Q=�)���=r�ǻ�ͺ)U<�P/=�9;����l�� <�H'�if�Q"���_��M� �=P�������y�<H <MD�<�k:ϊ鼯F=n�P��N=�	=����;��~�g���f��=��f������9�yk��!�Sn���KB�RZ�e�<��=P*l�3�,=/
e�تG�0:�=~�g<O�O=���<O]y��\��� <*���g�<�վ��m1���e��<̱�;<e!���:�F=�P�<�Rd��Y=39=x�)=9�<�s˂;�N�������;<�d(ݼˊ=�Xk<���� �yO�<Y����NU=�V%<ʧ�<�:=<��j@�s�<rYZ�s�J=�����g�/�!=�\R�7�����=5���gr=f�8=II���~<Ӫ��N��	����: =@�׼X��<B΄<r��9�F"<��=�룼�VE=�<8����I�@*='��<�G��;9�ֻ����U�K=��M;�,C��Z	=<�<�A�<�
�<\�3<�[U=C��;=<~<�e&=\��<�0��Z�=�:��� <i����<#]���b�0Z&=�=�<\�J=��f=��<|��>�M�D|0�Qu)=���=�<D���&="V7<��#<k �����Q�<"Xż��C=!=4�1��V?��I�%�!<�����R��$;N��<��<v�f=Ay��ݗ��޹<U�O=�49@	G=��!��3^�	�K��{v������	���u=-W]=��k=}㼁�=	m'�8�=S���/�?������]��-l���|�Q�*��(g�Nkټ5�Q=��	�.=�)�l�Z=��C�M�q�F�=�	���=�d��n�
=��e�1 =�^<��5=6�y<?�;X���?<�ND=�h�s��r~����=\�-�A�Ǽ"#6<�6�6)y�j}N=���<��<:`=F�i=��,� 10�l��<�����*=m�!�0w�<\N�<����+��<֖��j�T=����������<��<����Aü�$����
����h,g����;���4�o�O��^X������4<E�=J#Ӽ�
�n�}=��W�n@�c5��������;��=y���W]ȼ�߼f¼���<&��<{|<�5��3�T�G��t��zL=��Q���<��C��Ȅ���&=����}�=�<=���t����׼�<�pм����H�"����{�N�N����q�6=��<u���}=���<@�D=��7���0ł<3ir�<���IFF�w�=�W���<�*=^��<[޼:�ҼƆ�<�襼�zc<xn;����=��#��"������p�<V�d��i���˘�_K3�������Ԛ<q&�<D.�;	��<v�(��=S�d=C��G�g}üJ,�&G�;­���F=қ��]����<�弶���n�)�1�/ �<7Њ;U����F�2-��&�y/��CQ�7���Kw=9v=̱�L�$=n��;�� X��5�M���ʻ$Q<� �?�V<��=�-������Z��������;�=������=�=��<j�L=�`=����a�Q�F�ڻ���״�;���<��м�m��iF"�3.�φg���5�)�؃7�F#����*����<�3�<���j�=lv�;���`�l�
��<H<""E=?��;S<��F=��Q����<�8�<���J =��/<��.�<j��<�=�����<\VH<ׅ������b=�==+�<��=KUK�m�Լ:!
=�z!;my=VEպ����+��<@�q�0�<�(_�V ���<4��[����4Z=��5���Ӽ��<I�=[�d=qb�;a�<���:�EF���g��H�<Jt���*=>�D=B D�*��<Z}���=���<�UҺ,i�<xt�nTu�U�(=�4�<�_=<
v=U�<�c=S=;��̼W=�<���<��Ɏ��~�KtU=)�}A�U�O���<��X��n =m�R�W	����<�����;��<��� G_�b��<z
m�v�%��ҼO3=�Œ���?���>�����6�;���rp�<w�E=�k.:��<����j�<�=<�,=#�y=d�I=tS'<�J	�(9�ͅ�=�_�B=2�����U=�t���F=jtn�$Ƴ��f#���޼�eO=Jw�=n��&O��-Y��ɸ;r[�./�<y{=��f;�P�>p��S'~��Ԭ;�..<S�<o�Ƽyv=d��;/��;b㐼 7M��#<����<��X�@�R=VuS=���ԙl:T_����J���6	n=~-�<�x
;N\j���\���!=7�\<�6`�Qa=��<�r�Y�=��g=�a(��,;=�Q/���һ7�ں
X=�
ϼ.d����/��ˊ= #e��c=&�c���;���<�F[;��4����<�#��X�G=��Y�����5����&=i�M�ƣ����<�+=��bņ<%�y=8�=B-��P�=r��<��#<�=�J�􈘼�_P<(kZ=���"��<C�<��G�bn#=_$=���y��������p=1�=����B����=.E�<�M=�Z�O�ɺ�\1<�1���`b����<�oH<H#=���<]2=�'�<BOm=�ʨ<Q;�ݜǼ#� �~=_�@��ME<坌<N>*;k�<��3<_US;���H��~H<	�@=T�4�'=�'ML=pq=�����(�y!=�=���=!����⼀�q�C�@�G<G_�;RV�俲��"���/=\�:v:�@�z�<�u��pG��E*z=�b$��z=��G=�>h���z�D�A�P�����G�	8���n7�[�$=�n�<=OD=�p<�B�kA>=� ��ؼ��
<��μ;�����Fȼ-S?=�4�OW�<��?=7R`���V=�"D=0L=lH=��5<f�5=�C�<r�Z~�z鷼��o�1��:<��;�P=��_==�<9r^<մR���<<+����s�p��<�Gb��»�μ���"�ӻ�<=��8=�
�<�j���e_�<�5���Ct=����
� ��=+�@�����M���=3�)=
�";MT=�Ew���=u�<�=�ڍ���<�I�;xx< @=W
 =�d=��=)L�<�)
=��d=���;wl��D�w=�-=�"�xVԼ���<�<�H���f�����<��켂��;8ct��-�;A�=�_=9�$�*bʼ5��<��q�%�;��A�v�����=}�S/���e3�
�="3J=�EJ=E��<h���=�+����<��m������<ӟƼ1��O?=����k�<^�=3������;��a�3T�)�[=�4�<��)��"6����<� =���<гJ��I4<�u;�%,=1�B;�ἧ�����=�?��ļ�-B�ɧ9��_���޼��F��n�q��⑸�E=)=9큼�bB�x�s��Z<�E�x=�D⼤G�`��<Q`{�]���7�;��<�`�<R��=�D�k��<LP�;��3���<(i3�2��;Ɔϼ��c=�%��� �9�O����;�K.��	��}@��d==ʸ�;�F=�K�>��J�*=�$��.H��<Ĭ?�C�=�>=�b�<~�%<�9_�}=o�C=�����T(=�ٛ<+��;�e=�Æ.���r��n<q�A��w��wm���3=Yn�/F;�K=�S��K�D=��P�%G7d=�'<������7�_�v=�a?=l3��H=���d=p�l��H�b0�RK	�:V�=��Z����<p���=���I��焗;��K={.��s�_K3=�*<���<��L��G����<�8#=�DK�M��E=��<И=(/����:0�<�L�;�20<�>�<��[���V=��X�=�F��ۡ�#J=|��<ǭ�<&)������f_�6�?=�<�<�6X=S�J;��d�fw�������lH�WՆ;�6(�o�����<�&�;�	��V�r��إm<RmŻX���j^;�6'=�Gj<ӆ>���<�=,��E�.�6= P-�:%��.�A��Hc���-=�=�k�`{#�B�m:�t<p�x����<�:=�YX=������_O?=�����ؼ��6=��<��=�d̼�fc���R<�����4=���<TD2���ȼ�d=w�^�/Eʼ�#�<�J�<��L<�%x;��1<��<���<�)<��D����<�h�;$��G�U�zb��$�K�=���c�k=����e�<�EԼ�9���db�O ��t�!������< K�<�A�=p�9=戒��\<焧<��*��������� �;2�=�Sy=x�Q� �]=Ȫļ!����L�������<Es����<�����aU��z=���<ER�'��<p�/��-�a/����R��c*=���<���</8��*ռ;�c���C=j�$=�a=L)��$�<�Z�<U*K=��U��K=rA��J=��U=2�R������ʟ3�
��</�޼�*U=M�),W��k�<�$=̓�<��j=��X<��%���+=׼S�=�&���(��ˍ<�5$<Ҽb����,S��0����;I���95 n=r3=���<���:Ǻ�;pH��_�#��:J�S<��!<!�����P���� =� :=%R=`=�<����D<���;�]<c(9<7p�q�=c��N]T=/�1�K�,�����CQ����<(�+=f@ =��N�<�#�_��;�;ϳ0=0�?��g��#�<"l��U�<\һ�6=V]\��dF���=U�Zj=H��<k8K��Hһ�p0�ݮ	�r���tY�!<g��U<���  ���:��2=�����7#=��y=����~�����������;Yc��企�μ��6=b�Q��M���O =Xq�����<{9a��=�t=�<뎁=���<�����X<�GK=s=�,I<"my��9��1�k'}�(�w���<GZ������>K�<��ʺ�����qI�vT�<�`��=?C�<^� :<=e� c��#�0�]�<�f����~���<�贼=��������	=�=<U�м�sv=�.���*=�0���/0���<hY;S)�<��2=PF =��<R=�}<?;���/�<��P=�fA=;�������
<t�U=�_���<suD=t�1���/�% =nh�N=IV�=<O�<O�.:߆�< �<_o;L�'	����Z��=@�<?���ۇ='� =�����A�:}E/<�k)=��E<�F<�y	����h���<z=��=�Lz;%�<9}����<�O �I]㻃v׼�5 ��L���c.=�(ռA�=�u�<]���ط��=}��-�<���0V�����<���Q��5_�5LX=*�<3�^=�~.=���;%<��]�0�Rږ��K��!4�;�;R��;���C����I=�9��������<?0�s����0=<��>�缈�i�� =�ĻqJ\=B��<�؆��c,�!S�<�����<~9�Z��MW=��=	���e�=ѷ�<�z@��_=eA�U�s<�N;kٍ<zT��4����;�໻�Sw����D=��R�̯��? F=:���c�y���?<�V=l��.Lϼ���_$=��<B�=���<��vu<,C^<q1==�+��щ7=���Y���~@�S�r�rwI=����K�=9W#=����#o�i�@<�r��2=��H����<���%��< �H��}<Z����⾼�"[�h��3�����!_Z�H ��fo�:Y��/��<�'�<��g��x�3�=��Q��I7��cj��4=��������9��CC=�M@=�"�;=�=nPʼL����*G���+9=�Z�	A=�����q#�<�	 ��L�쳼�ed��%�<�*=J�Q=R�=�|�;K���~�<�1ɻ������ڻR�;��F)\���<��0=�����:9��=+iW���o=��)�;A?=gB�<��r���c=��1��%�:[!�<-Ȫ��<���<
w�<yť�����f�<�@<���<�q��=9`=�dܼB� ��F=|C�j=Z��)���I誼�;>� <�H���G<��<@Z=!� =�=UN=�ە<s��� �g���=bB9�?<&�<О</�c=�M2<
ɞ<&�;����'2<�hy<t"ʼ�JW<��Q=��<�1�<"b=��<<]F<���e=�R8<�6���3�ZI^�sk�`�=��b;r)�<���<�/=��¼��#�@2v�9�b=�yT=2�[=�8���#<��B���F=�P=7���9vF��2��*E�?��	<��<F56��6<��)<>�<�#>��*=`��=ѽ	������<%��r.�ޑ�:���m���-�ӧ�<���<�A����Ą߼n�==1m�=��=KC���:=�r%���'=,\����jVD=x�<��/�糖;�	_={y^�4(����+�Fm<�؝�<L� �+oN=[՟�VlR=���<���VP8�r��T�<w=�� �+=�m��Y�Amֺ�(=-i/��l���:�<A �<1沼��*=O�"�XQ�A�,=)�.=QR�N��r�<�D=��k=�A���(7=+�,�`��<
"<vU,=�D�aa�ye����%=���]�6=��E�<��w<�!A<�(H��Z.�X�s=[2=�SY=�������w����=j=d�=��
�R�W;�X;������=!4�(	6=�F�9�U=*�����d=q�E�7�6�a�<O=��=*�0=7:n�	=�_c=���<�=$��PӼ:�+=B9=Q-��;=lar� X�<��;<�G1:s�Z���]���ͼ2�@��=�IS���m;X}���J=����9 H=��l=,HR�h1<�&c=@Y�:�\�<�%f=C�"=��Լay>8_��K-,=���;����M�<�k`�?֊<n8���=0=�n9��'�<�����K޼�m%=-� =���Y��<�AG�B�.=����v�<0�L{�<���<)��<��r��$�����l{=*s��g;�x*=:n��w-�_0���3=�ޢ<�ż��T=���<΃�<�:=F6<�E]��.˼=�&=0Q=�V=�Bn�	�W�F�=k�<�i�QP=F�߼��!�,f���=� ���2=^L=��V<��;�T˻$Z����<�9���Ŗ��	��D໻u����D��#�޼y'���p�tj�<��=&���z��H@���T�=��=UDԻs +�m^`��_R�	�s����-B$�S�μ���h�J8�=ڻb�<��S<��Ӽ��\=ƃ�<Dn�<�8l<�YG=E�7�8V�<Eo޼��S=s���+��݀7=.��p=���q�l�d��=�w�<PrB<��<l�&��+=�&��aD=�FN<�ټ�l��$�нy�~'=n����t�&�<t�?��%9r<����Y��r4��T���j�Av�<>�;�dL=��:=P�v�a�;w�=݊�<��<+�l�Z�><����xC'=;.�B�u��e=:�߼�<?!=qv<�bP�$�����
�����n�e���c���F=ೇ<���t�l<-����>�'::����<��I�]�X=��&=�5j<z�=�/ϼ�vE��t=@��<�>%=���˶;��=
�:=�W�<�F�<�qż����G�=����'=H9ͼ�{r;��n<v������<�������5=F�%����<
S=�==���н��]�,����<��)��j0=]\庘=XY�;|6;��H�/Ȼ�'8��G�<�bW<�g�<�H���<�<�{��L~<��A�b�����<��1=��y�j��;�]�=�#
��]���&ݼ�Q��=J;�`~��Ҽ�$F�ύK<����L=k���<Ǚ�{�4�u�Ỡ��v���Ѽ�-���<[=sO���=M��A�߼M��;���'� �i��<�a�<5��ㆽ��������ּ�d�<ʖM���ɼ1�i=G����0<�<0<+�%=�o+=.�:~��<�J=2�=/=%R�=��c��5_���=?��7���c=�<f�Y�D<ҖY��jZ=>R2��A�;SQX���=��=��\b��V;=�~=�k�<���;�\��"J=l3=Rz��e;=!=wy{��xA��;'����T0;������:	y<_S�<����7�ݨ:�S�)==�*=
s�?+=��-=�l�<S�/<�|R�"�>=�;c�P���<o�����c=\/'�=�=��r�;�=��B���D�����	�Iń=ӻ<����?�9=�8*�&��;�p�<|Y�<xA�;��<��n`e��n�;�k�<�V=��<�}���;���<���<�y;<�8�<�/>���*=�'�<Hq��:�<~�˼\Z���3�;ے)�D���ܼYVW���"=5�,==)ּ��3�]� �u-�;�4=��[������k�z7�<%CH���Ӽ���=���P�(�w�輟�:; 5a�]S�<L���P3=��E�K����	�;��6�,�'<��;����o���XZ�ɗ�EԼ#�=6�x�똙�C����=�=���;c��J%���=-3c=�yS���<*�q�k�D��v�1I="�=��J<يP<v>E=E��9	���Z]�Fф<V5$=E�]PX<F^����N�����<��^<W�缿�f�s͑<{X�O[�<2����v�2�4=kݲ<��;[�&<u�=��h=B"*��\�<O*�1Wc�1t=XU�<���{=���92�=o��e}=G�;4i�<��i��g=C�`<Q�s=<�O=b�q<��w���=	���t9���@=��%=R}=͞K=��`=F;����i�����~=��90s3=E1�V�;��K�)�<b�:=:y�<�w��gi=�� �a=A�=�cm<*�ؼ�g���|=p����=G�;1�8�y�U<v��	��<ss�_s�0����=�=G�$���=r�=��]=�>!��c������=���м�X�<�I=6 �y�-��T@�ZRy��]�<��Ҽ��="%��{���=tRP=� =g/G=c�������m-�-ȼ�#~��ȁ��bs=�8���R�<O�G=���<9c=J����/<\mQ=#�q���˼��,<���<�6	���i=������G;�6z=T�<����xK=������d�LK]�*!���8=1�<��Ճ�`"=��v= 6T=�f���C��%<��*=횭<��G<)�k����<jD�<cO=S;x;��C=�N�=f�7�`/�<�=bO<Lc=���e;8=-^�;[>�	=	_�
Е<����b��~λ8;=1�l=c 1=�D=R�мx�z�x *�V=��<K�κ��B�X���y���BF=�6=98�;::<
7l���輰�4�>�s<�	x���"=D8l;<c3�����=��:�mм�+��;%���I=i�P���������j�<�g0= �<��x0�/�h=�_�<6�����<�^�=1����t=�2=L���0���PZ�i�T=~�Ҽ+���7�#z���{�<��< �s=���<�y�����T�;�R���zZ=�i�<őj=�o6�Q��<����l|g����	�Q=�=3^�;�pG��qR=t�!=�(l�$[=<M��xX<|P<�q=\�n����<�Fȼq���g=J�'��T��!�<p�ؼ�!=�피������=�û�*��Ex	<�1�;�z<=
��<�ߓ�b�=��#=m�z<> �.���l;��D�<�;*�
�`g<�ߴ�<��6=�w��[�%�l?p=�y=%������p�<����JQX=�G׼'�.=����M=Oi==#%=��+<8����O����>=\pU��
R��=���<�L;���<�G'��k'�AW/={p<�V����(�NM�;u\Q=�lx=ǘ�=�|]<(�=�x:���j=�g�;H�9HԼ�o=-�5<�S%=���<�yQ=��;�1I�F���p�L=�� �,v)=C�=!�����q%A=��<�T���=�=(�����窒����;�����<�x�|�$=@IF<y��<D��~:=����>I�;����:T@=�݆��N=�]��lG����%c=�h<<�9���ȻU�s=�9����}���7��W���\�B����=�?=��漛���Y<�$d��G����<�p<��+=���O� �Lm�<�HP��5��J1=9<��J=�6]=ƌB��|�B�:|$��N:͂�_y=8A: ��<G"�d=5����t1�� ��<� �<�}�;$�<
�U���<��?���<='A��[=D�<T���t��<�hE���F=s��S(��L�<x��=�����n��G����=	�;j�<D��<���<��:P=���&/=*'��cX���L<�<u�t��<M_n=�&z=�;�<+�=�U�ٲ������7�E�j�ɻ\<"�|�=$���O�'��;������"=�ݾ<��弢!��0��r��\>=R�,�KY=g	�~=<b�F=�I_�$r=�=��;���<��"t�<��S�$�<;n6���`<��=#���LU=� ��M9=�������;���<���Z�<�ɼ
t�A��f����yH�")��=u9=Y�ݼ�,�<�%���i�:��<w
��b��[�<��=�0��W8��l=��O=��߼t[=�����<�i�,�V=[r��K�=�BE�;�;�����<�{E��w޼�8=��3��^>=$�,<U�7�c[
9�W�<���Q��n8<��F*<�y=V{���f=�G[��)�w���N�=S<�<Qm,�u�K���>=V�j=�%;�U��S+	��u�H=Ы�<�e=t�»��H=	R��L��;~�Ѽ�߻��<F�R=��=X氼��6����=޿=(0�:̮i=�<򼜎^��%�<�]�b��<
)=�_�Oƣ9�0<<�y,�\�
��P=�"[=90���*��m,�q~&� t �(4q=��;���O�o��o=����]�=>�#�{�m<9|�G�<��J=�G%=hs��M�<�b�;Uh�;a�^�>3�;?MQ�j�v<�d�B��<�=��=�r̼��=�&U=h~���z���*=y�d�	)ڼD>=��мd�W=p��<Lv�<�t���Oh=�m����-��(��cʼڧ;^����+�Q�;{HO�11������	=&�<P����*�I�N���W=��U=�֏�:i�<2�M��0��2�9�NO����<J$�;]�@�=��oM�*;���:=��=U";<2�ȼ��q<]��<��<C�ؼ���:ȵ�<JK =H�i=gbǼ�I��#=�o���̼�-=��j�6��<��s<�T���
�C�u��h�498��1Y=M8��ż.�R=�[R�%4=�f=	;��-��<>�=��:Q��a'��ZR�Ec���&=*�0�N�=���:�G2�87뼖� <�p:��<�6g���=0�q��e�W��;î<g�H<������e��ۼɛ�ƥ��W�Z��t=<�;�*�E�<6j=+L����<��d=W�=���<��<"�-�_j_<C=����ƻ�:�;�W0=Ӟa�E�^ʻ��żf�=��
=m5j<4���;��<�N<?iY=&|g���<� f�S<q�4���n=�U��Ȼ
u�ڕ!���]��T=��w�:�=y�=�@q���ۼH�k�tޙ���\=��k�$\=���$8,=�,-=>CC�.�H=�xb=�B�;o�2�Dvb=S�=ϾW<j���'�<��s=��;�G=�����^=��w:K�!;��<��R=�x>�N#��c%�G�=�M�<ug�X�
]�<�F�<r�����g��N��'���63�~��<�m��){Y�:�����s�ܻ"�=kR�����*�� M�cGG�K�e<���kʼ��;aD�<sNa�5<��>�=���<���<�4����<��7����<��y��_�;,R��W<��<s=����Z���Ӡ��ng<�L�;h�����-��)}<1�o�NZ�<�HF��X��w*�o�_=�<�[=&���ϼ1Z2�a�=�i�eE==�H=���i;�]=�9ڼФ��w�;�)	= �>=��/�~���$��j<W�I=x��=ſ��ʮ�:������˼���՞
=&�f�g�(�y�i�������y<��:� �<�F$=UN�����B�;C~@���/�7MK<KcL��AG=��<=b�:���&<�\��Q�E=��Z=�M̼���:�2W����*=�ڼ��<E,���2N=E�r���N�=��<�>J=h��ȩ=#� ��A=�e�w>q=�J0=b0�b�D=�t����:ji��q1==��F�<����Lx�<�=KKs<����}�]5ּ���< �<K�ψ�������<szü7�T9��%=��G�J�/�G���<��;�!�=iF���k<=~I<��;𕭼h�ܼ}�=Y�aܧ<H c<����� u����=��>;�f{={�?�c�%��E+=R_��?��l=`�`=R�ϼ�&X=vn{���<KX�;LU廬����B����.�����!==�B��/{3=�`T����;�S�<�7=�A}=:7d<��N���
<; ����j����Ѽ�z����^Լ$[(��l��$G����uA�>�<�/���꼘R;��`��I�^������j�ຆ<$�C=�}<�Ƨ����;��?��웼1Ƽ�/��l������<�l�<�9���
軼�0���@�;䁽{���fA�j#�=钅<6	=�9�;�Y�,�=e�0;c�J��wE���!=��!=��J���B=5�;)�����e�H%=;��m,����<��0<������t�H��<�S���<8��<eE�Wys=Et;�0=�I�=	T�95a�<�R=B�<vQU=���<C);�y<sr���/=�=	S<%�G=C!��*��N�$;�������R&�:�<��1�Q��<���<���lt!<'hN=lƌ<�r���a��� �v���i1<�ǐ���<�Ρ�F(�:����[G�:�D<]T.��1���$��?�k�(<K�����I=}�U=��o��Mf����8<�����U=?c=d��~�<��W�a>�<� �<��Y�~7p=�������6=2<����<Ս\�>=�;�<ڃ��6;�
<Õ<9�g="Ҽ�dS<{m<i�S�����KU=���<�c�<����?K��*�␫��f�'i�<s:�gO�=8����<DW*:@�4���i=f_��ʐ|���3<�g ��H�_\�<�U�FIu�;�8�oM�;�r;=��<z�<��7�:���o�.=�Fr<�X)�~�;��o�ؼ�l��9 o<�:1��k�:0��<�o�D�~=[�]���t�����;@-=���~�<P�S=?=�L,���|<�+�#��igQ=�=����I�O���]��5�&d��`s<?�8�A��<��V�bu�:�.N<˅]�����(G<���<EB�<��<ܑ�<�oW��|2<Pv<<�����K��Q@=Y�=nE���<^��D�򪀼H��9R�����=zW����<��<�O=)A1<C/ɼRk=�ׄ�U��l�̼�B�h�a<h��C6���5=�#B<��1<L(D=�m��>���W=j�W={��<�G�=J�;���;�<�M�61-=h�=����<� �Z���e=����m!��(�<��t��LN<��<�5�<(Q ��z<g���
'�Ƿ<=�%�"�e=�c"��ռ�|E�-��<7!�<E��;�-��:i����3=�p=XI�%�.�p56�3v�<�;�;�p���Ƃ<̓z����8_�<�*��o^�eQ_=��a�("�<�]����������)�z�g���j=/�< �O���[=�WC<.蕼 YW��5���q=X3,=a��<]uV���A<OlC��k�;��<iwh=�Ac=�=�b�<�t��_��=uм'z;�o弁U�<�f8��μ�q<�;��%=	�E=U�"=�g��H=�>5������U߻��V=GQ=�ղ��?u�<.*ؼl!�=�f<l��<�H�;�*⼨�����<꫾<�ej�h�)�)� =�:�\X�5D=��8:�#O�m��}� =�<�*�F��<���:�v={�s��bc=�n�<jNj=Wu�<�O	��]0=q�6=�(����$�[S�<(��<�-N�Ѵ<��4;p� =Ν��8L���#�+1_=i������;�7���a�f+O=w:�<�:P3j=C�<�[��Nż(B����0�k���(��J�Rb@�o4j��6��<��k����<y<��@�Q��<ä��J�<��<��s��=�I�7�&�DG=��q=� =mN�}ɻ�D�;CI���,[=˶^�r�C=�g <��{�k^�<�M��m�=E�:Wס����<׭0=��8��	=fg8=��<��<pL=G�<���<,E=����#��C�/=�P<"�&�0d��̶����<��ٺ�W=R+�� C���K=K��%&=Ȏ�<�ۻeU �%�5=�"�g���u�<�r�n������<�މ��I=�*	��3M=�c����<?��<�P�<��\=f-�;t�1;#��2�<
:�=�E�<!�<(�<�.�8H]�W�]=��-�ީ2���=>�)=��<�T={��0�<}S�<�W������:=�=���7ƈ�'�;��=,u=��#��Q���3=Gn�<��<a�<˄*=1)��T�<��=;~T;�6�:�m-�8jl;�s�;�~�:�<��\�na=�^���n�<�P=P��lC=��<&�f��ӫ<��<ゼ��<�DJ=+S<�}=����W�i�gɄ:FG��a=Nt��4� � ���<���Evڼ:/�����i�<KL1<9U�<��+�\�P �<�S`=��V=�%��R��<$�6�Z]���6���z�לJ=O-�F�=+pm<#�=#��:W���BF��od=��;*�Z�-K =J~�<ӺO<\x�;4��vF
�ԡ�� �,�b(Q=�k��bI<jS%<�?=o�9="_={=-3@���C���}���C=�(<ON	=[��i�w=!=�ܸ<��[��E�y�;��
<n,R�Sw	���=W�?=U1F�.)l=08���g~��q=X:�ے���6<W�q����a�q=��
=��s��=v��w��r��d��a����Q�H[g��Ul=�%��{P.=�XA=v�
�Q<�&=��V5���޻��<�&�<���<&����A�#�x<��ü(��<�a7��o�<���[�yז=��e;�F<m�=%�ҼP�l=�h�;�F��nd=,*��.�����л
O�;�皼��D=YD=����D���E<��(�=q=^K=���<:R=�=��8�84�U�B=��5�l,8��j����8��<��?=w)�<�{<5�(����\u<��X=�K<#!=l�ҼS�*=��=��n��z=�r�<%P�^���ؼi�Q�w�ļ��A������Y�<�f�<r B=�4�<�0P�-�(�"l<�zS=q>�<�7�X~������2�	üڔR=6+=�d�,�F�Rd��k��r�<�򿼒������n=��@<�vG����c�]=���	V< �=:�M�`�A�d=D���.�7�=�3�o�l�<*#=��}�?HS�O��oO�;
es<��!��; �=MC��|���<("Ҽ�e6�r[������ *�D�n<�9�=Y�_��}L=��=]]���%��P[<����<=V�z��K���V<7A=�}=�U=�'ҼU��:\�<ˠ<�J�<s���(�B$#���<pD�<���;7�<Wle<>C;�m	=+x���%=����
��;��tg�P�"<�S=6���dc�I=��1|;���<�̄�(Y���+?=��:=.�~�v�"��pƼwB����V�M�h;���<�nv=V0@=�}���0=�Z�:w��<���m|���9"=Gc3=w�;=NG=6����t���̼J�<�Λ=�13�5ؼ��k�4��ۼ�Z=>��<���=�닼\~f�~�:T�M:��;�D�;�e<�P�<H<<Fo=yg�<L0����<����xmM�YN����<�w;�0W=~���B,=+Ϝ:]�B���Ӽ'��B������Elj�a0t;`+ٺm�< ��^C=�sx=g�O=1�'<矢��=P2���s=1`��y����c��O�Ҽ+̥<-�G��0R=7��Ì><�ͱ<7��m=�z<W�E�]ڑ�#�%=�+�Q�&=W�I=]��<��I<���<X=���<��ٻ� =�mO�r�������<�%/���{=s|=6�)�("����';��#=i��;�h仔W=�=�Ԩ<ʢ�r�O����d��<X=W���ﶼ���<�:�;K�B=�;<�>=��=h��<>Ǩ��׎<>��>=�p=�G	�z��睗��P|�'j��/%��-���<��f�XB����=�Ƴ�'n����3=>H�<䰱��[�;���';<OM-��r��#�h{���{���,�<'(����M;��=��=vZ�<�T�<�፼�����P+=�w;� ��s����<�v;uW$��.}���`<?��O=p�f��(��*Ҽu�<�B==�Jw=��7��S�鼜6�;�$\<�hg������]�<��>���(=�<��=0�P��X=*r��[&=ޔ6=� �=WS=�a�*ni=��^�#�G=����q}��V���!9�G=��9�������`���	�n�ϼ�[ļ[62=*=�<���*�<t,f�F<�;z߼�2J=�vQ���<�l"��a=C��<�%=C<Ĭ�<��<��*��CƻPU���s=�c_;�e��$�:=��#=
�<WЌ�a�Z=��k�nTy=?#=�2�<��>=C���u��P�=����n�A���<��(�&5=Ĥ���b<snT�Ё�>�񼋆R=ή��	#�;�/�����N9e�5��H�=ds�<-�6��c=��0�2�*=�������4�<��z��V��=��_=��m=A<w�W<������_�X�E~�;c@�<rw:��9=��<�ߥ��H�<�|:=?�a;� =�4�<���`�u�&����뚼�!=��̼A�=m#;k���w��z�-�'���==,���>�-=B�<�b����(����;�<=�9$��{A��d�;I3E=�]L= ���|��O��w='Q��<3�P����<E�V�Ŏ==i =��+=�?=M�<:f�96�=��D�����	�лu:H=�1���Q=�ȼ��;�EE5�'^����6�	�;���x=�����<��;<��-<5������z��Ƃ�<C;��̟D�J٢���<8�mD<�^Z��d��2:������{X=Eg�6����A�N��<˖*�!�����~��b�a=b�駉9�[�<1U����-���<R���<�wX<���<���{)P�B�?3=��%�^��:z��F�ʼ��:�<=��(=�=N�V������<��w��v<f���a;ςW��g�<��p�>�=�l2�<���<I}=��3=���T��<J/�X�<W0=���<e�:���I�w<?=�E��b�
�jT;HF����>�;�HJ�<5i[;b��o�;�����<�=�k[j=�l�;���%=6�j��D�<��@9̞=~=��=���:&:�<��E����ֲN���b����"R��+=��
<P1_<�(p��%��s�<�*;�f�C�]=�<�6�/|�^v�@��g;:<�/x=�e�!?�<�vT�.��<e��<cjN�ٷF��=�����3X;w�P�B�_=�������<���
�����)=˜/�3>N<&m=�'`=�=�	��(�
�6�%�ƩQ=�!0�j���
�%=�n�<Y�<��߼ڑ�</T"=4o伆C9=?He�7r�<k�E��	<-<ּ���{�<�:�;�U���	=���<�~<6u�떼��1��u=U�$�[V<�7��<��޼
PV;NB:���<|))<}=;�=B�&<�,��q�L�<�z�8�xɼ5�+�.���U�#=^�J��:�=�A�<~2�M\�<P�k� f���JD��2��¼�ԓ<���<8T =[=L=S����A=����|� =�|T<�qu<�f�f�μ�켳9M=W�^=^J ��}������Ƽ����<�i(�W�'=@ؼI���k�4��<�� }U���<��K�u� �ŚE����&��P=�$�u=$��;���<!����e=�����P����;gu1=��[:�=��^<�ga�i=��!��B;�|H��R1��<HP:�J�Z�|6P=�'S=Gg�<�G=���;�lg=�4<ā�{�M��T&<i�<3i����<'c9=&�<'� <��a=0kZ��+&=����g
�<J.= �$=��3=z䷻�j���u�W:�;�P����P��{(�%�Ҽ�
�;�p7�j�(V=��<ei�;r�@�p�=H1�<n}<˩.=_=�����gy�T��;�e=pv=�����=�Mt��U=��=5�Q=?+K��iK�9�<�6��(�=���̌�<� c�� ��ޯ=F��<��<e�U����;�Y+�H\��ܐ~��D�\D$�˃���Q�)43����1�(�<M�QR�9hB����;�e/=A|к'׺Ɣ�<��O�P5��GF<�7= +=S�?���u=琪�~��	�d=�(;�2�<� G��w=>�!�Գ7=��;�@[ �3��;�M���=��;I���駼� �;c�!��޺; �=��=J�)=��#=��?���<ÅR�@�{'�<pL�;X�z�։�<`��;p�,;\)�ZF�<7`a����`��<�Q��9e�<�uN=�o�/TY=r>#��	�;;��=��M��eC=��6���+<�*�;kQ������W������.���:�w��2��M�8�#=�y;�;�]���h�Լ���<а~�+��<T���G��H��N;���<#�<j�9�ި���s7=.��_m�:��x���;=��=�i�<b�B=�KT<�ٱ<2`x��>p�2��*s���9=��»��OO=�Rz��9<�P|�z5�f�����ǻ��R��M�F����.=AFb<�d;=�\��ҳ_�2Zi<�M���%=�k�<�B��T�6=�v��P��5�����T<�!�|/���2�<����HټL�#��7<<�9�8vR��;.<E7��Tぼ_�$=g���_m;i�;7X�<t��<L�=%#=�/"=�t=���Lx�:�=��g=��S��n���(��UǼ�l1��<W=ڌ��͆��?���x�f�<��T=��R=��=�v�������<_����	���	��\=S;����׻�O��mk�<�N��w�<������*=��	=����M<����e='�=��j��&�oa����=�D=�0=��9=��$=��8��Fj=�]<�w�<5(�Z-=��׼0�;cC=B�9��3ȼE-� 	I�y�7=/�)c��U���,�<�>=�伮q׼���<\ �<���<�V�<�&�o}I=-
<������b��?=	�w<�<:�F<� ,�'"=���uG�<�cS��o�y�y�p�5�]dm�z���<�����7��G9����K��<�c�2	�;E~=е��_y��N�j;��+=¹��5<0<�&=;�¼	q<"=� =V�E�; ޼� X=�=��b�r����;=F�<���a]�k����x�^=�W�<�����,=�tF;�@<�i�ck#�p�(������ �<(=	��Q��a�F��{<���<d�=�e=�W����6�GZ=�*�<����~?�<7��;�k����9暏��4�<s��<.1=�̜<��o����;�����bR��Ҽ���;���<�r =��Y�v=�٣��F�|�J�<<E�=j*^=9A��k'�SY�;���<;�F=�&׼��=�t#�#�{�u�1���
����;9�<��\�n��<�OD=��;W(�<l<�<�����%��-�S�==ȻW�M=hΨ��,�fߌ;��ż��=;V�`=4b�yg���8��Z�<B��
�=*	J�0�4ﱼs=5���e=+�*=��,��H̼�N=OTH=?\s<����@7��ۻą><ԙ=5
b=T���6_�L�h��<|4z�o�,��!4���N��.���Z��S/=O�M=j�3<yX0���(�%*=�� ;	&=���<yb�$�Ӽ�d#=���ܹT=y9�<[�p��]O<����
=]�!�`�3=6@=��?<�U2�ٟ�<�=a��<s��<Q ��)Σ<m�J=���5��K#R�#X+��<<�%�<u���&�<��.��M;�ק��;<��4:�9�<B"��b<�«�7�-=�Q�<�f�<ח*����<�
w�G� �s�<���޼�I�<{��<ӵ�<�;��?�5o=�	9<]*=�2�=@l�<�3<��H�� =@�x<iLi=�=,=8~4�JN<	�1=��I=�]=,���s1�<N�O�� �<�d?�������<=��=D�=�0s�a
��ӆ�c7[����%<U4�<1:�L�Ի�e�Y���=��O�c�2�{0=1��;.�;޾�<�R�;�>�<�j�<w��<%T���NY�t��;zp�ci,�&d��Z�<'Kl��mA=O�3�����xQ��x7�xE�� �<.�V=��<>&�;2p�<�m�,z>=�L��v\�'��<Sf�*0��!"���,[=���<�?�<T�"�C��<��[8M��x�c=*4)���ټh��<�og;��&=چ�*�=?�=�a=�����T�<	�.<�7�T==;k=�^W��Sռ^�h<�K`��� =�<Y=��e�g�H�Rv=��L���<�8����ټ��ƻ���Ix<�2�9č���=����>=n��[�<��=T�_;,n=���;�SF�e�=�v�<.�;
�	�'@�����J��1���D������D^�тl��t<�Tw;LL�v+P<���<�DW:��H��b�Z9�;��U<nܙ<����;�K�09;����h���wjq=�>��#0�h>�<�=�UF��l�����S�)9=�Y=����Q1_=$��;�z��¹=�4��
r=�$�(-��G�m<b4v��F<'<��M�ǌ���FE<����"��a=#1o�6�T��	м��c=�Xl��d_�b��[=���<�W�����}=��μ������@=.c˼>l=^c<`��jA��e�<��K���\=@8<��s%��� �������ػ�1�|�@���Y��o=�r=�h�<v�=8{M��K���Ǩ�s{�`=�;AD==l��L�D=�����NU�_���/�;�H9�h8�`́<�Ѽ�S���T���=Γ)��)	=���җ���r=x���G�?%I��VU=X"V���{=q,����G=����1�x��Q<'�=<�p=������=������<���!�+�9��=�C
=z�<nò<W��<%3�H0����w�n�����ԻM���=8b.=Х�=�'=� �ymW=s����2򼓥���)=��p��<��>�0=��N<� �A�]�6=��t��R�<,D�:s=s��դ���<9;��Z<$�:=ZX1�,��<��7<	��<G���O_�>��<��?=�B�<"E��K�������8=V��iq='2(=yYa=��<��7<�s��^q6<��׼	TN<�v<�tUl��}ļ��<�|m<G^n�Hq��G�=ǒ켍�=��:=~�|<��e=wK���ʼ��P�G2u�:�ܻ� =��ڼ�]=uq�<z(<� ;�<�<-Վ;��;��x;=��!=�(�;[�=��<���yp�<B�=�켺{���U4��W�<�L)=�F
=L�<��������.{�<���P,%����,�<��]��z�<+z���1d=|B=�:����y��<ي=��=�q4=���<��?<n��T�<��<툸����:`h==ր�<)�%��	�=�_�jiR=�#k=|ͻ��/����D=d�+��U?=�:e��=
�<�Ģ<Eb��+Ӆ<�|7=J���u �5İ<���<�[�<�l��t؆<H�?�C�<�R�<��¼�G�������S7=Ζ-<��=�KE<ۇf<��<���C��k<�'2=H�.=���<�ڞ<�I�����t���L7��k/��o$=�f��.=����]=��;��B=2��;Z>�(CQ�����8��;�O�<���_�g��@=.fK:��	=��Y=��:�W<�b=e腼P~@��.����;��e�Sn9�*���`<R���5� �V��;�{5�<E�:=���<�(4=S��<���f�j�-�C=�zû��=��<�ak<��=��ϻ\*=���)=��
=P!%<
���~*��=A�%;a=5a=��M��`=#*0�Э<禼����Y=۬�Z69�`?I�������<]<x<K%3��$:���]��,��y:�ۋ�;�+2=���G<�p��_�<�'1=`���X=��<�����<M	;�n�`zټ�b���k=�=���͔�<�M�<�&��ܻ}`)=E�2�86���9�<ի輦;=������<���<�rG=�b��J'�<�ĺʰ�<�X�<�S=ƚ�IǺ[=D�%Lo;6-u=Ct�<&�/<s�4�֐�3�򼼼����A��\�<�5=�8�;��=Z��uSO=��W����e��<Y-=Ѿ��x9�<��+��0}���=+�P=�V��)/�?��]���t<�7;=/հ�5~q=�[T��U<yݼ��ü{�m=�Mf=��;Mr�<˱�<@(`=Z�Y=(&��$�;����T=@�,=�(�{&<4�B�?1߼F^y;��=���<#�$��7���\�Ck\=�f����<��)=t�&|<��ɼo��<JXj<pMU�X��<��;��b�����ҍ�<��5�.���T$;���h���d=Q+�<m�[=�<��<��<�)껷���F�G���_��v!=�Y#��c=V{/�Ѡ���û�5�<�*�l�ջ�Aú�@=G�8�&=3�<�R���@�<|��pKM����;��<�ļ���<�#�<�?=��<��2<�LH=1B���<�s=��T=�����%���p=�Aռ�亭��<�I��T	��c=�}���O�<����o��I!=�J=�4���++��z=�+m;��S�{���b/==�X�!K���#<	k�:)؞<{�&�o�;���1=�w=�6�<PAU=��v�_D=�8c�y�f��/%=QP�=E�<� �*4�1J��=|�弆�=7&�<-�]=���7:Q=D��@'�)-L=I�ؼoqt����<�G9��=���:&֖<[�M=�)�� W<1����w<X�~0=s=m=ԇ�<�hN������(=���;�ؿ;�ļ����OD<�\�<D邼tA8= �:=}-2=-�=*�{�6Q�<��Q�}*=]R8=��g���^=�c����k=\Q�k%G=�?R�-�<e�	��~��a+=o��͑�;�Y��Z^��$�<�<��<sj_<f�V=��>=�C~<��=H<=�ּ�<�*=#5���S=�p=�#�<�fK=X]f=�S<a�C��8�35�:Q���6,s<�<=_$�;E�;���;��=�_�<��}���'=�2?��[�3�<��=y��<�.���J<a��zd=��=�W=�1��S�<Ϩ�<�u�l��<X�S=��B�Ἷ0	�W��<�R�<|w=��Q= �a=�м��<�B�xDO<&���]����'���I=�\�A=����&���&v*���<{j����k*g=�v��K=}6=��/=Q�n�<<2�A���0
��$�<( ����u�+���<!�(�c�<�AG��tp�`1G=��<^+f<`�<�Լ��@�L]=!q==�y�c�D��E=��<����0�<W�d?C���<p��Ic5��pc=[�=+0=P?�;Q9_��O��}\�>=���<����K+=���<a�<�?=�<����<�ݼ�Tn=�gM�&�:��ϼ���<+��ћ<�>/=�>H=9�ѼU�U��]���|����0=�<��<�߱�R�<�QR�*��;>ȼ��#���R<��T<�X�;B9\�"|ѻ֌"��x�<P������<�L�NU�<�ɍ<�)H<��@<g�<4-����;�u=4����<���<��>���"��7��CF��C����<����r�����:-�xF��*A=���_�H=aC�p�=��އ=Yy�`^�|$ܼ�S�;ӐU�׵�gۍ;d�=ƪټlIZ=Gׯ<�0�=����=+��6�y<����"j;�tY=m�^��Y=�<�}V=1�7�Dݼb�ۼ6�����ռ �<��$��Q̼͆i��Y>���=��r���w=�^�<D�eN�<A�<������&����}��<DWI�^Jh;��&�.����=��O=-�I=��^��-N������X���+=��<gV��fb���Z<'Z.�� �R�|�Բ��3x�vm�$��e��;��e=p� ��
[=S�������5=�<=m;���`�⬻j�W==�>��xh��K=�=(sy�9�ɼƨ(��z�<�Z�k���{���%f�Vݻ��m9����5˻�u+=@�2=�-���;fq�<��<F�)��b<���z�<<�<�����[�<˟̻Lt[���;8����=y&��%"= 	�*G�=Y���;��i<��V�9BF�=F�;hֈ<v�*=D�;R5o��IU=�S�s����<͇<=`�=�]E;jv��~�<³�Rk/:�f(=� �<D[��L���Ǽ��:�{ֺ|�8=i#��N�v=� 0�N֟<[�;��|�g�.�g��V�;�P,=�^�:�&���G�]���Z��J�o���>=ހ޼v����~<��<�]M%=�T�<E�3=�t�<8�y<��<�8]=4�n�*�Q=wʝ�c��o�>:���A<kZ���b;<�[��=\�ڼ��<RI�j�%=�fX=�b���X=旣9F��<�!H;��I��A�<��~��1ҼSܼ>O��"��ݝH���"=�l����x�`K='(K<�!;����5�&<�n��	 =��5���߼^����Y=�_�<IB ���<�g�;�g��KҼ�cg���.=�꼻�T=��|=SQ	=�V5=!�4��н<_�l<[=n��k�Q���!�{j̼��K=��/<OEd�� ¼�L��t�m���=�"��t�����<��;��ͻ̣<.s�Z
}=�?�<��D�Y��< �<�>^�@�<gͳ:�AS<���<қ�;
'%�9��=�z4=]/���jZ<����P�����B�ƻ8~�����f<%3=/W���`5��w��{�=�H]�8�߹�t=��&=�T�<t��<n=l���"=F!; �`�ti�V-]<
���>6�<��s;��*<����=�T=��5�@=��ۻ�/3=.>R<J_4<r-�OG;<;
=<Q�;�<o'���;�jN=d�[=��!�v�⻫����2�S���&�=U5G�\�\= �-�xeE�i�<�4<n��<(V:=�һ�	=3={�n���z��2�;���<l��</F�v�t���Q��J�P�o<P�4�t!����<�C�<��=5��<�J�<�Z�<���r��<���<E)�7��)Q�;�u��@bt����"���<Sz@���x�!^$�7�H=���;&4<<)�<��(�ۺ���?=�}L�{x9��o��E�=ም<ͷ!=��"<�Y<G`ԼU�w�3`���lB=�IG�}@&<#�ۺ\����=��F�lZ��:K�BDO�i��;��|��<ΘV=���<]fͻT�-<S�޼q�&=��,�P��<�e�;FU���J=|�.�0�<R���ļ.��v<|>=��<,�M��z�<N6�>�	;+MV��`3�<���� ���꼁�(��׌<�q���h�s�d���5=3��R<��U<~��<��8Ŏ����=�<�#T���F=�:���=z�<�!M=��;|3�<�Q���g<��-=�#��#f=�?H=�� ��؟�2�<͋D�j�ؼb8���ڂ=���՞<7^
:4�B�o^�<.,��g�殜<���<)'�Fsi�X�ؼ�쯼�?-<~4>�Q����2:=���,5x��
�ݬ����T<iΠ<�[���>���3<=�;<���a�:��M�z=�;��C=`j���w=_ԧ��ݼ�/��q�<�aV=~e��,&��Ϻ�H�A��F?�v�0��:<lg=�=�^��H�<�Ҥ����64p=��<YR�lCټ��x��W�7A.��&��Q�=@d�_�<���y�\{C���_<��l�r��;�a�����!�[a"=������<�̬;�zO=���#���C*����<��,=�3S���&<+ �:�=�CE����<ݑ�<�tC�5:==$8��M:<q
ɼ��8�~z=-K=��<���,M�;��<���򍊼)���X���F��@S�'	����<��J�rp;[�(� �L=6�3���ּ�Hk�9�u��8��n�G���S������Z=�d|;�Ȉ� 3�<�v�<�!=��=��� R=��3<� =�'C=�����[߼u�;= �w@�S|���<B�:�i1=��<feT��%��p�;����BS=¸&��d��F]u=ۍ�s/�����\,I= �C���z�'=�e<����^�Լ��5�p�W��n��\e=i0&��(�<gX'���d=E<k<!����I��Ɏ���'=�o<���<����qz���J7��g����<S4�:��A�
=��}�8�q� ��1S�6ͪ������B=.G���d��2��!�6���4�<�Z��"=_;\��<������ɼ�x<��1=�=���<Tn���7�s����6��n�<�Z �ˮa=L�%=�;�`.\==���Te<kz��F-��Na���=���<t�3<�#޻�m;��d�;{�#<܆`���"��:�i��ʼ��3<�^��P
=u�@�os=b$�$⩼MQ.=�����Ȟ8��j��T<c��<�������%����<�#�T"�B"�s�<�e�0=x[żu���g#=��"�B��[�	��슽�Y[=�;<�!���E;5<��'=n8*�,%u��㓼��.=j��;K���K^=�uD=N�4�;TY�����Z�A=��#<�@.�$��<G;�|@�{_=�֡<����m�$�%JA�@r�[8R=5��7�`=�y�<Wh=#hT=$��='��<���<&.���cE�<�x=J(u���^�]�2���	����<��Q�y
 ���,=��[��ݒ;\!�<�Ԩ�*<QBu<<k�'�<�~$;�@=J��=nW9;r�<4�!=yqe��`=�q�<���	:hO=�j���P����<�y"�
p¼U1<�|4=�:�=^����<L��g-���k<9P�U�-�*}:����<�)��Û<�����b	=�\=�,�ٻ` <� �<��޼���}�<����^Y�h��*�=��3;mR��/�B�t�u<�,�q��:�e�;J:ݼ����k(�N�f<�!t;O��<5������<!�`=���<��2�{?p�ދ<{㼅�p=h��<�Y=��	=�9E=��׼��{��<-UY�K�=�Θ<�^����=����s=��`Y�:�\�n;`=�vx�;T��_K<��wK�b)=p`�<���<-��f�<k��9�\�<i�J��ZJ=�e;��=��=�v��Bռd��<!j(��[�;���<~�h��ʌ<\�ʼ�oH��%=nk��U���>I=���;�#���QP=��6=f�=$��n��ͻ.�Z=���<{E��;�;���r�F=�EP��N�<]n;��=�2���C�2^���a=p��<^!$�YX�<O�߻���킟�J?��r�B=y�<ֶd=^�˼�ӥ<ö8=�t�<O��<r^1=!�a<��#��E!��,�{�<�hA=hM4�I8�=^�P�;uJ=ll0���<Yu�<O旽GSɼd�~=�j�e��;Ƃ =�I����\�r-�<��<a�׼�BO=�I�tO��� =�{;�����#=���;�v��uj��������<U9^�=�v��9��"���"�B�;�}\=
�R��m&=l�v=��=a4)=�pݼ�h�AxB=��<�[g��Co������[=�E�<�,�uBX=���f�==9�<$�=��|<D"c=�N<��ۙ<�*M=v��O�=S=bd��NL=W`=v4�<�u�;h0~;���<��9=��=M0=�m4=t�B=S�� R=F_H<$���j=<�gK��<�J<��Ѽ ߺ&s=Rs=�/�;%vA�*:��j�輠�6=��ú��>�wa�<!S��?��n =ɺ>���[<�1=�����~�<ڀ/=&J��|����}:�ۀ�&z��R=Z}��X,��T�R~L�����(��I]���;=��)��N=BQ=�xۼ�B��͵�w
�<�bʼ���#<�;�: &(��K=֧�<z����α����h�l��7����<�?�;m�<<�<Eo!��0&<};�	�<��"=g���E*�S n=߿��Hܻ3��<սF=�
�տ:�$;[��;3Rw<L'��"�<� Y��S���W�9?=B{)<��C��;�#�3�X�����<��V�	�!6=�.b����ڙ2=<�oY=�������̼;�������U=e=Ǽ�A���=5�b�8=��Ⱥ*�I'���@=ip�҈&�_(�<��<��%=�3T=ギ<��}=�]<z E=�W�2�[=? �����<l�k��=��7=L^ݼ��=(i��"=�9��!cd�N��<��%�wȉ;To���j~<�C����w�����Id��"��"���E�Ƃ'���z���=�_��?�v;t՝��;q���9��r���w;���g>�$�:�v�<�m���%=u�L=�G��Y<�X�6��<���HS=c�����4�N�	�N2�;*�|=�ɟ��m5=
�%�� %��H�g6��#i���H���l���=|����w=��`���T��5:�4����X��N=�Ȭ;!�?���ڼ�񥼆jg�T����vP=��a��m=���:�J<��5Y=2��dV�9>m���:����'<��=�(:�u�<9:2=L7��*�;��y1=/,n<��(��*=m]T<�mS�A�F�z�=�+����<���0�a��B=/�n�ۗT=�<xy��}4��r��<�) =��<t|P�ŀ6��)����z�r<3G;�~si=�3���L��P!��F��\�<z=(	P��ǩ9��8=AU$��y<��@̻����n5=D˼�@�T��5���v�H�{�=8s�<@]P=���<�턽
յ�m��t���ո��,<��<arq=�w���-�%��<�zؼ������חb<�<6~<�5=�䛼&|}�8|�<�鯻 ��:���;����м��Z� �<!�<��=�PY�B�����;A>��G<�&\=�f=,�ҼIu��֗D���6=�>=V�6��6��r(��?&V=,'�ug+=RbU<�$<�9�;�2�X;=O�6=��-;&�<-(ɼ�{��OK����<��<��&�9�;:����蜻}SS��3�<	=r&B��V�<���#l�r��;K�W="�W��D �� �7䍼�1�<7�.w|��.ż� �<���[�C9%���޼!��<Dm=�2o='�v��5�£~<��wo�;&����|<P��Li����ԋ;M��<� ,=o�}����<(BμY>J=��<��G��bt�sJz<`[S=��;�3E=C�=��9U=�F.=��e=WQ���Y*�MW��zB�<�p��Խ����$'=P޼�H�_۞�e�5��<
<�<���?�I=bkG=�0-���<%·�?�<�t�����-$<Vt�ZN��Pv���<�=|oV=�K=��2�}�#=��S=��=d*ۼ�a�<$1��qa�Q�����<q,,�0eۼ$&>=6#9=�B�<��<sjF;�q���'Y��\=v��?��3A��vL���X;���727���<�Y��{�w)(=B\O�>����n�	)��P�-� ���1P!�g�u�H�=�̀�j�&=�li=Zq<�<����K=�|��`�<y?=�ء<�9ټ�m+�N;����;�2�<��"�=��j�=0=ƿk���;O�<�mG=8����;'f�<���O����;=ɡ3<��|�������X�����uv�1$!�v���/Q�����;��'=s��<�v�;� �<B��<1n�7����o�:��7��ha�c+&����<r�U��J=��a�����e��M���⍼бƼ��J��O=k���I=��ǻ��s=�ϻ�Ѵ<F�;��<�'=� �<��B���Ļ�K������;�G�=��y��Yr����߹/
�<�(��hy=�n=���c=�(�:=5=�5$�_7�I���o�� ��:��C=I|w���8<�D��Q���m��������;�A�C&\�����{R��߿<�DC=7�Z�Өʼ�.��Q�Z�0=�0�<~g=��C���S�%��8���>��O&�<��^<y����R=c�:3 b=�"=��<�(��@<�9=t}<�wG�A����f�<�[��È;���<�<�:=D����P�5qA=���<��m�wD���;�=���A��<�M�a��������_�.�L׫�y�!��V=��$=�|==���B��;1\S��7y<$p4��i��
�N��iL��[=��=6����_�"�=��=^���5=��[�s�%=rJ��<~����*=m�<=�S��!�'��t^�i�=qo��o�5�KO�<���Q䢼
�=�x_�	��<?61�n�r=�x�<��	<�W-�,��sV��4�S�N=��?=�<>���Ƽ,d�:��$= ��O2��7�L�����;�{�<2IZ��f�;�Mܼ�U=��i�|����UE=0w�<&�=P��s�;��.���=�]=�F��v ���d�c(T=;�n=2m[��8/<�I���n�<��<7v��f�=��c��'[=蔓�h>�&_���<�<���]=�����<dJ�<̻���<�"=�c=�.���6�J}�;Uns<j��<Xa�<ҟ0�w桼�9.����"E`� �i�pW��������Y�{v�!�^�b)]=�r��$�<*/Q=�( =�ށ��n�Y��
ɝ<�	�"b<��WQ��MмM��<���<�0I�_��\_
�d�p��`�;l���V=�Qu���;mT�<�V =��$���fܽ<>��;���<�2=�`�dl��k��	�g[=��ּ㚚:��Z=�A���^<��G=��v�4���l�<:�#���;]=1� =s�ɼ)����<��s=��]��$�;UĞ<v�=O�P=o�
��Ӽ�OV=L#��3扽b�C�<:R�\8�Q��<�;;�AX�cY�����=�1�< jU�����<�<�\_��}4�#=7=q�X;��<�y��z�������ؼ�^�}T0���Ӽ�k�<�[ ��4=�~L=�M���갻$��,�>4)�o$&;p��D�ɼ<dV=:�]�m˼\�ֻ.�/<�W�:L	I=&�R=\v��F���^Q���A<��=�6�<s�=��H�S�Z��z��; ��aL:���(=;#J=יi��'=�)�<��N<�/w=\R�;�}/���"=�,�<J�R��z*<on=-�;,���ő�;��G�PIq���:5��=��<�`\=��P�]=F �:U<�*>�<�<u=Qb=.*i=��Y�K�0�sۯ�D�9��}=��F=�G��F�R<i	=��I����<O�=h��:q:������ټ��_=t�\=��Ӽ]�*�'�I|3=P�;�Ǜr=��>�L�㻌j׼�CN=���<�;H�eĽ��".��x=����<���<N��+_��,�j ��-�"==+�<��1< u�<��Ѽ�t���b=ʔS<�u������
O=���+=P<;��<2�k�U���p=�:�9�.�[�󻻪�����<�;X���z���<΋=�<�<=��=�Z�����w�=}�=��e=d]��<m�Y=./==G�¼1=K*���p��+<=8�<�u�;t����+G�(�ZL=* =`�<��
=�X���;.��@�&=.��<k��ώ��;U=�;P�#=�pc�.gU�5�;�ȇ� �=K=�_�������;�Q��Ϗ�e��;�MR��3�:��<�}==lz<B>��~N=z��C�V=��B=�wu�l{c��_A=E�?=Ǥ�<�J�<D�_;��<Հ=U=p�q���!<���<1= *@=5~=W�4��+�; 2k��g�<���@�(��u8=�R}=4м��H��=4��x/=t��<uZ=ͳ�<�W�;y ����a v=з�<cʨ;ӡ��������<�O8=$�����c�މ*<T�t�2q�<�m=���<�_��l��:"껣)��͚<�+N���*<h�v�S❼/?/;
���tW��7Q���	���>-:<MJG��
.<[�>��2=�*��������Z=��B��Z	��l<)���Έ7�d+B�j�0�㷂�lp��"=���<㑢�:h�ǫ8��g==P9=~ڻ�Q
�����A{�FS�_!�<��4=Q�6����m`�KS=<)��;6K"<�'+�b9=\k�� n���<�=(>�/���l<]@E���<�߀<��R���!;�X��`7=/=�<^( =���HE=�<;�{~�%@<��u��=�<�{�<�q��k|��h.$=܀J��{=$)�:	�����;Nf<%G>��Pt<vL}=���<̄T��r=<�<���<Q����<Y��<z�b=��8��AR=�J�q?�<�<<�'���<��=e�#=�!=�@߻)z<�N�
�<2~�2���
Q��_<goi��/l����<��F=�i��;���=�MK=�*3�B�<�ܿ���<钼�����{M=�!G��(�<�<��<�\�<�7F��
<��ۻ�p=M��(��<��u=�+<�"K�<!��<F�YG��kȼ(�� �;U����`=�d�<�/=�jc;�c<ϋ_=���m��pM@<���<<tg�ń
�B�=�N�<�Z=�����&=��<�^z��n=��1�1r��;��\%r�%�%�U��;3�����U����{l�<�[�=���6<L�R�N� �������_�_��\�<���;b-"=;�=��u����!�ü��{=��2e=I�<�z.�z��;6j��-��V^�<7+�<>M+=��»��,�Z�e�����լ1���b�l�*=NVt��r��;�<�d¼�*�ifu��{b�6�=�b<O��'=���<`
�9�1�<\�9�ٲ2=&��:sѡ��I=X{��/#\=w ��S�8����,��L��ZH��h=�=ЍV=��T��:�'�<4y4;�q�<o�5=��U=`����;(��<}�����@=�]=�z=�洼��"���-��8_<n# =����� �\�<��%�yl��"B���]���s���ۼ,�S=��k_=�r^<m�;	��߅�<h�;����u*=\�<���<R籼����� <���I/�#�Z<4B;�Oj����<C>=n`�<��F=4
�<ߜ���9;
����_T=-V=���<�f�6�V�����o�=��7����)%�����_�;nbܼ���1�8��q=� =g�;+bA=J�mO; Z�:}^���#=��;��8T;v�o=�sK=�N=�0=l�!���+=RF�<"z�=�E�<FJ���J<#_)�a�q��w;WŻ<�e���<��|����	a8<y�����t��Z=��)=V�&<���=�>T;�[I��_`���=OW<�*b=�i=)�h=rH?���9=Q��<3�l<�Yw=�&= �%���<M(`��J=�{�<'�<Oȕ=�'<y	��ח�m8s<��?=��<f��<R=i��;]�E���<���<�yԼw6�Rֺ���<�B=0�=\ko=�,=���<����Vi��FN��hX=�E\=.=�+���=��:~;b;���H�83G=�(��I�=#���kx1�l�=o=���;٤G=�*�<��q���>���=q'�<�pe����,eG=�-c<0}=��~:�k)=���<����XѺ�)=�g�<���U��=_���?bH��G=� =����+R��\����C=��P�RD&��m?=;���&�"�Ⱦ�<�봼�e�<�|!�������<Y2Q�t�9����<��m=�����ǻ ��:@� �B���\���3�Y<�2��8�)=(�<�)J�yt?��b=��K�􎔻��=�lZ=��;<is:=�A=��k=}c���#=�U='q<��#�2t�`x7<=:��MW�>�޼?�<4s�<��H��vT=�6i�FS=讠<�&=�[W�j��a�<�a=�!��{�_={e%��A�:�h���/��v�?����4��ST<��X=<ς=�܁=pil�2���&=T>,=p�g<F21�~su<(�M=�h<�'=ˤ�m���\=:�:�s���n$;�(�w,=���.�泤:���;�<}��;`��	�;=N�$��強�#=��;�ھ</�F<ʦW���ш=ؖi���	=u7�<Q�T�jE���z<;�ּ���<x�&�R��=ӝ�<���)��"<=5~�<���;�Q�����=�� ;D� =��=s��<�VM�֒��4B=�䉼��o�����Ă<�N�3�F<�q��>��]���c�<�-=�ж<`5B=d�/=�?��������� �p�=|���8�ۼA��C��<�yU�ϳ;���'<� ='������û@� =TY =�<�5g=3-�c� =��D=!���]'�%��<�b=��.=�r�{T:�c&�$&�;/Ǭ��K=���nޕ�T���/���Ҷ<Z�Q�N�t��d|�=�W��2]�ߴ5�A��<0��?ؼ3��<S2�<����5;=���<}��<e\D��wv� �<��<i�=0�����"�=zP����;��<4�<�iq=k�.=�}N==p'��E,���b=�\�<� �<��u=!=�>=� �}��<Z�r�N.4��qT=cG��˦d� ��< h�<;�ʻH��;1�=�(�=f�@��Wl<��Ȼ����d����-�=��\i=3�>=��v=���Gc<0��;?�=��y=�r<�2�gJ�<�}�=Qv�0�!�u�=�d�;}wԼ
`�jY<��=~3K=v�o��	H=1�=U%��;sL��,�=(�<�Y(=&�м��%=���������W	<O=�Y=_��Ͱ�ؤ�<QL�<�
�b; ���;��'��ea��D`��<q��2;<��bn��W,�<{��;�z&��V=�M=�����E=��<r�=J�L=�"=aoԼ:B=�J~=��
���<0�=�ͼ!����传K޼	��<8� <Ϋ>�J�=��(=�T9=���y�<;�S=}��9�Ԍ<n�+��b���xu;�&��B=���5��NR�g��2����S=�l��KU�<o�|���=A���K�<���Y��6JʻGF<;dL�<S<��=i�Y=��� X���q'=���<�X:<#�=��I����<�PQ=��c=�;1���,�6��<���<0S=�+=�ܦ�LHa=�9=��=�Y7��Z�\9K���I�'߃={���H���.���;��&=C����B�o��:8.��<gaI��O�<k�=���;���< x<gR�ޙ�;���;�=�i��}��V=4'����"��q�<m3-��� =q�,=l=�&�<��Q��A��F��e�k�B4=��L�n��ڧѺ�����N�<Xz�#� �}���q��S�y�Q��;�*w����<�.��|��=ɼ�<�J�=%{���?U=��<�/ּCJ:��!=R"���R��y�=8KB�ZV=�v�<��%;Wd=5s=��a=57(�p)K��V�:&B;�ٶ�<���<��޼��"=�;<kZ==�V���E���<8$=�W�Ѣ*=�J���0�U6�<����׷n<oR;��I=�@=l�=�@<b� �"=��i�	HG��:���@�!;h<(z+;+�+��v，�����<!��G�G��=y�=�2���3�sP=ď����<�+=�W�O�<����N�����<��=��<=�_+�׬��8�¼�Լ��;�G�4�,��qO����;���i�<��?��9K<*~B=	�Ļ���;�ؼ8��Ĺ���2=G�e������K��X=�/��};�<[D�<�ܷ;�b�<��v�R�O��?� �*<Ҭ��BR��0=m�=^<I"�<�E+����<��(�<�/<P�=-}=����ż�{�����}�D�N�R@�p�=%\R���#=8>���]����_�;�ɺ9\Y<J=�/=׵\�$��E��������f�=蒐<nA<�E��<�#M=)[��\=�j��B�<����g�Լ0��<�;
�&<��-���h��<'�w��ׅ��L=�PI�1=�����A�<���<�խ<��<@E���n+=�Ӿ�F�ʼz%]=��<H	�v�X��>�<Hl�,>=dS;s�sP<>r0�<�<sQV�.4=�f.�s%=��S<	�=�z�<�g="(P��(=�L�;��Z�^;��k���� =#&ܺz���3˓�'���F�=R+�;#=#�&����a���_���K;���E0�<d�=�/=��H��i��c_=n�<��<�d�5mi=S4�"1�<��=w�/;�����%=V�꼯EQ���]��,,�,�8=K��\�R��ǀ�^�k�����;�=�x�<������p<��>=&\�<b�nY�R�<TH=F�<G�F��C:��»9��<�`��1l;@�+�F=�i�<�wi��e'=?	>��]���<j`�O�<�ٙ��� <��=Q��<9i=������"�k�=����O�H���8��B:=�l���h;B��<��ļPC);��:=����{ջ�-�<�'4�]M�|]�<+P=�����T�*%�;9�(=_�S=by<ʦ5=.�ҼJ#=�W=�I+=�Z=j���슼n�5=��=o��;H�=$����=QK����i�X=;�$=D��� r�f=�"�w=/���<�=?;��@��;u�<�����Z=��T�\��Z���/'=���;�8����/:<q�:Q@����?$<�J=q���~/��u����*};8�=�U�O:�<յ6=�ُ�8َ<�t<XW�J�7=���<W �<�ͺk�<��=|�F=��]�EL]�">=X�b�10�Ȯ���<��q=r&=�ώ<��H=pv� H'=�:Z�0=���<�^��{�d���w<1��Zb���<_���>�vRR�
�\=�E@�L���x�����M+���N���$;�i1=��C�
0j=h.��v@�ԡ��~=�~�<��(���2=kd=�
A��;D�7�8�&=��=�#'=��弬��l��<���<������'�Y=�i�cc���==�b;ȭu=��ܻ@��<�R^�LO=B*�Ἀ<:�6<t=��\�8)=���_B�<;�Ƽg�K=�I;=��;��,=f��pi]<$z9<\�ּ�5=$I�< ��<���b%8�ҖH���w����O�BŃ��`-��.�6Y�<�4ồ�켺��<���:���E�<6=�8=�=�;�%M:�@6C=���<��S��쒻q.H�&,˻q�<�l;�y�>�Dq>���H=ٴ�<��=����Y�L��
�<��=U�<Uo;���Ѻ�]-=�<e=����^�=\h�<+p�<�eQ�F2	=OT��ˤ�AY<Ё:��`{g��Q0�耚<�o=�|��% ���=z�<�Ż[�g� ��v���P�㼃��8�Ѽiug�)�!��ea�aIz��0�=*�<�%�;.�ּ��=}���g�'=��B��a���&,=Ȕ����<|��<���;^@7=UIr<�;��?�7񚼆2�@'?�O�R�_4��N�;��`��f녻�9=׼���H=�"'=�,T;7Q����<��n<BX ��t\=(#j�Z��<ݢ���wB<]�*=⻼y�ۻ-��;>P=m��Pl��)p=�)e��G���:��ب<�?��~�(^{<�e�<:5�::=/��;����ܖ�R��<�̼�$B��0:ʟO=���<:'L=��;=֋��Uִ�#�ʻ�ʽ<�g�6N��!�<�꼥��<a�Y��.�<՛=�=��={�2<�X�gV�;8c:=�����2��7�����J�ǁ���R=�VU���<S�s�u��<� ���<V\� %�<�{��a����<�@�H����< jz�ǁ\��qμ ���K�<z��Z�-<J����<=��<(=���=1v_�'�<zng=j���i�;��ݼ���=�==�qD=���<�,D=�Y=\$5=k䰻��N�W|��bУ�u�L�����p��,�E�D��<��9=i�����S=�"<��
<��+=ҩ;�J�=�6�;Gn+=%���z̕���#���M��*=p/s�'�\=<�`�=h��;zc�<͓��%=�Z=�C/�gA�	<�ͼ;�y������;�yǺ_�]�(GU=�6d�W�k��=��? =X֬:��7{��������/<g���5�:<���Xлy�DH�;S1�<?�7�BD�����\��<�>=H�-�����Ar�<M =u#!���=e0<��`=�G;YK2=��ּ�=�?� T;Fg���_=��u<ոJ�5�`=$zD�E���s�X?�z��<�&;�L��>�;=��3�~�E�N^=�1�!0��t{�DO>=�tF�/���mY�J�"��K	����L.�<=�D���n�5<�|=߻Zn��@��w����<�q4��,�1����x<<4H=�=�n=ٞ�Т�μ"/=��=�x�
����󼮥6�O<}�;�1=�2�; ٥<�L� �5��Ƽm���U=xv��)�m�>�zq=��F���ahb<0i?�&�3<�0���Z�<�9A=�`_==����<% ��<��<�=s���^�Gf=��y=%q?��05����;sM;lkx��&K���1=+"�;M戼���<.�^�$�LP.���D=��,=���E�E=�����S����<o�|�j<<�i�)�<5�@�7k='ۼ�g��6=*7<��=��m=>�0=J<!�$�s�=2�y�S"=���9�6=λ8�����~$����<�,#=�"H���<DO���}�=W=�=f�;<��B=;a���4ZR��b=kA�<	��<�"�<��d=�B�����E��� �U�_�-P/��h4�Χ<��K��Kʊ��c-=bV��/��*ȼ�	+<�+�<Nba=��ûRm*9r�=�8=��;p�:�f[=��S=-��;(D���w�<��<^;�;����,vH�$���R.���W� `#<<~u<R�4����{�(=���:�Z&=~`=5=>�*��C˼ޝ=��<F�*�Aπ=˸u�TO�^�<��C<5z:<�<=%��<�F�;�������<v$2�~����&l��	��"%=[s+��q�9&�Q���yQ�5EP<pÔ;��~�&%�� K��o�<��4��=�=��;�H��V�]7=�=;�<����q���Q�%M	=y�-�~�'��c�)� ��?��S=<����s=�.)��c;��ӛ�������%=���n�<����wH�F�J��;n<m0���>���;E����J[¼�
�m�=я#=�h�<��i��;m�M�d9�6�Ay�L+��,�ڼ�Ԍ=��S�9;@=T�¼^���R���:i3�<0����Q��b4=�/�d�=�����<#�=3�4�^�7=����E��Ka=ɟ��P�;A!�tѼ0��<�B�ny�����<��<���<s�j=�kE=�8���I�P��<$S�<�f��''=�Yn�q�<os';�+=D�#=o�
��|ܻb43�����9I�Q2�J~��|�<����<��%���9�.=��4��`=ڱ<)��<���e̼<�/�<�&=��}�	��H�;���F�K�#<�=��=�4=Z��*J��)�Py=��d�܅6�Z��;F1����L�_���켜�^�T(%�AxO�����>��p<��v�X=�N�����6������=p1����;1/_��N�<).¼����m�=�˅�<�[�۳<�d���-�<�z=����Fo�W%
��qV=��.�Tz@�p�<J�<�pT=c��<Ua=ϽX=++=���<�[�ͷ�`�8�⤇��L=�U1=5�����C=�c�Q{�<��;�ii9Y�<DL��/�����	=v>�< 2м<e�C�;�"�F=�K�<脤<:�=��x���=u�����<��������=��<��a<�=�!�=�65�a\@<�?���h<)p=Ie=��-=X�R=�|=3��*f����<i�����)=�� &�A�<�aZ<�j�;:{t��<m5�</�;�+���q�Y1=\
�kcG�MN=�B�9wռ,*4����=/� Q=�� ��N�<�����<}<\f<h�˻y=6�<@�k=��ȼ�������%=p��;��o<x=����8�<�@;=��<?��<��iD��/�<"C����<B�<�;k����<�v���E4=��a�;������ҥ�fg�;��`�@����f�c���<=�k�����<����Bfd<��"=W��<1!= u8���I<�#F�������<�<=C�+='q?;6'i��<<��[M�<��#���)=�N+�n��γ7=�B����<,��n��nxF�u<9�8��<�_��]�9~�/p<��u��<�s =7ֱ<`\3<\��ݫ{=�Լ���9d����ֻ��J���_��P<��F�B�B=XT='KK<h�;�c4��zC=��9$�|�ׁ���:�9��ȼ\4/=a�8��<��M��9{<�7�Fc.�p����Ӎ=�<ɻF=��r�y7�y�<��Q=�u`=v�n�ir�;U��<ڣ)�f =���� �lN���m��PE<���5�<<v�===#?=��6<*�A==E�<��;ϥ�;����Y;3����b�3��)��'�櫅<�+J��K�D�M�a=<Y9�<U;V�>S�<�ȭ<)��<���5����5��<��<��뼞(-=��`=�?=u�c������W<כL9��i=�t�=l�<
-y���w<�3	<�y~<��	����ЀX<��=�q�P��-���޼P"0���,��{T�s�"=���<x&U=��ޯ=1o��Џ�=�\��b<��j����*�O�<0.=��l�7a=�p=�x<p�>�ы#;'k���;����_|��x�=�-X���ün��p;�]@��f6=��k=HR<=	�I�i���4�]\_��+�<��I8-�m:���9_�q�S���l=C�<9�v�˳��y[=�k<Drr� M���Ҷ�qrʼ<��>���=��2�O��0+F������c=pG<ä}�v8W�̚��ٛ;�2���ż�e�o� �i��<�VO=�c=�Ё<	0<����㏽��=(@ļ�y=GdB� "�<�i�<�p=8�z;6R ��=3ٕ;Ԧ�<�6�=��2��.��� �d:=� �����i|���=�idJ���`<�M����<j�<RI�<�p��OI��nD<%��;��a�F�ż�F"=�p<��f�<ME<_�]��~�<�K���S��MۼӚ��(�)�v�Ί=_��;�߲<��<%b�;��
=\[߼*�7=_�><�w��=�"+��ۼ��==Ķ�:� 6=
;���|m=�8K=�m=�1z���l<5��<��Ѽl�4���=wE= O)�S�~����; �I��g��d=3�<~==z&�yJ!<�5�|Ի���B#��r���`�<̅��ŭ�<�1��q�<g�8=�1�<qܕ<+O�3�_��>b<.c�<06��m�#o����<=��<cЙ�=y��<��<Ū;Y��;���
�=���;e�B}�<i~�<� ̼�f=`�<��E��e=�-�0�]=،:��k����<=��ݻ�zڼB���GԻ���Ԋn�B�=Zn,��v�<j�Ѽ�1k:�<]���<u�< �?���Ⱥ�0�<���/�=�s�;��l����D����<�QT��2=��=�����I=z�	��z=����<
��{[=��="�$=F�[��s��1=�c=��e�g�{�4�=1�.=��K=�:��=4<��"�����+�;�5=Q$�=�=�G��ϐ��G�<I�������c[=E�<=V#)=b<(��"=="�=]n�c9=�����e��� �:��1���:���O��o{��F�=��>=�! �??�vO���;�'�=��F�tA=_JJ<|߼�ƺ<�b>��?!����<��)=IC���6�-C{��:2�E硼���<���<�G��r<��<b=��!�^2;��%��jG<��3=�����<D&�<�=��߼�q1<��;=*��<�;3:=#72<+�N�ժ�<ۖV=��6��}C=�׼��(<������k�e��~�5��e%=�ʼ)�{=�E0�L}�<���R�<=Eⱼar^=^��z�r=�Q=��$=6D��~�<C���4�,G=���<So(��f��%�<<���<4Y\=Y���U{��Rȼ��E=�����м:l�<a����e=�,<����<vxA��C��<��Ƽ)��I\=̤��@��?�3=c�=xr����=�!;�td<RL鼐J�<�8�<X�j<�Gm;D�H�#��;{�<�Z�;���<��D��k_=�0���]�}f=&<^��I��S�={:�==��<5�9=k��<=�A�>Q"�쵳�+[W=I"[<�:���O�,V$���!�o��s���!=W��OX=��=�B-=AM=��.�!=��<�m�<�a|;�wT�#�ٻ��"��⫺"�:�!_<��(=�j;���<@A��|b��C��;��d='n=*��F�7��&Y=R��<����Ӽm�<�G�<͠�猋�O�~<�^�;9�w�ğ�<��=��U=-ZO=�@�<R�������<�c���G=�Gn=��c<�f^=_g�/�u���ݼ���W)��h��������t��Ԑ<w���0��]<T<��j<�ڛ�1�o�-���{R��zSe=;6=��4=�a����<��ּA�;R�o:������?*!=�>Y��p&�R���mo=�A�C�:�]<i����5;G�=��5=Õ��kwL��e��}Q�H��@)D�
Z=�bX=(*����f�ј鼆�=$�&<!y}�,��<��y=Im��=�6=͟= ����G���a�g�H<C.)�Z�=]S�	��2��<$�G����q��<V=Ľ�<�H��7B9��<h˼��:�7�	�w���G�ּ=�o!=+:�<�芼R���I�*��0=��n�'�������]���&�v#�<�R-���ɼO稺Q��<�eU=Q<���<�iM��ټvc�<��Q=��ʧ4=�ז��	*�l�z=r���z=��+=Ǚ�Mvۻ�üjHO��A�;�@���T��S�M�l=�B���X<��=��=�r�^�2<�,O=��e��*5=�ܼ�;��U����=B=�f���������<ĥV��������S=�)����Ȼ1��U^}������P�����<逊=B�(��<Ʒ"��c<��W=�{�I�Q�[礻��)�Z�=�Y���л	�</oP�K�;`P&�8jI<}^������Ɏ�e���W�7���-=i�c��9<�p<�6a<�e�:W�5�X	�<�iw��� =���I@=ܷ��i� =9��!Qf<���(���h7�.�Z=��<
���U��gɻ9��<�Y��=���s�p=��=w:��ߑ���6��f�Jݻ�
=ť�<�08���>�9�w;�=���<�)==6��jn�<͆���j=�>�;��Q��:�콻Q���l��<�=�ػ-�<�E=�x:D񄻭��Ϩ8�a�/=S�����<b�G=�Dv�;)�j0=��<j�2��u%=����(E�={�1���=���:�Z��]M���=�v&=��=i����j<�s<~1���<�i�<#b����:�N�I��<�����o��i�<M�<�B<
���TG\=�	�%�I=�D��<��[<���ۼ���K�˼ԭ�<L����=��N螼l��<�@e����)��m��P�O=���<�	<{�;� -=��F:uᚺ��>�&��<��<'V?=�'�ȍ0=��@;,�:!!0<�29<�?�W1G=oӴ�
�����;�{�<�u���=�m!��8���i���=�<=+�'��ܷ<�q!���6==�����<|(E=�g�!�>/�<R�=}=Q=�^o9�.��a�4�]�=�n���<�m���e�]C���&=�"=#X�9_�.�)5��r�����@; ��p�I=�RI=]�O;��#���>:k�g=%ӻ;K�===�<z'=q�	����<@Ϩ;(h�����<��S=.K߼Y\\�,!�p�=m$M=�m�<f$e�W��<�����H<!�&��N�dku<��M�Ƽ~�2�����ew�n˼h��=țC��!$�����0�����<.�Ƽ����R<���<�A���m=N�=N�/�����`=>�=�L�r�}<��;�o����;({�<H�J=��S=kx/���%=_w�<}��� -�lU=��;W��;��<7�=�=M��<-�?� '�a������d=v�:<?�ۼb�\����<n�Z<�n=ޏ��x=��d=#�7=ޛȼ�Z��'DK�_��6ֻM� �q�*���ؼ���<�ɻ�1�<�uǼ�U]=*�^��=�;6+(=�u�9�<k�$�z��S��;��=rM�<��ʼ�!k���#�W=�N��U�<:h���=��<�z����8=��#<\�=�4;h�é�</g1��'y=B���k�����<��Ԭ1�;,�;�尼��=��?�$.[=�=om$<�1��[|<
�)=�7T�H�<�\p<p��=��=�LP<�v�f����2�Ki$=(#���?<k-=Ԏ�k �<��ü1���=��� �(�ȼ���u�"=u�<�lO�Կ:��"�9I��myT�f�K��Q����<Qh#=k u=��ݼ�����ƫ�Yf�<��2;Ԑ=��L����b��=�)�?�A�!�����;&�Ѻ��X=�z;=�U �C�h� =a)|<�c�'k =�������ػ�w�����n<�j$=�0;��Z=2� <  �l���x\=�H�����<�-H�g�<d��9�!<=V����k^�=2z=���<�X���=�yR<��$���><�o��Z/</�u<ͭa=,�<N�������gL=$������ʜ,=vQS��U=<�d��D�K�&+K��9c���y��=$8�<dr���h=`4Y=#=��Ӽڬ =���<8(�<+��W�<9�f=�׼*B�<Kdμ	>K;�g�<MC�<����)/M��8=ȕ���j��=�`L=�R=Ll2=U2���1� ����1<�˵<�y̺:X=/�\=		=؀<�=��<�U=���<����J�<��<=��ü�¥<礋<"S#���*<��o<�$=r2w<�ڼxV�L=�*E�NQ ��?�:��<���P�<lX��=�-��u��缿�:�0�+ӊ<������<MO��<�<�s =�&���<ݶ=�=�=x 0=�4W=��=���%���4�;���=�8@<�Y=�>��l�Z=:�ݻ\$K=��0=���<Utd�%�+�ZgC�.����V��<��A=�m�<��=|��<�r�<�#�<��!R����6�<��!=!f�=�C`=�F�<��E���6=
��=����/�<wG�<h��<������k�i*y;��b���9��,��.M�(A={����h<�X���K��E=�=�����U<	�)=(-����������<��Ƽ���6/�]T��X0==Wr�<���N�.="r�<��J��r%�wӅ<=9<x$G=��ʼ_T�[!�3Z#��v>������5=�M=+��˯E��@=@�'=j*��=�2�;^�G������I<?�� ����UV<�+p=��<G�O�T����ռ��R�m�s�*��;�\�ݼ��K���J=���<]��<�Լ��<�'�:a˪��5�܉,<M%=
�@��!e=��-�]B=O2>��鴼�C|��@M����<�Y2��B���c=D�=���<�d=�=T�
���ἁ��<wg���ټ��*�����m�S<ܰ˼�UG<�/��<G.;��G=d����=���%=)j�;���u���k<:��;o��K���TռsЄ=��;e��;�P�9�#�"L<N��=��<f��=�}��	n������;#	�smt=��j=qx;([���HH=�U;�dp=ܼ�Px��;=��-�r��<� =��v�<�q=r*��l~���Q��9K=�橼qG�<w�J��%���^]<F�= 2�<����8���B�.�����Q�仐B�:y~��l_�,�+�6�;�:a=4u��p�;�꘼�C:����<�on=�ѫ�z�}<� �;�00��3=�o=lѕ<��V�y#���E��,�<��0��+�p��8���<t�3����=�L-=ĖA=a�F=e��;�1=ǵ�<]�'���O�v�X=�����5��)���=�܈<Wp^=@�M;���~\=7-�<�a�<L��;[���8�����=�	=�,�=C�K<��<�3�<���=��/���K<5�&}=gk<��X<9�A=%E���+=伀���];^c'�7����f=FdE;�:�B���I���o=)�<-͎�Lْ�ݩ9=�E=�=ݧq=}�Y�(�^�J�ܼ�"-�g�<�]q�<_ �mD!���=����P?�<��;o���P7a�}&�{��;��t=�@��R��k�ļo�F����<�k)<�@	���k�ɼ�[�E�=Xl���)��e��S�<�꼌�N=�� =љ��۵��|�$R�<���(=-iN=Ml����<:-����X<J
��mC=ݧ(=�g���V�;8��<�yI=}�`=TO8=�|U�HH��/E��n�<J�G=��v=���H��%�Q��
�;	�w�c��cJ�<��#����<L��q<
U�������<��/�Z���P�<G��Q�<��J=x�G=� �H'=b[���-+<fx�<�aȼ�J�;�:; r=�\�oc���Z4�0<�J�<��<=��	=r��<�I]��=n�`=b?B�߳t���'=�߼�gI<�=��A=�~=��<���<�����<�(I������<[컑.=v]{�Li=4�?=y�ͼ����/��;�C"=��=]Uq���J=Z=���;�7<=3�	�̼��>=!��;C�케�G<��<�R�Os=P�<�����h<,ܣ<Z���~Q�z}������%=]�A��㻭P=i��� Ӽ,��<��9=���<!{G�m�#�n��8&<�Xa=Ӹb�&Z�<��N;�)���q=��;}?=_w�m:=�Q�X�S=
V<&ȼ�q=r�a=�����5^=����.!;�V��s�=M?�rX<h�<=�;2_ټ��=Ѫ����ym;�@&�=7�<W��s=��<M���U͇;MH����a���<0L��j�T=᪭<s��c�j���n=�`:���6�W4#���;�t^=|��<��<�7��o;cܜ<���R�<N�^��N=�g�<���<�:�8:�<V��s�!�8m�:nG�]�:��������u�'�H��;��}/n��근�V?=̍�%�^�q�<Y�>�:�X==V)=�y�<7�/�����=�J{�ޝ��-�t�8��{c��GI=�@G=��2�����:=�+/<��޼ g��\d���7��$=��}�,/=Hu=a�:�g���<Y�&�b{<�٬�Q�9=;�^��i���h=�f="3!��t<,������<� =��;����h�T�C�~R��1�s=#i	=�������<��a<��8�e�O�T�Q��==;};{� ��=''=6x�<̴���P=2,.���<�3m<�dɼBW �|�b=��)�V��;�0	�%��<��(<���<dgn<?w=G�E<X�_���/�J�<�\�p��ۥX=��=�A�
�jKD�,M=� )9�{�<�Yj����;n=7rļ���<�/&�Mٵ<աD<W�,�z�A=��=a��<���<����(E���I<O�ļ6��<nv]��2T;ba��`n=�s]����椫;g�d=\���L���=@�@=�-\���=fCݼ�A�=Xu�9�L����;@��: @�<0�¼�k���[k=A=��O=��A=U�<��;��3=��绹�<�=5���c�=H��9��,=J}s�wм��-�5��<�O�<��<D|�<jC�=��<j���;�i1�uvK��_*;�y�*L=�E����<���iB������h=}4X� ��<��W�~�_;�z= �F��Q=	�<ދ<��)=a�6�)_F=�5}��=ʔD=��ڼ�W0�U����`\<`׼�a�;C�<p8=�4D=�-=�e&�/i�<�EA����<'�
�9k1=F�Ƽ��R��%_���5=e���r=�<�<��$=���=��Z}�<�Q���q=�]Z=ݲ���������0�׷M=�0%�G�=)l�G�x�'�=�J�H�Z��W=�J˻�����O�=ž<_R#��=#�K�h�Q<d�=�=�_��&A=$^C����u�=o$W<��h=鿼�S8=)<��_ <���<�(��@��-<:����4�h��<C�.�<w8�����ei��a:���ӻ��7��@(�dB鼏�¼(�ݻA��F��<��Z��u,�X�.=OL[���s���=���S��<ZxǼ3�g�sd�<��@�U�>��xQ��E�<hFd�)t$=P �=(~�<u�=��<��c����;7==W+<��=��?=�=5=���=���T��<��_�<a�� �=;E�9)���;=��;�t�<�SN<�X�VV'=!���y��KK<�=��$=
��<�T��9Ỽ���;�����d$=	�<O���P��<bq�<��=d=Ъ�<`'g�_�K�� �<Gx��ܮ��)��<o,û{�x<R�=T�$=�%K�}�1=��=^�#�	�)=_�<)�"=��e=��<O��\�B=Ge2�*Bk��p><�����2%���w;��<�7��r�:��=E軰�\=^C�~ ���
=7L/���꼲k��f��o��<+�/=E�4=fs3=�z��U��� *�MTg�.2	�.���p<��<0��<��R�$2:�b>�˸��!*<?�/�f�|=�v<�!��< �;�d�<=b`�w^=�@w<@�<:(仨�;=s�<:c(<|2h=��m�.x=�t<��<��k�sh_=y����E�j�.=��Y=��x�\/%���
�m�=��=ҧ6��y-=�1�=�."���%�O5�<U'����Y=�~)�#-��]�<�J=��M�Y ��ԁ��%���'?=�4�<�5��s�r�\=ĕ� �6���=Y׺��=nA<8����n=��==	Z=ށ�=�R׼s�<r�b=�v'<�5T��㈼/Aj�7P���
���d��JY=�/N����E¼���}S�<W$=xr��4�S��pֻ ���S��<�<�Y�W�T'=�V=)��;�@=�%<���<O�S=��� �=�9<A��n\�;c���ʻ5-ؼ�?F=F�<	�4;��s���1�b)��Su���q=�E� r=�Fϼ�L*<�ݼK�-;�<=�Z4={���m<&�������Q<��[�JՄ�X��W��|%:=7V
=<0<�(� �Ƽ�t +=��ɓ���v[=�W�cV^����%L��<�՚;��;�Yk<<��K��(=�qy<�D��ĻT�����
~��G�'�
=�~�;�az����<�"�;ZJ���
=3�O<k`�=��F=��4=�<^d�z#/=at��X<��?=��<*�f=���<���;LO�?P��������=�.=�j7=:B<���=&ϼ�B��9Sv��!��Qa��SN�<L\%�J��<�ʃ<�3\�m\��z;�TW=�dx=�.q�{���0 =)û?���X=W�<'Z��xq
�81���=������< �<��=���<�U�;4�;��/=�k���/f=*6<j&U��^<�������Osn��ȃ=z�`���t=�-=)<�_%=k><�i=�}�<:!=�.4=��<��ټCRO=��;<�K\;���<�%�<���<扻M �����Z:Y}���Q��ʺ7s!<n(���׻,��<ZG���=G̱<UH�<��9�_�ݹ��_B������v��ԂR=�{̼�����=����ܫ��0�C9�����!�-�^��e�<���Z+��}J���� 4ɻ	)���L`���<�8<=���R�-=҈=�fm�T|�A"$=��k�]="��:7�9��<���;a�g�-=�̝;q��ld<=[Z��Z=�Q\=3w0�6���R��._=�A<7�6���=�>����<bN�h�B�݅���,��]��+=��U�y�D�`�0=A�����̻���<�Ӑ���m��C��K�� I:=���<Մ��.��;O4ü"=;+>��(<��=�|	<�0¼�%�~��tv�<�@,��f=��L����Q\=W��<(�ȼ|&=K�	�gݞ;R3�s�8=�F�<���<Ӕ���D|�Z�=)�X�B�\G�"�R����������&=�$�<K���x<��0�\��<Q�<���<��=��R��3�;�����(���;ѼS�s�=JP{<SUZ=9={�s�P)���R�������W�F��<b�<J���:w����;c�(�t= �H=�\���jz�<򅎼�ȕ;?�z=Ț <o(��I�c��=�4���~���ϻ-�<L�=O\&�QI �@�L����Oa0=R��SgG<���<���!=��)�������<��<�V�<�)'���\=.�=[n�c�����<�/.=@���=��Q=ON�u��<I���W%�Tq���E=X�e9+�G=�ۀ��-i=W��<��ż�J=[���i���<3t=�4-<	�O<fZG��BM�J�v��V�����zI������}��L��������#=̡��UUe�F6<�p�<���)���\=����!�tH�<Rۋ�T�������!%�jO	=4�=���k���=3'H<2�<V�h==+�N�����.�<]lM�q�鼕��μ׼|�{g;�kP< fp�6=�K!������3:��<�Q:�����G��oL����<1�-= DA<?.�����<���<X��������?�O��
./�:�<�I#�k��*|<�A:��N��F�{��?؝�dk
�������<˽B�Ҭ!=��K�<g,�����=jc�<kdټ��x<�j.=��<�u=���;S�<<g����<���<.4��8_<H���J0=mu�;{��;a4�t^�<�;㛼��ϖ;�mʼ���ڼ�\ =�,=��|;��v�h@ݼ�߁=��;G�=�bZ=6�M�� ��XMm�Y)J�� =�:=b��<!�ϼ�@<�}���:A<E�Q;Z��2����y���@=��h����<�l���<�Gü�*&=zl$�4;��G0/=-����;4�w�,�
=��D=�HѼ�U4=����Uh=���<�D\=�T=��I��h<�u���<������.<U<�"����t��6=�L=m< �d=��#=�x���9�ؔE�M�L=��d==�=�W
= �&<�N��μ'x='<� �<������8n�=O����$����~���> �]�����X��;���vbǹ��K��	z�\��<e9�<:�U=�഼%/=C�(�[_�����;�B+�O�;�� ��=4<���u��� $<+�V=.�Y�Myl����<��!= 6=�iG���<�� =5�=���r=4��<JR$<VtU�Dy=4�'��S��r0 �ꮳ�$��<�Q3<�-=��p<
�Ȼ"�<i�`�
�=�̼�<�^R�`�+�eFD�T�%��o�<vqX���μ�鰼cl��=�
���-<A5���=n����<����� �G��<�p� �B��:�<�65=VM:�ü;�<e٨;�����]��������J4;��%�k���H=�Z��h =�8���~�=3w=u��/!��j��$�'�Γ<�K=+�G=U�2=��G�u�{8�P�z�k�δS���'���b=X7$���o�9�=k@y=�x�W#����<�C3�ݒ<���;�M=;RӼ�0�<{F?�Z�!���<��^=n� �ƹ��4G�Trj���Y�3��<I�5�r��sU<[S���=0R��5<;�p��fS�\)_�!�<e�h;Ź �!=#��<�YK;8�;=���\Y%���V=I9�<�f�;/�1��X=�:��{��%H=Z�4�#�X���<�wG:ۨ�Ø"�	�q��dK<�%P�..P:"�;��E��5�<ٞ��	$���<AB������/�<,��<��%�l<wE���H�l��<e6I=�U=�<<96�ևn��|==+��<�*�<�; ���'��C!=��;4Ga=���r�<k�<�7j��}���������������-�==��<�]9;�t�<m+~=Ǖ��qI�Ԙ�<�A%=��j=��q�Ƽ&�R�e�R����>׼)�L=[u��YD=�i�=���<��b�[��<���`TּE[=O�|��C��AF#=�[V�u��<p����fh=�i��A�Ƽ3?=�D��X=�t`�PVӻ��<c�6�t�R=�_�9=��8��=�������fz�sA,�{?=n�E��<�@�;�{t=��!�DQH� A
=mWc<6�N#��>⼗�=b�<��=���r�+=���3>��,��b���ѼD���e�vs#���<7�`=~��<�0D=��p�[.�;wW἟(<=@yO=�R`<8���$5���]<Q��|؇<"�^�<��<ɂ�<�QR������6 �U遺
�	;q��<Z=��,=�����ezY�q��:�9�<�(���'꼡���F�(=�� �V���ğ�pB�����=�2��<�g����Z���<�g8=��:���==:�<x]��M����;=3��tȬ<,P�<���<�dD��+�X_�E_���x{�T㍼��ż���刺�*.=��" =S��<8;U<_�=c8<`k=�޾�<�=���3¼?`�<��	=�c,�W��<C=�@�<��O��c�^�ϼkE=iҷ<�j�/+U��>)=_d!<��ݼy4=(Y=��<��3=;0=w7�=c�]����7�<⬟�q��<�
�<?�i;���a6��.�t�<�������*��k�;�7<e�|<Q�=�N=��E4�9�B=�.�f$�<B
<]Z�<ғ�<�1�<U;7<��.��<�4=	̭��h�<�=�,<���޼��Q=��<z�<�K����)��<^;yJx��
d�<� ���g���Ǽ¶=�g=���<��#����H=�K�=�"=/��e�<(��9c�<�fH����;�tռQ�꼜��<��R<7f<��2=�&f��|�<��O=EYC<�º;��Q=�=�F�g=+AQ;���a����ȼ{�=����<ܘ�<g��D3�<�*�<�	:��3\�!l��۵,=�ͼsWW=��������ƺMuk����@�J<e[Ѽ�	%=$j�*��;�����s�x�I��4�<���F��3pA=����g��=���=s�>=��=�lz=��<z�⼕�I�,}<[�<��A����g=�<��<�G4=�W=��Ƽ3s;< %�0BU<S�=i}�����E�/=/cQ=��_=]߼��=���<,�;�LJ=����j�j���A���G<�SR=}���$���1=@�<8=���[c�*������<ٝ������z1���A<y�Y�>�;x�$=�<��q=;F�<�^�(ŀ;eZ �|�<�c����B�F.,���@���*;�W��7:�O=�T�<V�6=��<*�=�?~��ռZ�(��=߆�0��<>T= 
�+󻂌r��s(�^*�:�}j��'޺��ۼ�q��h;X�Q=9�$���<%�������`=@$=�z]���=D�];�����H�	�)�^�/�Z�=.��#�6=���<nS�<n���sH��j=�����]��b=� �;"���?y0�Ӈk���"<
S<ּ_Q�;5�j�Or�<q�ݼ��<��<�t=?��/�Q�`��<r3�l� ��e6�eę��୺�|������6� �=B�<�m=�j�;&X=6�HME=G�N�=	<��=3�=")=,B
���ȍ3=C��;U�2=5SA=��z<@f�<��<׶b��U=�˗<�����;�}���7���V�H�Q�����=�O;w>�<�#=Ӗy;�����迼��D:ݨs��M��<]�V2Z<�S=������=��O=,l��)�R�[����T=�a=��KZ0������:=e�Ҽ�aX�t��K� =��<M*���A�j�O�E�"=�����E�s=�@����у�<T�'�x���bD� �=O���2��u׼��D�	醽�K�`�����e�>��8A�0��<\��<��x=Z�[�B����:�1]<��<	�L=���mC=��g=FR%=��8+E��޻*r�z�c=�]<@��<�〻C#�@�@;�S��4Ƽ1'I�\N?�E�'<3U������8���<�(�u�<�Me����<����"=������x�#�!5�����T�<0GJ�Z(=�/Q�w��� ��<�z*;>/���Q=�GJ=�ߓ<5��<P�]�X�1��J��Ԧ;���<%4D��$�����a�<�==���6>6=T&���5v�n��<�Q.=Τ�<��!���=����f�W='�F�C[N��S��M=��)=_�N=)���RW�<W�<?6=�����������Sl�VP=�B�<�����躤����BA���]��0���;��n=G�o�������=ǺX�^h7��?U<9�P�&¡<��<�W�dl=����Q=� �<�*���(��re=����2��{==O�'<��	< ق����<Ӏ�<܏>�L���/��<}S���,=�Ņ��C@<�H=-�[=@��2�< =x�����{<p/"��z�<F.\=�Dm� 2���rn�����!�P:}<�`$=������ռ�j�.����a�B=V�E=���P��<l���7"�)����?<a+\=q�[< 㼏o}����$��4���=:��<��K����<��A<�-��팽��<B�H�e�M=�U=��}=�N�<��;��@��/�� )��N㋼MjZ�e�[��@=-�ϼa�<<���;�-���=�m<�`�<�B=��<���<� �;���<~�<#AR=�#
��W=�^Z�d�n=���<�G+��#=��ļ�Z=U�.����;@a����0=eg<=�^�<�,4=��;[3�<�-�=4=���<�##:油�C�@�ݝ�m4Y=�����N�V�,=k�:���;@�<�̌��P=��3<\5����=H�'�	<u�	�\���[����;H]=��U=H΃��tҼ`�g=2WV�|�K=\N�0�Ļ�KS=�+=䘨<�	���Ř<�:�Co��}�����.CB=��˼�U8=ґ�<Iq�Rڎ����;9Ǘ<io=�wZ=JX�'#<7��;=���U=�;���d��ͼDUk��9v<�T=ʰؼ�@2���<���:� r��%$��Y�<����8;=ӵ��t�;:ּ
�<AJ�y�7���8<e�.<�:�;�0?=�i9=�;�T<=� ����h=��b��4�<M���ݦ9=�=$AH����36���p���8=��9�Ձ�<iU�<MQ��hü�i��en����P
p�T�W=��/6����<o���>2��Dh��'='�=�y���1��Ѓ<fa5��~�������<=R<�:�+��
$=M6�;8)0���I��<����<���x="��k�W�&@M��l����<z*6<�C=V4`</u=<����<���;���<�&�<��<�f��Pj���<�P]=�+�;�G��"/=e���r|�<C=�f=���
6�<�bZ<t�=32���,����׍n<%�\�b�����)B.�˳�<"Cz���<%b<=]�9�T�������=b1��������]1�.��;�[X����C/#<��ĸ�9=H�8�j�=a1Y=���<�kG=}S���\=��0=��2�z�;�vA�#Ua�}l��$^<� =Y:�< �<�0=��<�i����6F=�r�R%_=����Œ=͓�<�=pڼ���}�=�P�ź)%����<��Z=+(���#.���*=)�;:RO�V������_:Q=��<\�:��T�����<�ݒ<�Y�;pAD<�U3=D�<�\.=u�;�~�Y��K��xi<��@=�ͼ�kK=���<{�G��>�<�Xs=:+=U4=+�<D��6��;ux���f���{=��3�m���b�<�I���޼l�.=}�=��{���<��
�(=��<��м�(���U����J=�7�z\:��8<�N=L=�L�<-�;�g�<0�=��l���w��#+=po?<pYӼ[6<���<P�Y�|OZ=q%��Y�Y =V���;	=-�=�nA=����Ҽ�Ǽp��;�1��0�Syf�+���=.#u����;��`<i[��Q=O�<�?W=We�;�#<�'=A'����ܼ@#;�Ӷ<�����O����=oO3;���<��M�H���}P� �<u�7��J�<. &=hy��ړ<��<k�,=-=?�<����I?=O�*=)y@==�H��	�0u#<�Y,=��[�Տ�<�RN;߸�<�/�{W��
=�r�	��:}A�<9�<���<B�`=Y>�:����=G�U=c���x� <�!<�r=T ��v�<���q��:��J��y��g�h�<w���k�S����-<S��dR�=W�<���<$�<�h/��<��/<OhG���+=J�,�P��$���I=�::����y�f�F=��0�� =BỐ�K�����G����Ƽ��=�b�<��׼#�;��_=0[���=�'s��3<��i�lX�N�<��{<�U=��Q<�޻��o��<=�o^=���N7������=a?���j��S�;F)�<�*�ڪ���T�ͼ��<�AU=���n�9��;�5@=��='1)=?˲<u����6�;?����<�2��ż̬��>�[=C��<�¼�ex;�
t�o��<�2����I=8�==�ȃ<���+�a�<��*<u���*==��D=%a��kZ=��P�:GY<B�>=$00<����+�"=��D=F���&鼆�м`���<�1���[='.W������/^=c{8=~o�<�,8=0W*<&�g=��[:R�;�0!=����8��7�<o`�<~1�<��G=l:�"��?TU�<�]=J�<�8<����#r <�F��X��v���;M�T���<��N���)=�8;�%z���<A=�*¼F���"�9�<r6��0�4=Nf�z{7�x��
�*=�B�����=��<�R��K���[L���9= oC�"�8�R	t<�G�zf ��/.��ĭ<���^(f=�2�&U��ǌ#��u��ڼ���<�Fk<	�m=,A=�E=��<>	��E�BDk;Oj<U(Ѽ)G��/�'= ��<�-��``<X���ﵼ9�<��: <=�����C�,�5=���x=JZ�<^F5��t��$f=�YF�ϥ�PǼ�' ��Ӽ��c<[6���;�d�<ɠ@=?'���&g=�q�{dG=0�=�vB�^��tD��Yd����=�f&�̒5�����E�@�<�淼Ҵ�<��*<G�(�]i<�żo�2=N�P=b������6Ǽ�<G�4=(sG�����9&=��|�e�(=�膽:;�x���c�����%��m����@�+�~<��ּ��<fC���
~<��O=A-�;Ēм#ּǒ=L�����<&*,�;>���$d�������<���J��Md�<ɱ���_ͻ�=1��<RX���:=�����H��P=�N�<���<����=Ɋ<!#P������[��t+��f�;�!A�\�'<Q\)=z�޼�DC=�]C����4=�R?=�F�m�w<rR=:rJ=�������-6=���;�=)�T�R=X���9=�댽0@C��=h�i����W�����ia�6<ͱ �5�<=e���o��;ŷr=%�~�8�:��\E���=S=ޜ~<')5=-B�����=���1�<߮�<)� �t'=y�=Sa�<�e�bb=È;�\ʻ*DU���|�6�>��Jʺ����<���<m�Z�	�<�ͷ<����S�<)��9o���#�s9���r�<*b
�$U+<1+=Y�(��7�;�.I=뒑��H��_<N@=��c:���<�G<��:<%{= 8a=
�=)2<g�0=�W=��{��q��3
�a��=�R0=̟�0��MR�Ё�����<������<?\r��鹼_�!=G���$�8��a��p��=�n��]¼�k���<����d��<T����<�x4���4�� J=
�_;P�);��$w��{��<Yz=�iM���	=Y���=��=�_�e)f<&d�x�-=P?��f�tu�����;�C���[��⎼��<d����5�=1m=��=z�<ݭ����U=ߢX��E/��"m=q���x����=�׼-:P=]��bgӼݼ#�nD�<�5��V=���:#jq<�V=�Q�S����A=��=���<@hؼ�p6=J�h<*���63+;� �;�X�:�2=�>`�h�<*0<=��<�0������= ��:�L=��ϻ�^+<Vk���Y&=!@�6���>�ċW=*F���<J\,=����=J�:=��<!��R���.�>=mw�<�VM������C=�_�F�=Lc��Q���<�=X=�� =Sz�*;U��h+=P��;�;,=�8�=By��[� ��<�yY�<�F�<�U9:�o׼a�K=C��m诼~�_<�Qs�4츻|tT;j����=�h��9e==��<��=�d��Z�]=Htּ���L�-�c0.<�eD��#L<�%��<���7�� ]=K3������?���4=]��<���T���5����� �L=~?�]@=B���mE=Rv뻲��<G��k�	=A�;����~A��f=�|���M;�dA=O��<w�#�)�F��TP=�_�� ����s�<��:i�<[�a=pF���l�!S�|�C�#{�<�J�<*=S_�<h�<�&��������<|SH=R�<�h;cꮼ���<N��<[%�<���;w��;@��j� �T��pp5�D/$<R�C<z�[;9V�<(�����<���<g�Z�~�'�g��<�r��E�j�^YQ= �d<��d�H�oq�<��&�|K=�=$���7�L�����P=ܼƂB��J
�{M�<>�G��d�<>^=�� ���A<AH<��׼�a���R�O=��1=-g<�(���]=9q:%!���g�"�;��&��<q;���;�ƪ�;�nں{�ͼ*}{<�?m�yA
�]��I�<ҧ�<f$S���<��7�b�$=��"=�(����<�����;m<(!�=kF�4��*=|Y	=�_���¼3��"{?=�ȹ��|z��KX<4*�<37<;O2[= vJ�#�*�,�-=�.��3Gc<W!(�A��;�M=�<�<�3ļ��û��6=L�l;{PL<��<-��<�+0;f6=C �<���x�|=1�I=Z�9�ןϻa�<�����=T��<Fˉ=B(�;n]8�\�<[:i��{S�gI�������d�<�>A=N:켇�; Yr=vbG�S`����h�P =b�|�,����_�(=��
����<����:;���O�0=J�p=���<�s=?AG���<g=�g�o���	�}�<ջ_��,e=��j��<�NT�D�T�DF�I/=��=�-�""��A'R��=�,�Cay�)KS=طD=�P�<��<9���/e�<����⹿<�~[�J�u<��ڼ}D�;��K���b=rd�<{=2ot�X�$;�3�<��!�wa��q�5���	=Պ$�S)9=6^<�f¼/k,=��+��)�<�n>��s#=C���0L�J���(J�x�O<R�W<��;w����,�R�;-�G�=��Y=���<p�<����n-���1�;��M��<�F<�xk�ų}<�߯�.����P=e�=��E;=Z);��i7��	=�^�<��;�J_�iG=���!�~�Yw*����<D� �$�E��EZ<-�:^p,=�	�<��E��N�
˾<�rK;~Ms<ܖ!=w�~l$����=zؼ�:<𝲼L��;ڿ���a���4�����w<q
<M}5���n=�Dx;e6���J=�W���E����*8{�Ň��R�=� `��wؼ�� �[�<��@�;�)�/<̤=�jӼڽ"=PμBp&=~�;��9=nE@<mt$<eH3<�;=���<v<q�J;�����%�<�+3�˥<N�9mÚ<��
��ڼ�<=�{�A��>.����!�B�K]�}L
=����@�O��0!�2��
-q<� =����Vo<+��<'w=q��MZ̻՞@���$=����!�	=tlB=�; =��b�i!�<*K�<�J��'E�",<C��;J!j���L=Y�<Q��<��;h�λ��<w�M;��J:z�=��W=�a=}L����<؄�<�8����~=���<HSC��^���J=��M=Xٛ<b;ӼDo�L{��vk5��B��"��Y����((=G��t=$b�;��>�K�z=����5�b=�#�AO�<��i�?�{��Њ�ư/<�۵��{I��.c=~.�<7n:���(�圷��׿��:���ݼ�k<n%���Yw;�ܻR�L=HH���c��<�<T=c៼�诺Y����˼lϘ<��S=�;��0 <`�<��񻶭(��=:�;���;��<i�K;��)�Q$���E=�Y;F)�����<|��I���*��黭,=�q��At=�o=N��=AN���/������<�3$��������2����¬�����7���6�K�O=(��<g��<�I_=�� =3:{<���<�:&=cp0�~�<&�(�:�<r_弮�g=�<S���"����>�<=���=��)b==A����U�TO=r~^��R��DL�;��=�ҡ��ۋ�T��;�>a=�Y-��w��Gl=�=���=	�<�y���O=n#Լ�����,�q�&<�`=�	Ѽ&�%=��=t�6��<��Z��n��S�<&M= ��:U����N^=֏;r|���=�H���;. <��<�lM�1<���;���<���<<�Y;X�\=ө���P�<w�=_�����h<��=se*=����#����͓�c�ּ�ð���U�q��<���4UV��Cf<8��=�Q<=P�;ř8��$��삽��o;��=?�+=�Ax�K��x�<Em=���<@���9��=�6m<~d�;�n.=z?<�F== +�;��E��V��z�m������<;»���c�D���N��<�6:�i�<�r����}<�lE=���<s*2=�l�9�R
=��D��Nd�Z���\*<�p[;y�=o��<�ZY= /�:��[��W�=�h
=䛨<L:E=z/n�oM��eH��V�*�1��������+י�4;Vj��z�z����=�m^��7�<<�ͼB�=�_J�ɭ<�^���=�r=��2��;�����^=��e�t9�w[S�:��#�9�Ҷ޼�m=�$=�L`�U�=Xڙ<ŸU�A�5��4�;6�8[c��I�^����Hl�?��%�׼��ۺJiS<�Ȗ<�Nu��ʉ��*��86�_*����/�1XE=:M�_=�lS��޼��*=��B����<%�F�0�< 1Z=�R==< �<������>���n�,���;�j�5e$�wi��m?\��[3����< ���E=-�����ն�F^��9=�eJ�m%�ڷY�W=�Uc<P�D=k7:�9ռ�.s�BY�:3��O�� q=X��<6~��on�)�~ ۼ���#�G��<����,�=��&=v|M=��)�4%�;9!�<|���l�/�5���S7P=i�<�U"�a���.>-�U����vp���ܼ�|�<ʗ�<�U�=MT=�+=���<����s���}<��Y<�j�:��G<ג=��=����q;�/��`DA=$�%=ý�<ׇ=�C˻u:�-���?=��(=��&<�����#=�<w6��G�E4�<����,�<��<��3=h(�mv���oH=�9=7�j��$����;8�D��蕼M�c��<%�8���O�(D�<@q��6y�<��伴�=�ü�. =���<��>��P=�=<��T<�U���Q=�0r�	�]=�<2�,=`LG��=�o��<Zo#��º<l_��B�	.���׼�f4=�=�;z���R�<M!n=1P��0D=����E�;==ZT=OMM��Ձ<`��J�6���b<��H�<	2ϼ �]�r�����u<,b��1�t=dF=�-=A=�I���E���3=��%�g�=�*��i��<���<�!�]=�/��'=t%����_;���e�<�a<�
8=� f������<�\�<�!=>�=xO�	���R��<�2$=�_z=�'=�
`=z�1=z;=vM.� �U��a���<���I�<	�<���.���=S�=��.��O�<a�<'�_��s`=��Y��qb<��;1sF�<�M��L:�!���ҼG=~/<#���w�;�D��\W�{�4=��Z<i�)=�1���po��F�<�܊��A<Q�)=���<V<6=�-��v<6=>=ԯ�<���<�<��*</49������L���6�%:�<b5#<Y#��VY;���Y=�Q��䁽-I���v==�t��-���[�:�	��7=��{����;OD»�5�;�%�W�(��o=p�}<
���D=$΃�s��,�0�K�=s�<}��9y�=�q�<_��<8U?��9[;�!m�Bd#��zػ�8�q�H�Dr�:�Ä��c�<]�y��=��n=�=n��#��;�<I>!<�'!=O�żv(h���L���H��揽W:-=od�<zn�<-��;q��<$t{<j�=ܵR=KWO<�UD�ޕ�:P�=ל�<k�-�g�$������=!lO=�ފ�Co�옷<P�8=�I0=%��=�Ż�C�+U'=�~v���g��ӂ�/�I������$��ST�-V(���;��J��P����5 ����go;;��+=�Ex=
�|��b+�^:I��O=�!��"�-�v��<�̙< �4=�]l<O�n��s�<�ӿ��D�<�W�<U<�n7��W��,=#=��<.�;,Z=dQ=�<���F�>4=���:�3�;"j<���Wo/<�<f��)=RqD;h����I��LT��x˼��<�u.��:l=D-�N�=S>M=��_=�Ub����<J�r���w���J�O�\=Q��;����S�;����l
�7�u;b�=�=�<��=�r6���;��=�X�<Te��"�F=�z�<v��R�L�~8$=�%�,?�bPP=�[B=Rg�<��=D�׼]l�viJ<(��=���<�:�=+3��w�H�Q{G=t��;��a���<�)p��c�<[&�<��X=�1=��<1 J=�b9<�>M=)�0����;W���� ���Y=��#����� <��=2��;!���g:�<q��S�^�-��<�h�<t�R�f΃�]���Ux�R|S��寻��'��0K���@�,AǼm����<�{<�6B���h߼`gU=86f���g���7=��*=�L׻1�]<ե�<Q�<ۮR���G=A¼	D�=��<F=u/=R�A=�(<_De=L�<(n�U���"���"<(�����]�=����c
���=��<ʽ=�s���������X����ܺ��������\S=u�'�/�*�[�-<^�������=q�d=.!p��!=I��<�U�)��;�=�	���f�L���` �6�A�֧*��>�<߱g��63<��Ǽ$�B�J��:��)=s�{�4#�;~��<�=�����	=�{7<��W��K�S7��ou<���<S�۹5��CP�.��Z-=��5�޳�3̾:*)h=P��<)
�"#���=��L���<��_=��$�+[��Oڼ �;�?��;�H_<%#='z���;��K���&=�˼"�U�
�_=Q!�<xmh<�4��Ѕ=إD��l7=0�(<��r=�=�����G=$��</�<V�N��S�a$������j�<3'<cko<Tt�<���<��#��D%=0uw=�=V��#��<<A�<m�=�M�<C� <ņ�<��<�E=�Y=8��\n/�Jw�<���<�c�/��h�:!pz=r=�P�<mUO=/>�<\lQ=E�&<��'=T)=��=tV>�('=��<$뵼�L���v�<P��EF������~;�Vܼ���:�)<=�|M=�&����j��-=��=��4=�_��L��0�"�o=���<*��Ռ��;p��2��/=�''=aD�����,`��7=Je=��A8*=J� ����<-���06=v�(���}���U\b<�����kC����Y�"�;;ɣ3��$<��ü91��us�;�*��(�<7��< g=�C=�"���~=���<��<�K4<�P-=����k��<�M�=9=��<o2^�� =�<J=��?<�����e0<��`��혻J䕽�����0�,�?�����i�<���O�:= �I=HKֺ�/��vA�Ɍ�9.c<WU@�{ӱ<�~p�o��==��<��z=w����V<�҅<S_1=�ب<����A��}w���`/���=Ӽd=�p��{����Y=ǧ<��*<3e(���2<-��<����-|�<"�7��<=/]C�3R�<��2=E�ɼ�垼a2>�Ki�<]*�峚<Z�ͺ�>���Ҙ<'5=
֩<c;;=jO�L�}����<��@�  ��:h�t�S=���Ii���A�;��V�<�n�,��<"��lm=������=��#��e�<*��=fI�<���Y��8�$=r�D�܃����\=#��_/�h��<�|<�΅=�6=�XG=���<'�g�	0b�m��Hb�<[2׻�l�;1=#��;��<�0��S==�B�<�b=��;�-^;���;�&�<QL$�k[;�'�Ǽ3U�:s�7���J��_��g;ߞ�<��,=�g&=C
����<R�`=�I=�n7��`�,���]���kG�q"=��7=����żV=A��e�ֻ�(=i���hM;��;��<NJw=:��<���cM��}���<꼋��e�
�*K|�MRT=��=�F��=�Ӹ<Q.��.i�<ؖY��.�l��%�ug�<�-�����b	=��7�S<�}=���5����<� =�%�~)�<�A�<��#��λ���"�e�<خ�<6����g���<
>�:T	�������ϡ�sa=�UE��ɼ�ӣ=@G�<��<�T��=���;JI=���v�Z�O�;Le=,>��%�<d{�� 
�̱�<e�ы��C��EƼ(�L<-�-<�U =�?�ҁ��*a=��Q=2�F��k2�{]�<����3���%=�q�_�F=φ=�6�&�5��R��H�< �x=������t��<n-�����R��<�x=���G�<��=�"W9~�.;g= �x�����n���˼/���la�<�b�d�G< �7�q�^�;=�S��ǩ�qD�=X�=}����+�<�$k=-+�a9�<L5)���<�ph=�*-�#�;cj5=I�ۼ��J�y�z�;=8m��./�9�=�М�.B��C��9&��0�<A�\��Z6�6}=r��=��d����Z3=��\�<�|���w5=k8�� ��ׁ=��6R���$Z�(\��\�<C�M=�K�<��S�>M�;����н�G���K��<9��)���[�1�.��.=b�c=h��x�κ�~��Z=k�6�P�����<��t�(�耨<z#W�WW�܂)�O뿼:�9��Z�;����Y�+�����2�s==훾�N?����H=���dA2=�K-=�%:�B���;sB�<V�<='�>=v���~D�ȶ=d��������>=h���D��:j���?�N�;�+@=��(,Z=L�<vz�hwh=�H��/=��:�災9\м�J=�,�=��<F��<I�v�l�T=��<5��hV<���K�<��P<��<J�t=��ռ=���*T=�~������V�;"��<˫���<$������<P�C=��6�8Ƿ<�	Y=ȫ
���!=.�@�+�q=��H��C@=7\��`��N���*=��9<�I=�.{��7Ⱥ��_=o��=��a%=�<S��S�xvQ=u�3���*�R�f�f����]�������^ E�d~h�|�w��FL=��;h�t������i�=�G�앀���0���o=4���N==u�<&Њ<�s,��%�у�<��J=m��<ߖ"=���<�Z�<�f��ɼ�y��x=l��F)��{ʼ�p;C��<@W<=��|�4S6=?=�j�;we.=r|޼�Y=�s�H�'=_`=�6<�⏼�v0�j$=Q�J��z��=�}T=�(�<�6���m��p���N=�F=�e�(2=�#���<��ɼL!m�Z0�<L�<��F=�35=��{�J�Y=�6�g!3����:�
=e�i=N�-���)���<w6<zٿ�T-==�dF=}�5}#����=s�y��}�n�w�Yr�V�<	O��4=�����\< f�]l5�+���%Z�����l�����м��c;(ص�R'=7k
=~��@*l=ͫ�=)2=��@=&�\=�3<��2�Н�;�����@���a=�"=�g����;"��[{�<��<|��<$��<��=��&;�����ʼ����_�|="��|��y�ռ�F�<��=��=���<<!`<�>��Z ���@����H�X=�� =8j��с=��뼎����r��3&=[*�<���us�;k!�<�c�%=�y�Ӻ�����Û�����N�;�/�[��&�<��=����B�<�T0�|��<c�_�<WV=�0��K�<��<��;C�;0�_����硼�68��b�nd�<?j=�}_�)�L��,������㼲�=��=��ҼnT=��;�V�3;�l%��FG=�"O��0���B�,�ɼyV���<,�a<c�8=��I�-���&�{�:�&伯�Z;�LP<���<��<�==oQ���=�_�<Z;�<�ޣ<.�8�'��<4k^=N� �kr�������_��܌;�yr�hn����o�qB=��+���'=m�7=��C�ȳ���s��.t_=�p�< %��\?=P!�����>���M�ز.=c��<�E=a�@���Ѽ��<����e<��,���<�3[=��,<�Eq=��!=��<��=q��<E��I�O=��mi2=�1�<kʐ�P@[����25�q6v<�0���g���l^<���<	��%�!=C'���cK<���<bV�<��Z�b`�O�	�y��=x�:#�W�F�ط�<k��;~os<�Ǽ��c=ʣ�;bT�<:Z�u�q=��}<����S=�h= 0=[L��ƭ:V�V=��<�Y=ь(=-Ӏ<�OL�
"ʼH�p=�Q��dO�j/p<-p�Z�Q�;[��y%�1-=�<f4M����L3V=��'D���N�S��>�<�K=7�;(�7=�`8�I�1��<+=�5K=P���duR��Q$D='����|=O�<@0B<Ya;;��<k7��\����L�"���;n@��S�<�|F���2��~��e�<���GA�<��F<��[�w']=f�=�E>p=���!ng=Z�<��<�[;�%=�*�<c�M=�=��Y�	<S����#�=���B�ѼƗ���;P�<�?=��P=����Ƽ��,=��==�o<�m�$�<g/���<��J�0�<�ϝ<�U=��;M�%�q�C��/=�h����$M=$�7=+�-<i?�<Oh�<�	)�D6@�"�=���<x�=o�<&�s�94=f��1�R�}�K=c2�<?3��%�;�簼[[��ۜo<�y =��S<��=))��=���<4o���ꦻ}\�<Jgz�K-�<<�)=�	�8n�=h�<�^|;��@;� B��q.=_�_��W�O�=�Iռ+Jb=8�%����<�G1=����V����<�=�:8=+�$=l1=�|t�h�5=��C=������1^-=d��;�I����)��ꙫ�_=�<��J=���<^��;��<pPԼ��<����=y޼��=�+�������>#=מ��Ô;��x�����0@�i���Y<�A(9_�<��=�ƴ<����G�=^WZ�<!=��=s �<x?��8�_�0���� ���<��2����<=�[<`~�<a|J���=a`��Ɛm='��0����<'�u=�Q=�'9���<��\�*�<B�S�Dо�h���&�<: �<�>�<��<qԄ�>~<�٨��Ȅ�۔+=��<=v�D=�{-�T��<xa&�Z*E<�l�<��K�i�<0��<��6=I-"<�����Ժ�7�?=�&l�]��<M�a<$�V<=��R�7'c���<�tQ���<D�r=T�ļ�-�K���===c�1�����<p H�N�i��'�� E�;�\+�u��E㼮�G�nW!=A��<L��<1�<�2;:M���f=oA=��n:=��1���;<<�.�kޟ��Lͼֻ	��ف�6��O[4<����`��@=�� ��I�����eR��{U��):�l8��Z��O3B�-�I����a_�<�F%<����UJ`���<M8���;?��<�u.�Đ�;��-&���ͼ��	��$=�n=���g��<k	'��U�<yc:ωn���<%�%=T��`bA=WCr�ֻM=(�#<9�b<c��<��A�<����Y =~�5=�X �(E=GnO=/IX�X�p��]�<��e:�_q<RYG����<�ڮ<}:�<�D7�_�=��J��S �L�k<�	�;�=��[<`�K��)��^�<;�<Á���a
��,w�� /���<0��4Z<�(=���E�E�-�4��I�<}�<[�m��m#=���<�n=�����P��l�<ځ&����<9�����%<T�'= =5��<۔�<�;�[�"I�<����~��٪=�ҍ<n���R��~�<�\޼�t�;�#�>�J�q�<6ވ:ɧ	=J|:���<�Q����"�G��<��;��E=mx�< ��<�\�8 m=^D�<����<�N;��	�)>&=�X��=h��0�-���<Q�1=t�<��<�/=��,�~,=�<�=�}: �Y=V=�������b��	�<G���ZѺ�JH��閻��<9e�yo�:���<�tW���<���K)�;[hw��c��O�!�:�����X%=,!����<�i,��Mļs*���P=H�;ˈۼaM ��gS���<�N&=�s=�n=ȧ	<�%��<��S<��W=�0%� at<u�JUZ�4Y=F�/<��%=l�;�-)��H���P==�x���Ѥ��<�2�<�˂=����Hɼ�Qf=86��x�0<:s�<�c��[���7�n�0�A�y=�3�<�]Q=�Nu=Z%���?���������ѻ�S̼H�=��"=�)=��_�	�1=t�+��1�<$S�;�ͼ�O�h:�:�5���R=��P=��_<�.4�.39=���;��;��!�  =��:�Cк31=i�Ud5<
h=5��:��<3�m:

`=[��<�%=���BV=�A��Fa�����~��*������o<`��ɹ7�A�=��=v��;�;����ʞ���I�ȘR��盼[gH�aH�<�żi<u��^/Q=z���啼��7��)�=�=�M<*@8=U�g=�X1���;O���J�<+��V��f�<�Dq;���!�����=��ù&f��B��<�K\<@�9�Xc=+�߻���΄=i�=���;�)�=�>���;����*��wJ����<��d��G=�.5=���<٣��I�|-<�7i���<m=�Z�<^�?�] ��	�4�1���Ѽ�u�=�~�
cR�����}�?� Dy=&�X�E����b�Y�Ҽ�=д=`i`�(d���)A<'���z�ݼ��]= $�<��^<���'��$s�:�}�V�I=Y-�Q���t�>�u�<g�,�v���@=<�"=�rU=뛓��^c=,�,��7��>xؼn�=�:%=��û ����}��W�<�<+�@��bD�V�<Xq =Od���m=N��<���<(D�kY&�p��4=�8�g�b=EY���Y�?'�|���$���U�H=��c��� ����:��$��q�<�$Y=)	=	Y<=b.<={]]=�Q\��
���xӼ��=��9��z6=;3��>�^;��4;�h���'=��"�n���q^�ΐ	�e�T����<�DP=N��ڟ<@z����\�9،��L=�����H�M+2=�Ҋ<7�`�kݡ<!��<�ŀ=z�.�I��<�_�<��1=m���&�<�)�<�=(m=����=g��1z�<�j"=�(�;��A=T��<_7=No�;tF�E۴<��лfCW=�V-�η"=#).=]�ܼ�?���k���߻<!5��B���O;��%�t��<cCG=ߠ<����H��E֎<�T��� = �u=�E<�����==Q������Z;_"���+� 8=T�+;� ��7���0G<��<�^C=�����
�<�-=���<��s��s�<+��<���/�-; ��<�5�;�H��5yO=%¼"����ӖW�y=��\���,�弫��;�� �v���� �Z�&<ͧ��2>A��(=�>c=m~��SN��{�;�'���?�Wi�<�椼�EP=B<=a=��%=*�V�8)�p-=z�^�D�<�'�;�;��B=.���%-=6�����@�=�Լ�@"��);<� =�=D�;'-Q�tk]<��/=�O�<s���G�<�ԅ<�=�A(=��;_��<��<�+#	<�PM;�_G�3�6<֠%=a�D<���q�%=��)=������8�6�.=���
u�I�0<#uY<�ã<}�I=/}��RR��C��V=���<H�c�2�<�B�:P[�H>:�=�jH=
�<�J���T=����������$��:V�]=��R<(����j=r��<�Q���SQ=U?�<6Q(������2=ՈB=��S=�� �n{��\:w<�S�7=j*=�A�<�"!�n=��<?��<�~?�h�{�����=XO4:�<G;�Q� ���^9�#�6;���怼H�<��"= S�'��<3�
�wGp=�P�9��E$�t�T�e�9�=y�0]8=�">��!�<�<r�,=�w"=b"�Gz<�S�<��+<�$>=�]T�Ć+��^7�ћ�<$7O� w=��G��M�y�>��E��[�<Bt~<��܏��Ώ�����`�:��]����=���<}F=�P��OK=�7<45#�.BS=��=��@���=
˾�q��$�;�D�<��~��� <�b�����3=8�.<�G+=�W1=-M��6=�$�1��r�O#=R��.�f<�b� �O<"|=�#�<�2i�ٷ�<���;�9p��']=	`�Bi�=�<�h�<�Ǽ�FF�=���F��<��˼���� �	<B���U��,=���;+AA=��<Y�Z=Z���D3�~��<�S�<v컼�
ݼ(�D���m:0��E���P��v�{\���{���ݔ�KVV=�&��D�H���<)�{=�+V;�tS�4���=��/< �=�)�<7:P=��$=4�7���<!=��4��@W=�w'�4��q��<����� ~=ke;=�s:���%<���<O�<�߳;Q ��)���������4"=��9��,=�{a���D=Q�=�M��X=���,A<��<����{z�<��üy�E=��`<b��3S����6<$�o�[3�:7�E�Xx�=��<I�J=7%�q���?t�xe�d�<�b��Z#�<�(:B��<~���b"=8T ��/�=�V����%=�	����=��-=i8���ʣ<vpb�X�n;��'�SB�<�E��G�;`=���<�ɼ�<7�%�<W����寮�������kX�s��\�;=�r��<R%(���ü)%���_=�t=
�R0�qŉ� �=�"w��9;��[��{'=k�G=�`�.�;{�<�Ly<?��J�<$+= s!� �T=��G=�`�?�=��=���98�;T[=�V=z+��Cr^=k�\���<r_H=vEI=�9���/<�K`���;1�=P��@ )�_�G�g'�<\�R:r����F�8ѼW&,=��%�j|$��<�;���;s�<��0<I7[�^)��D�<��:L�X��<�?/�g�=uN���[M=�\�<p'ɼ�ꝼ>z���0=�?)�
���LJ�9�"�=E�ڵ=�b�š����E����4UG�Nr,�����	����F�;���< �<s?��g��J=ŜӼ��<��弻<���S=k
����z�4�i<�O�:,��ʙ@���h���=�|���S=�W*=`uļ�������1��<W]=�03���K<�|=�!d=Z��<n�5�&�u<,�\�3Q=Sġ�H���c�=AU<�b<�x�����;����2;?��<PI�0@v����<��������;t��b<��,��E��=ӒU�`3����=�-�<]�T=���<Z�� �;�����'��lq�<�$�������*z����<��<��Q<�`�,!���<;
=�:���;�o�<�P�<3ʰ<�%���M�<ΟM�fZ�<E���B*���f����Q�I�A�<�;�:?je;��%=������-�쁛���l=�U%=`�=nUI�����d�E��g7=��;A=8�m<�4w<�kC�J��:�'i�<���;A/=��<=��:��==κ��Y<�#3=�3�<H��<�zx�"�=���N=o�3<{[=�M�:W͡:I��<tkȹ�́<��P���<�����<�#�<W�V<�����y7=z�:`��<�����=�7t8�`S�[9U=��2�[4=����07<��;X�k=���<�b<�{ؼ���=����,����}3��4=�]�RM�<��=d��^�$<-��C�<�)j<!�m�����!���<�������!�����<������������\='=��U�<"IX<[1���h<�Z��e��?��;8���+;IW<�p;=#A���T��O-;�=H_G�
.�ĭR<��<=�=�y=!T�H�=���cX�<�z�RK7�'���B=c��;�s�<����U�����<�W��>=ڇ �_.U=�K7Pm�<v�=�&8�  =_K?=٥�x����ڼJ))=W!��|	�z�P��F.�䯞;00W= 4��ˌ=�=��ռW*�=Q[C=4=V��0%����=�;����GeZ��1�<�F=������a=]���6�9����g�5� �|R�<:�� ���d����<e��:�iA<�pݼR�'���	��m#����<w(0=�T9��]�A}��=1t=^�*=����鶣��H�<���Y~�%.X=q���<�G�[�5��g �~:=2�I��B�=�.��c���g=�-�bf�<[=+=�����Q<n3=��N<��'����#:,���<��=�g��Tܼ�$�;���}��<ӛ�62�\W�<�uh<�*�;k�q<��D���A�l�h�Kx=��<��ݻ�w�r*�@��<@TP�k�@=Z������Z�μwe�<��3�ټ�"�:	˜<��s�G�<�A�<Z4B<H9��J(*���L��7�N<T~,���4�rY��=��<���<���;EN9�lU(=���<�<'O��d)����J];=��	=�Z7�~�X=j���<�z�����<=]��;�Lѻ\̤<W�8=��̼l�0��̃���R�I���b#�:�*k=}?=o���c<^�=�b�I=�ļG
3�3�c��v��s�<U�@=%��8Vl�퍖<|�<�R[���N�x,>=��E=����Qe�r��B�Y�iZ=B�\�D7=�W�w���tL��B�<�q��m�	��4+�������=�=рQ���<Wڼv�J��c3��jܻc�/��P��w=�뵼��<9�O9=V�o*���.��.;��=�b�<��
�t���	V���;P���Y�=.!�:�|<ܾI��ٴ��� ��x��<e���<�/��N�Ǽ�l={Ӽ��ϼw�9=A��͋�lZ��f��9���<}�J�	�;Z��cZ=�fV=rXB=�#�<�jd=�@�<�Y�;��μ+_={퓼�׻�E����]�����ܑ8=�e=p���m�9=�%=d����=Ԗ�=٤N�s?���5�؆d���;|E�����ﻀ�{���</�l=�8�<x�v�E�����h9=4��ã�o-t=9�<YtK��},��Վ;�Q���;�z4��,�;��;�����<���t|�<��H<)/'��?<L�ʻ=��^W�}f輒=�0=+(���c�<��=�������1�)=���,��B��*���Nռ��Ҽ�6R<��<ѣ=8#=��7�k�B�1�</��<֋�<4�<�Q;�2t=e�=��+=��Q��3=ԛI�4�l��(��������`�l]���'�v� �C�S<��A�
���y|=��E=x���Y��P���B=�}*;�{>�+� ^!=8��<��Z�ޢ~�!�}���-�#y�;�N&��n
=��������<����6}�<1�<]�R=%�'�叶�R��݅�<R�-=��C��I=�J=�N�<��)�����:?,=A���c!=06��J:�#�a��ƭI�u\l=��6���*=�5��O�7���i�q� �&A�:w4=F=��$��nݼ$HK���9��$~=*�3=��W<@4�<���<Hj�<Γ�=��3=��!==�P=�H=KW_<"����Ȇ�۷g=��Q�׸=Kh8=k�	<�]=['p�����xU=np.=j�?��:G�7i�<�<`8�8_�y/�?���q=�i=��G�����<��V<�6���0=҇
�JO<E�	=oM��*��\ju=`��Q�;�#���2<}�j=��¼������.���=���<�õ�ݐ2�ş���7�<��5="8==e��᥼c2+�&�1��$ȼ�3Z=][��R��<�x=��a�bٌ<k�g�����=�F;R��:"�=�<�*��<�Б�OZ�B�J�Ӧ#<1� =�ǐ<���<����.����μ��<�мk(��]���$=�S~�i�<=��=SlZ<y�v<��=E{���Ѽ���, ����˼w)�<�Qa��F���=����
=7s�&�\;s���KH=�=�]�<�Y����<�<[�-=,�=<��=m���H�=�=z?#=����{��<k�U�ʇP�?}<��=K2< �K<��=,��;��<�l���ǻP=���H�k�:..��O�^#����<�ˀ<�1��x�<ޢ�<gF�<�-6�p]�<."��E[�<�`.�fT(=s�<3}���uS;�X<v�l<ܭ<�$=��H<��"<Ϸ=�iX:ߙ3;������<Aμ蹳<�2�<ϼ0�J=�N�<���M��ٻeX=p��<�=�69k����)<y�h�1=/��<V�A��<[f��!Ǽ��5�r=��=q�?��/�ܯ�<ҩ�<�[=��W�t�=hV�bc=M7=��=-<T=�\�<�W���O��>��~/<g�6=�1b=֊�p�;��]<Ԟ���y<E����4�D!<��=^����d=�K��}�&�<ɽ
=����Ŏ�F=Ļ��=7V��`ډ;)2+�f5���8=��)�<�ܼ���<��q<I�<����TLӼU=o?���=��H�N��Y��o�K=��~<Z38��6�s%=��=cY|=:�#<�0���>��
�<�Q�פ{<��<y(0=M���D�<��^=fP�<"�<_��=ք_=��>���ʻ��I�v/x<�=<'n��j<�����ϻ�W�����ֈJ=�dS<�ػ�$���V�<;�0�q�<���-dd��=�=x��<��f�A0=�Q=�m{=�lм�<�xw<����=K� ��C<������@=X{��Ά�u�t;���Gev=K�ＨZ�<��0<=@^=`=���4�"M�/���(=�ii�H����;�ﻼZ�@�#	�С<��J�+��<���;��_�����١U����;M�=��
H��"�r�c�B�=xڰ<���<����vpz;-��c�S�vA�rx���/���мb��;�d.;0��<}�(�d��UJ��;H=�P�;n\����&=�[�ሼ:�����:��q/=� 0�Dk <�ԯ��]=O�ͻp
�<���T*=T�2=�TD�+�H��:�<�
�;YKK���d=�]5=��k;�ǂ��y�<YWD�f={au���?;4��MyT���'=�3<db
=��B���h��{b�<�%W�j�~��܇;���<�lҺ�X��=��3F�-� =P&=�=�	N<S�s�k��<G�><d� s�	����Fe;~�<��;�4a=B�����Q���8����<�>,��&�;��<B�4=��e��e<��&<zki<ڊb���ڼ�6��Pλ�Fм*RG<A���m>=;�U=���B�<��<��$=���~P��Ps��=훼P1��"=��"� ���f=0�n=s�K���=<:��LH�f'�<��	�_{��)<*��<��<F�Y���c��YE�	�!�f� ��<=�Ma���R;��E=��@<�_�<t�=@�#��kü�s�~��<�b�����=Ru9��O�?
�|�D�(2D�f��<�
�<�����`��:p�<��<�5�j2z���#�$䆼�G=�4�<3��<��<}iڼ`�~<)g$=����=i���
�𽙼4�p���G�=Q��5�<n�=�"Լ�����u=���<��1=7�μ���;��@�$H���;&�p��k<����#i[="xm�*+=���U_)=���[p�5���W�08#�sY&=�YҼ,��<g:�<�=Y�G�<��;�� ��=~"=��9:a�Ѽ���=	"=��ü��{�,��e�=8ɘ��I<��Z=�4μM|Q=�z弬�;®�;[�<� 2��Q�<쥍��ຼ�V�< 7���=�iV<Cw�<�㞼�؎<�ͻa~�;��3=�s<��H<��8��4v=y�`hm;O���;�n����o��Z�=Wr=,(=��<h)=���P5�+��<��<�-�;E©��H=z�8�����u��^!ɼ��
�6ի�pI�<��s=�	��ૻ��J=��c�o�=�X&=^S=ĺ^="BP=��K99Iݼ'����;�		�0RD;�{%<E�׻��C=�T�<PeP=]�׻T�/=�����d-=I�;0������a�;�}���g�<�G��;�Jy<%��ǀD�������!=���<oE3=49f�~'��Ȼ<H^�;{��<�ˁ=�Ζ<Y�<�8E!<�lQ=k�@�6����==�rF���<�Te=�4={`�<5�'���I=�Ё<\yd���ؠ��:�Hh��[�7e=C#=Pl�O���i��=�-V�v�(=e9���9=k����l�:�2;�_�oUu�
��v�@=&�J<��Y���?�.�<�">=����-�?=���=�ؕ�r��<���g@=% <�o"��~�<E�	���=�9���;�	���6���*=��D<�
.��#-=^�`=b'H=>��<�(�;�ͤ<%;R�߀�ư�<vN�8����7���a4=|�%�i���}	�[��<:�A�kd�4��<8�G����t�u��a�<#ݚ;+.�]��<�`p<��>=	�Ż�*�<].�h�Ѕ�JU=b���Q�=�~m=�ٔ��
=/�>=��j=K5�:�2<M�Ӽ>��kI�<��<.9e=�4R=ҽ=���?<��E<��;��u<���;�I�ݞ���d�Zt�<)ޜ���ļ|%���u=�&@�ʧ<#Vp;7`<���;C�(��W�;�M���;��a1�7�ݼ̅�<;�-�C�=;$�]�g:�#�<
���n}�<���&��<��T�����<���T�R��p�;�)<=%i!='D	�az:�[=j���2<zE�͜M�ec�<
#��������A�A��<���<˾��d@��N��X@=!�=H��< �2��~=D�������m�s�\׼a�@�}L8��=-��<n���\�B�=�<�%<��Z��*���=G�qڼ�2�;�hJ<����S=���;��*�5z��f=��;�ʼ���H�6=a]�������U�=�]=������U�<�48=D"���==
?�<�?=��;��<f^@�Z|=�Z��e�ܹ���;p�N�#�==?�;=�TZ=�c=0:�(��H˼�8=������<�<�4Y<��=I4C=&`��丼'��<^��#��
��C��:�TE���<��"=K)=�,%��_=��p���=�Zo=�]L<���d��<����:�:��%L�=��`���:=���<PӞ<��<�;X=��<�Ҝ����qO��S:=�=���E=��]�8�<V  �O�<P�<��<q?��_�0=~d����=��J=��D���[��Yd:@gݼ��\I;=&�<2>ܺd떼^uJ�x5p�tR=j�<iHJ={��;�L�����(<A�����=0�C���E<�F�E|p�����I=�s#�S�ϼ{*���<2�{=mx�<���̫<�0=����<����U�:� �B-N��N�<���:z�0���<����*��~H�"q<=��m�,=��:=��2=�N<~!�<���f��_E��gC1�	�<	 L<{�ü"��<4� =
_�<�X=ص2=8�<ԥ�`[s��]B=%5<�)~�q�<��=�{�;��+���.<�vY�Z�=�K\=�1l�i*�5�5=�=ͼ)w�<�1�L��<��F��01;⪑=6az���弡V�J�K��'t�F?�Mqo�� ��w"=�|��~�����J=���;���;�p=T�(�=����Z-�<�'�<Ѹ�����<��i���F<\3N=�"������Լ��^=���K:
=@0�<�?0�������-=cA�ڮs<<���]�<��������a�a����ꩼ�����<�k\=�N[�k���0�V�u��;��=�&w=&�=�J���є�<��#=��=>�㼤6K;}U=�z��lW=H=;=$�X��"H=�\=����F�<P�:	;=������E���A=�+�;����TJ&=�W�<%:=��	��j=�q<Vt�<��5,=����ynt�Շȼp硻-I=�i=�}P;��B�T�=/
h<pt�<j�b<�n���r�<$��8��� U�<�H�I����f_�.$v=�q�����<$��<�^g������V=4|=�Y��1�kk�;��@��h=�2����U��N�"���s��pӼ&�z�@T.��o�<�9��X������G	B<�2_�xC�-�f�h�N���j�Tn8;ε
=)�
��.7=R=�ϊ�v�_<pN��� �����8�=��	=���;�Ȃ;�!�#�=m��:���X�<�ȼ͸ۼ���<7O�=>�2�N=�#=��4=cՄ=�#&����<�"���y��f������N�=�DüQ�{�d P<)Љ�Z�m=�L�<��p=*�;����3��"<�8G=��1<1c�[4<�R=4~�<��x�*�;�a����1�=$�W=-UL��y�� �<�	=��T��њ=�y�<�?=��7���[5<�f�P�����1o1�B^N��^1�!i��:���<<4<�D=�Ŏ��[�ܓ�0��<�X�<�=�]��ȳ�<�~��^z׼�=:��p��<;��=��1��J�H�;�4:4��<�!8<gς���"���a�xg�����<�<C輔k]=X�s<��������j��Tm=Ia*=�lt=?�U=�|=�H�<��f��7�0�$<���n��9�--��j0��ݼ�'s�iq�E���/�%��dbg���A��%�=ǰ<�~=����=;�h�v���&�<��f9+�]����=�0=8�ú��#=B��<�Y�-�<<'5�o !=1��(<�ދ=��y<��=%/ǼC[^�F�9=�B�c(Q=�㠼���<? �p��8�{�`;k�&�#�����<�m�6��<V=7���<�ɼ|_=�{r<���;c2���e���"=�x�ܕ�ϣ�q!<���=r��;�(��P!=B�B�>�c:ea��������K<�#ܼ$�㼈�=_r=I���n�<��2=Zh<<	�q��$�E �<j<K��<�D<�[R=����;�9�ǌK�����T=3�7�~w@�L��O������V�$=p�5�c=^?���=doU��}=�X��q���Y�k=ఆ�F�=gV�;D@.=c<��<F�<���<���cE�<l&z�<��<��<R�[=��<=8O��S��;H�E��6�NO�<�w�k .���4��b	����;������ٻA1��2�I��<=(	!������L�ւa=��<��X=��<=�c�-=��7��ǫ<'`��@=���{D��4=.'d<C׮<��@=�.�<�K==B� =��~=�<����邙<M�;��_=bR�<=�#h=E"�<Ź;oH�<+:�	�>�Й�~�F;q�[��s��ރ�F�<�@=:Ә��ވ;���<\��<T�'��֧<�F< �G��H���D�<�"�<��;�<Q=0S�<�OL<�Rm��D���$=���t.= &(=E���F�8����ņ<�q����;#==���<j�F���`=K ;Oc0=K�g=��!�Hva=�e_��쌼�R0����<_��<��$<���
�\=��6=2��;a��<�0����=D�F��68<�y8���=�5��ǻ�9n�g=�AQ=B�C=�\�~�"<N�/=�'|=�O=䗍<W=��^<e�M:oR2�mH�ce�<���<�Ѽ��g<��=Jy^=��޼��=)/I=������e◼B�iM�=�;/=���:=JG�����<r,]=���<�k�O���h<
$I;��G=z~�OL?�^!�{���f%\=��i�(&l��(d=���9+�y�/=�#=����=����J�<�s<�%e<�ɥ��gݼja�>�4=��<|&=_�R=�cO����;��Z������R�p߼jt���t�;�2H=�ד;M�Y�h,	����{}��?V�������tF^��o�4#<FV�;�1=�S-=�'�<>Q�;�,7�5��;9ڼs9�R��8�="���l��>���2= Y<�j_�>(7���6�RQ7�!�z=���<x�3<��Z�{:T=�4�I�6=>�Q=�Ĵ��<;�r7<�?�A��ו=/��OBQ���P�hhy<k�X=g�;7��&=<��eA=P�ܼ�%���}<�=��	=���H�����|=v��<E��=dST�N`/=��c�l�J=7qü���: �C�?��<]�<��h=*#��ߛ�m%N= e��+=��h�ʹź�wY=�>=�����j�żN�=19��{9�˾3��ޢ<L�޻��A=�x7���E=s=�D%�L��<�"�N���M�;$��<����<=�\<��;��u_��<T��]�<mr;�໷�9=�J}�}�;�;t1��P��� ����P=�&׼-=R�����e'Z���$=��=FFb��h�<6���d�<�Rp�=c�<Ttv�|!�7h��}R=�N�<m^�;����J?�< k�N�F<EC=�����Q<r�_��6t����<PW2�`�Y=���<G��<-�&�N=��"=��̼�m��V���u�<ߥü�l.=��%�y���r�=/r�<��R�L�;��L=�kh�\�b�B�<�����c=ũ,��:�<��<-��<0�<�Aw�=d	O��*;��<� J�_=H=1�㼵(�J�h���<��<�f��m{�+�D�[�@�/= \�����<�ǩ;"=a��=�G4�q��ę���z:���<�m=���՞<�<���#=�d�ޥ�')D=�..=h*<~J̻���<���<�^�<)Jj8�6=ya�<n�k�?�=�Z��Wl��S=cp�<?��+����V#:��:=��&=��ټ�V�;�]��J���4��#�O���EZ��N7뻁�J=�=��=������g;�ck�!�<�,c=�;{;'�+��s�n9���;a�"��j�<gP��$M����<`�6� ��<1�޼Ъм�	�����~�;��N�f\=:��.8���tC�WԲ�,~�<�#^��L�<��Y�ĝ�<CZ=%DY�m��<P8^��<(�8<�����;y�=�G��J�O=]m_9E�8;n�7=��1=����2X�A�"<!���I8����<k�T�"�O=Fu}��rk=��G�/ټ���ͼ	A9�Ų<Z!���T���L<�<_C�9g<�:P=L����<�)�<ҷG=ea�; �u�������e��<B;�<�*�Z���e@��J_=YJ�<b��u��;P��^�S=~�=-���D�r�Z;�e%=}=V����<����c�O=��;�-�<���\�_je��(�=��ӳ�;Y�:�-\��Z�<��s��}�<y�x=<�f;�vY�d���mp=:�1=��O�P������R��<�9Y�ݴ�+��Z��<M#���{	���<���f=j�]�-)L=w���i<�n=�==-<=���%I;�o=JË��R���<�se��X0=_n=���켼��B��<6����5���b<\xK��ȇ<��&=�	��<���u�������<��!���d�(=��<�6�;�.���wY<e=�-�׼�I<�|q:.�k����+��������Et���:�o�<v�� ���Z\=_����t���-�;K]K��9Z<���ˍ+��gn�������<�3<��s��g��Pq,�$�(=��6=�*i<x�"=�j�<���(�������w{=�c=6��=
�U���9=G�w�{�ʼM���ۉ\=%�=�6k�|=隿<MҼM�;/\<�"�B��� &=]Ey<a���<4盼�����D��X��֍<�ba�r���+9=����ktl�zl���t��#P=�U{��B��<Mk�<� J�����JY\=_��<1p$��|�K�UȤ<�y_=��<=�q�������O<҉-�K�m��ϧ��뇽0�<J��<;J�@�+��C6<�$4=2�&�+Oؼp?=�F��͇;�A1��v=p�<��H=B�=T����C�^�=���;���<��߼��ݼ�x�<��<�6,���=c=����<h=��z�<Z`G=�j��=
}0��&���+=��<�dk�ݪ<q�$�h$4=�˾�(��<��w;Ћ6=pT=CL���ԼL�y=Rhn�T�=��J==��ڼT�t�#�e=�q�<$=*l=��\=���<MwƼ�"=��=s�b=D����e�Y+�%u:<�����:�S@=󂛼\d� `K=�N�E��"�<k� ��Յ��>�7�-��� =�)�XJ��!��{�<܇���L;}/d�$�Z=ŵP����<��c�r��<q÷�+%��y:"<W2��G,�7��� ����<�;=n�9=2���P=Q>߼�HR��iF=O=�G񼔜����3=�>n=���;�`�<��<9]g<��<�qm�v�g<�=��T=M�	��+A=� <*�$����;-��d�?C<(D9=«=�d=�~�<O�S=�MV<�ɠ�a	V<�˻�D�<��̼�s��׭<���nB��A�`��<��Q=o<���8켡t��T�e�}#�<T����<�<j@��l[W�F&8��z=��r��~�<&�L�1=wP8=h�<E�@<�\����<vG~<�F�<�E}�5���{�[�7�<�==l���-0\<S=�:4=�?}<B࿼��&<k��u�5���S=�-��D���1=@f=>���~�<40�<�/��������96=��g=ܮ&==(A��R�<�?;�Q�<Gc�<�=<V!=5=+�&=2Q6=���<�㘼�ш<��8<5�� �,=�#ټԃP�����"�;��Y����=.������;�q�,�6=e�W=������)�ټ8M���9��|�<�(�sT�&�=�t=.�z�^��:�G=&�<�;�s��2C=%�<���,5�b.���<�Gc=�dH<.���~�L�h�����9��=LM"=!=�<Gj=�Wo�B(�<R9@�#;u�A<���v�,=��a������<&��<SFE= ��<l�<�ۼ����=�Y<ŕмGh=��_����pR��W��C�����[�<�p=�a =M��(�<�w�u=�J<���x���D=��;��5=_҈��<�<-�!=/3B<�O�+Yf�A�<6���,��<�����=��i;��V���n�TB(=K���!�N=(�o<� �B�}<���<��=���10=��a<���aO��LN��֡�#��;�%�<K����������W)�9��q=}$��a��� �c!=�x<m��Y�=u�ۼT�m<VI�;��>=t�p~<HK=U3=����8&�W>�;L��tt=����?~��=;J�<�]�<ԁ���K=��<T�=r>=ϱ<=�溼L���sN�4b���x��[��UE=mX�=������E�y����:eO<4[�<A�e\R<��;�Z���gػ�/k=�ƌ�k����p<3<�����j��`&<�5U=��*��	;�&�F<N�=9� �U�?=�ۑ���b��.�"#��5=<a�,��d�".S��^��pP4<�4=�������<�r����K��=~�/<	�:=m=�wN��km;	U5��
��f�b�T=�)=S���GH=�=�Ʉ��_�<~�r;[��;R#�.+=�P:���C=��4=��I��5��N�س���,��K��n�:߈0�ɑ����<�����:�*�;����0\���|�*	%=h��<@���t�ݼI�������	��@��Ή��h=�,޼J�p=��R���;E�<[l=�
^���
�75�;,.C���9��[�,)ż�W���ּx8�������<H�<��o�哼H�f���i�����(3[��D=Vǻ���_�����<�?b�KvJ��[�%��<HG��}2=�M�J=�n�<<�\���F���z�r���y��������� P�X�s��պ�e7<N��G��q�^<3�]=N0,��y=x)��߷���ļm.=�=���I�I&= Fs=*2�:�r��4=p�l;��Y=�4��<psJ�	�� ���<d�9 �q8�]��c�<�C�<w,I�#B=�F�<�AѼh����W�<s�=��<�R�<w�;垼N�b=s{f=��K��Y����<\�=d�� 7=c������<S׼>�k��M=k��<�#=�Dr<�\ż9�<� S;�<F#Z�P���j�1�z8��.��Ͱ�=�y���ʼQ�<�f?� �2=�`�<���"6k�{�ڼ}� <��:�hL<i]�]�< =��3;��=S�j<�zI=w]}=֕��䇼Z�i=Z
0�cؼl�`=Ҍ�+@c��TX=ZJl���<��ּ�=�@�=��-��e<���;��<Y?B����9=� $�e��<ף�<�\T� `==*��"��A�=��<G��<�	#=�E<c�d<�'����M�3�/'Q=�ϼ�'z=�<��S������C�<g��l��8;p��<��W��� �=��v�"� ����<��=nk��06=�z�St=OI$=[�N�=�<�m=�0<��˼�0=��9<��=[����_�m��xJX��bv��L=��7=�]V=S�<ܱG=JOػ׼�=�r�Q	�xm=ͨ�;q����;� ��[^�<6+��A�;(t�M@꼰�3��2<��D<�м�Y=�<W|��Z�˼]Ş<$�ƼU�=ctͺd��<�;�����:��<H��<C��<�u�F��F�j;,�;?�n<��;,�P�U0�;�La��0�I���Zb�E��$�&�T?ؼ��8=�S<L�H=�:�iQc��G�����u
�\�:��<�>�;�o�:�+U=�>�=t����k\�%��i���*=$j=���a����C�{�5=�a;��ܻ�v[�P��<���<{�H�3��1�5�i$E=�-� H=ӕ�<����C<&�X=R�;�8��N=�؂=��=^�=��N�(�^=D��<��%���e��*�=8��y�=͎<�մ�z��;�pz<�KK=ꇈ�ay�;�=�$<U4��L"N=��"<u�]���.�� ��#��;�����/<H=$�N;�"��H��<�*=����4��.�<�芽t8k=�R;��̼����,�� �I��<��0������e�����g�<�t�%6=���00=s�a����A�Ѽ�9���<.�=1�4��;���A�ٔ=s�c=;)����B=�0�����NT�<�Pr<+��+h�.=�μ�y�<4�@=4�v=�)�� %X�-s>� >D��o1��]ռk�л��<�����i=�Cx=� �<s��<���<�C=��`=���I���8<�M�{:��3�
�e<	p(���;��g�y�`�U��<�h����~��`���"�=4!�8|3<��b=�N�<y�<bI˻�HY=����av=�,���X=@� ���~=�ʣ<���c�-=<�
���/=N���+k�=��V=�2��-N�}9�L���7`<�oS=�N]��O�%g =�ƥ<�V6�T�=Y?d=�������<�ܼA	<^ �1�< H-���������4&�I[ =�ç;��^�D�U��=,��9)S�=ކa���l</�����\��3=\M5�NN=�H=�@�<�<}#���!=��<t �<�&b=Yﵼ�O	�����VQ<������5g�<*��;���^_:���<��T��
���O��$�:��<�1-���o�9�D<g�<��<��#=�~�<>֯����g����=�P����^=DP�L/<}�缝����(;�W<o�=3�<7�<l �L�|�K�=��`X���C��l:��P�!�H�F���[�;t�ӎu;��u=��R="��?������<V �8P2=������|�d��.�;9G��ռ���.}���6=�5>�(xV�`Br��u\=TI��^=+ZG��QV=�$�<{��6��<)��;����k<}�(��J?=ݴD=��>��mQ=aɲ<-�J�s�:�19=�X�~��H����<dP=	��<~�r�y=g����=BV=�@=w:���c�<�,�H�$=��<��<�(0�T	t�XR��VB=�Mż%���q ,=�G�<�6	=�<U˿;������˛�a.Һ�y&=�F�y��<���<l�8=�!=\Q��χ¼�뚼�޼ԑ<�<�;��R=z�<Y�q�h
�k$=����-�q��#���&�;Bͼ�O���A?=��<z�=�?��F'<��'�~Ƽ�d<��=����c<gK=���<ƛ�<@~Ҽ���<,<�C���#<wǉ�/�:�.��ǆ<~˼&:�6�<���<Ն= L.����<zF�8q�<����	�˼'���D
ɼEa��<�\L%��P�<o�����<�����`��F=+I��Hˣ<y]=u�G��<M`��<�� =�u�em;��x�8��9��<H燼N�
=�] =��?=Z��;�����<�D���=c�?=��=2t�<+$8�)_�=+=UH��~=?�~h��{��K�<�:M�n<�H{�s��<W�={ּ;:��X����'����<��a��К���=	�<5��6,�;�	X=�6=Bv><-3|��͚�WF���j��b+)�L����8�����{�����<'^0=�
=�`E;���R�=�㭼��<%z�
fP�m�<.�e�Ń=.2�<�OG<�v0<7E=�|�<�C�<H�<b�м!5A=}��<���<��1=�(P=$��<)��<�{<��b��=�h<�r�;a�λ�=��J�Q�=>Vi;T�{4�<[O=��U��$;=���� &=F��4(��,O3=�[=��L����'�A�6�\��{��C�����J��7v<���<��}�93b<~�5=��r=W==�0 =6�^�l����<弦3�=FL����<g����J���9���I=�Cb�S�r<��;��\=GD�<I#�]~�=���<R<��_�<�\=�ݷ��������H�=�k�<'M =�����¼m��A��=�U"�x���|J��t=�2�<�H���b�"�%�G�V��R����<��Ҽ���:G���	y�=~�����6�n,����=�k�;l��<%G)����B<)��;'y�OA=_b$�X�5�s6k=�2=��ݼ��a�-�h=�As��R+=s纻)�<}&
�Ɍ/���4<�X0�VD9��7A;{4%�q�<�����^�	���BN<~?���=0=�ea�g�/="Uϼ��A���<E+:<��M=��[=�:P�.=��������p�=�1=��_�ꑼ��=��<��F� �
=��<���{�����YK!�r <=W:�I5�*{� 4h=�@�;>,���'=���2���q�
�7;��q��<)�z��I�a�ü.�<u�T�N�8���=�3���Q=��=�'�<:C;�������ͼ�c������=�M���,����;�ӂ����L��ة&����m��;�&F=���:��n<��#��#!�e��`��:T<���qK=]��<��d<��	;�T���=U<);�9���v+=��T=�v<=�ٝ��t�<uIM�*c7<܏<Ӱ���|���a����s=ۛ�;+NA����<C����hk������<<�[=��Ӽ���i�K��*=AE)=:�A�--c�n�=�!=�v�z��E�d�4�ˉ=}��<�I��<�1=D�V=m���D=Pj�;s��;�u��T=]ED�n�z=��X=F�Լ�����׺<�wh=���<L᛻Z����:=�\>9x\9�4=��3="�-=�
Ż�B=���<���;#�; �f�aL-=80˼*�w<i�<*�q�e���d�C=�q<�=]���:I�y�<ai;�s�<���`�<s���-9��&<U���ڻt�=�2=�%-�)9�<�	t�N�s�f<�ό��o,����<�Bּ���<�憼�$����<A�G=�~v=�����s=l��;��%=Q-|=R�K<���<�<6fͻ�q7=>~���3�}Q��������_�� �i]�+ļ�����G�<� l����;R��:��<���<'T���D���7<QkZ<�} �p6=���d2<� =��<�$�]��:�=q�>\;v�Q=��fi������Ы�z��<�����l��D=��Ƽ�꫼�w�(m�`�<M�I���j���%<$%�C�J=`�����<K�z���<-�}��������t,�K�<�{�}
�<�?<Y�<bO�<]�!=�/B���ʼ�B5=5,�*�l�QU=2R�f�w�܉�<
B,�lv���8=dF��m��<"�������\8={���e#�<`�L=P��<�X�<��c���S����N`M<A�O��;z<�&)=��X=��=�RK�6h�Du���j=����|��:���D1<�E<hK��-D=�=�j=Ep=`�<��P���P�x�E�oп<��J�����s�����AB�?�=�+�:��������v=������.=���<�7���ee��]2�)1O����M��$��M=ם���X=�%��C��2�;�5 1��MM��:�mZ=
�<B�b�e�R���Y=��Ro=�6=^�P=��5=�4=�4*;�;=�(�e�<�f=S&`<Ԏ�<L�U��Om=��<
�=�־���O���<+�=0n:�9,�B�<XX�s���1*���5��A=�AԻr#=#���%���o:?Pl<O�;���l=����F=+sS�#>?�*�o�@�h=u���-C���E=d��<C�=ž��Mq�<��==��<�E�ntP�~���A����<������꼟�кv�\����r<ÿ���GP=ݯ���Ai�x4!=��=>�<L���p�<�$*=FP�<rj���k}<c�����T~1�r�n�}�׼9S6<�%̼u��<��<�<|
d�0G<�ym6���=�R!��\�y�a4m:b`�;�|��S�\=�1�s�<��1��9r�]��\�}Y��2�^=_� <���;fQ=C�ʼ�Ǽj_Ǽ�r�<�� =H�j<cu�:115�g9���J�]-�<�~=Q^��<U{�<��d=�e���t� �[��<�����BC�7X@=n��[�<�����<�Y��N�<��U=&Rټ�-;U�ɻ,$����_�N�G=�U�<t�����h=��<� <DB
<�>��k=��<�Y��W��>t<>�>���Լ��;"���{�4`Z=[��E)=�f�vT��Ql<�C�<���3}��)�D�p����J<���iH�`O�<	T_=&:��=��=��P<e-�<��*��0���'���<���:�����:=�d���6�ԧӼ�J(���c=X�N;��#2�<;�V���:�f���u5��b��y\=݋���ʼy
-=��<g����<g*��Y�v�7���O�+��:r��~�==r��<�H�;sY�@�>�+=0��<.	L��7=������a=�y�<��uB~<Kd.�9©<�m���=�6>�
=j�:�!��ⱼ�ۆ<���)��\ݚ����'q*�8U=]Y<�:ݼgW�<�@�<&;���1=�GZ<���'9�q�!=��ʼ]r-=�7�N=�-<<�h;������ͼ>���ܼ�<���<t�;Y1<ؑѼ	cz=��y��6�TK�e���H��?y���}�;F"l�����5�;��
0X=��ûY8M=~';,	鹕OQ=[�ؼbNo<�,�xW =$�b;r=u�M�Gڿ;�,=�%<�~��K�q�o��b=�E&<�cϼ|1���%=�� �"b2=B^P=�:�;��=�XE��$�;���[S�` <��Z�+f(=S���O�`���/yb=HRѼ�d/=��⼲Y��g��S&�aF�<��q��Ա�G��;��<���<f����j�<�V
��<=a]�<�����0�<2߄<��V��u���<؂�=�d�MW��he �$׼Դ=�U�=�M���V��a�)9^�����<�=��	^�^0�<��w}�<� �.�ʼ��m�3���]�a�;��?<�_<<3K_:�cK=����9=Q =�L(:%��_Z8��5�<Vs˼A\F���%=���<��
=��+�U�����<�]���M���;<��<}N��{�<�4.��V= ܔ=,5=2�<4=�vq<6��< �� �G<A�7=� =N�<��;Cu�<Ҁ���$ؼ|��;����IP5<��lz�:V<|c4��x���9�<Vy7���:օ�@R�<���<���qE=��=S��F�d=�� �(�^��D�󲍼�!=������w=���<l�ƻ�&�:c~�~�L=���� ֋=�v�;K���_�мQ<;��N9=3��C&λ�ѣ�H1D����m�:�>����<��<Az���~=�N���{�<zn-=��=�N=Fl=݋W<�8"��J:�玽
Қ�������f���%=%SU;�<䖿<C-��n��<�@H=/9��'<��^��}�K�k;Wv�:��?�U���؟⼘
^�zd4<Y�N<�$���<��<����V�5��<D�<�@_=��<~W��I���tB<>��D	=|�ƻO�P�xn#=�ɭ���=,p]��@N���,�-�'{J�Z�̼�Q@=��@��)0����+�<
�;�!�<ř$=��	�)ė�GbZ�Rk;�qI=f=̃�S^&=�q1=����b�=ߺ!���컉�	=W1�kׯ<n
�<�ێ=ӑ�LCY=�E,��������RGD��O=� =�i �J����	����r-0=�N<"|�ʪ<S�Y<3Js=HvG��V@=Z�<�+<�֌�]<Q��t�i������"=J��<��=�t��4ļN=��<����/׺�;�WH��H:�e�4�]�1=�~�H/<|���¼��+�kn��n`�<op=OO�<B����1s�<��@�/\�<��=�|��/4;ȟ[�k�.��T=|�1=�<�g�>'=����뼼[8��6�<�}�<�f<�����2=a(r=�K=���]�#�qf޼TW=��=c�/����ϣ]��{�<_�<��<#,=���e,��w�'�;V�;K���;.�;F.���%�L��<A�p<e��z��<�l=*���5�=��/=T9f�G1�}<]���<�[7;Ft+�o�<b�7=5�<n��9�����< 
<4g7�Y�<��T��=�J���f;�za�#h�<� �R ����<��n��H�<��\=��<�3=Ǐi=d�z��T�W\�<~X=@;Ѽ�H="gA=�>==t6���<����X���<e��<C!���M<O�!;q#F=��<SN3�5����т;�V��KCn<.aK��"h=��<}�"�I=�v���^$=��l�� {=o1ڼ;�'�z��<��e�d]�<w%̼��%���=);.���=Jd�ڤ�<eI<�=�D���鍺|Џ<Ո��L�=�U=F���#<���<M���+�<�c%=0F�<�T���,=|�¼�k��Z��K1�P�O<E�ݻ��<@�����=�G���i?�z �<�dM<k=��<)<8���<�U����ʼ~����u��i<�\��������;p�`;^�#��A�ʀ�<��&=Y��<�C��==�D�!�A=�?������2H<����8���0�'��<	�E�G��<��=�rf=*�~=3=�]�[eP<XZ�;�`¼0��x\9���_�����֭{���w<}W���x+�M&�����'F;?=�^&;�v	�S����=^���7<l#2���6=Vv|����<���<7/�<\_<���VG
:A;��~;9�I=���<�y4��]`<�8ݼuɆ�o.ܼ�cO=�[&��w=:B�='� =
=��<B?!=o!�<�1G<
=��O=�<k��I<{T�<c�弣�Z�lX�<8(O�hUo�n���P�=�-���q�zj.������#=󠃽�q�Kc	=�l;�&�
ԍ�[��;#��:u�Y:`�v<�+B�o�Z��T=e���b�<��ۻ�v����\�,�)�2�c<�o�VE=��Q=9ἒ�1��}�;޻:;�ټ5<��g�n1G<é�<��?=r:=�h}�����x#=�4��7;wڼ<l�=<װ�m1ۼ�0'<ŵ��0Ǳ<k]�T��<I츼p�X=�ݼ|�<�;.��'��kV="�{��ry��:=�x;��=��p=�G�<9J;�# =$�y<G�&���=~`=G�=|�T=Y��m$�<�)�8[l�W.�=Jx����=Z��y8=	G=\o�<��=��\<!I��v�߼g�:����gp���o<�<=��<魞� �Y=hƑ;T#d��ic�O��<�?�<�f<�&����<>A=u�=���Aq9��<��oQ�o�N=��,��+5�ܼ��K=��#=�XD<��,���;K����-�KO���Mm����M�	�KdƼPHV=�MA�G�g<0߯;K<��[���`�[<x4*��B ;�(�\��<��9�; y���-�		O��(=��2<`+��`=�A��5[��bb<�f\�un�����.}=�|�'�'��W��Z(�Kx=��;�+�C=*�=�[{��N�����ջ~Ƚ�h�5���<U�;=�"N��"�; [D����6|Q���j=��(�+=�� ^=}e&=�QL�]*��������V霼�J3�N3�<6=2C��4��<�5��N'<�^E=��;=V�!=�6�S*���;�ǃ���8�( <��:�ȼk|<J��w?��|�<�<&��qH=n=��<n�=��=5>=�wA���$<�oR<��ۼR{D�d�;4�<A7= 2o=��<�D�<=3��*;�^�<��ʼ�I=�G=)�ɼ�$=VT���,���i��i�u�L=���<�X�<71�tx�<��)=�.��l<r-=k�(��Y���==�A�)$=�	I�(K=���9��s���0�m��;>�<�~�<��*<I=7�\�"]W�#CQ=�^Z��Vj<|g�<1 =`�< �<-��d==R*<��Ǽ29<ĩ{=�.=�	`t<�Oj:>�<=raͼ�gP�-}?�M�_���<�H��=���(����%=�n�HX�*B�<��$=��~�*���gN=7�<L +< �{��
=��#������ؼ�q�~��<�J=�fO= ��<�!=��ټ�R�:����a�H)=<$V��{=٘��O���3=�i=?~~�]�=e%=_J_��̼�g��"�<�E#�8b	�Lּ�m����M=�[f�
�M=D"�l�/:V35<��*=�HN<���<���<B�c�]�;Xi�<�N=�Jü��̀.�Q|Q��'���>9f2=���)ؔ�-�E�ŋ7��a�<�ީ<��~<��:=m囼�I1�Ә�<�Q-:���<NK����<�S��HԻ_֋���X<���~p��v�	=��2;�=�p�k�U���3;鎼X�!=��μ�e����t�U�0<XP�<�E=Ϭ�<����W`=�1�ʎ��TT�<[�O���n�&O�<k���)�켢�+��[b����p��;6L��l8�ƃ���j�<�	K=��Ƽ�O<��=S,S�	�<R ���F7�=�<$Ow= �H<�J`�7�=��dz7=K=1��<e��п�Q��<�3<��,�P���>̼U�=���٦�<�x�<�v���v���8/=)H#��t��Д2;�s>���<�5h�#�h<d2���W1� ���Z�z<��_��o�O�`��`x:�f�<v4��Զ:m�<���<��]��������<���~Ӻ����}y�떶:��+�.L=��E=>D=����#&=�<���*=f�'=�(��ǬB;������6�](�<l�h���<��d�ϘI=�Lo=�3�<U2D��N5��O�<k�h���'��;
=m�=h��∢<�<��p�X�K=g�%���B<�|��&;y��hl=@���+k"=~I2<U�_�L
�<�=1=3�ǻ��:=�=8CQ�%��<,���n��	<�w=q85=��<��=s6X<&eм�==|C=��a��=pi����c*=-�»��Y�PWQ��1;�h��
O=�J= ���>=�*�<z�=��<!۔<F��<�-,�BZ�<|㫼�#�9�=|ݰ;�<�<�B"=f����E;-h���;�X��/=<z/$��6� !缺3���fJ=M�����<�v�Q�&=��S�pi=�<�:#<�]�r�@=˸�<�o�>��<A^޼1�� 8%=�ڛ<�g4<�P�<��^=��f���=7T��@�<��!�؋q=]��<��M�(�3=.�8=P��<7}T<S�P��IJ=��:@�
<d)j�.�_<��Ơ�;�;����_�:�8��L�ّH=K�<���<��=����/y<`c6<��;�홼e$�<�=�m=�j��=�/*�k���9����<���ߝ��+�&��]�@��10��: ������=�mK�˼;�G����<���
1�ץQ���/�o<�6r=�D
=��;h�1�02��@"=Nr��tU��bO�<�m
������Rт���;'-�;���<�/=j9==���+n�<8�<�3p=�;Y��M黉Hk=�$<U=�Z��Y����<���&�qg=�o�<g<*h�<z�=ѷ0=�(W��CT<e�f�	r;L�j<N��;����Xڼ�-1�~���he��gS=I�\�X�<սʼ�a�v�S����<;f�=&~c=!����=��F��+�<jv�<�"ͺ��)�dG=�h�u�<tJ?=6zZ�(T�;�~<�y<�"Z=<w5�<�`-=��?���[�=�I<\y����7!U��i��	=VY=�"⼋�I�d��<��A�Z�0�R,����P=ns�<b�z�d/��a�<�[&�dP׼�]�/��<�R��w�<��Q=lp�<��;� =9=��<.�k=�MG=aIz���*��g"��$P��I?=UKH=)��;�χ���d��t<���A="nټ͈)�`J
�d�6<aD�;��<M+�<ZĜ�ż0�9*������4����<��)}=z�
=��h=	��<�Z��򙼓3�<�I0�>?v=F0~�NM8�)B�v�4=ϡ=�������=�T2�ކ�<K��<ZŢ<�M�e�&�:���1^?�cb+=L��<l��� h=����������໧9^�D����X=� <�{Ἣt���=���I=��2=��;<T��;Fa��Ƭ�X�:찹<��漺��<``�<<�<�fE=#H��ȱ<6�<9,�;�B=�C=�a�<���<��G=��3���H<?~��n+�� �^C�<��#�� ��� �7R=����v.�Ҽ�6��>;�c��Zy=�LM<��Q�(���gu<��< ;�<"�𼦬 ��:����1=��;�,U<�+��=�=.=�����B���b�8缾щ=�/&=��N=�n��_���=�T�*J=ˁ��H��;��<g,!=Vg�O�3=�g=<�%=��Q�J9;b��<`Fl���,�="�<[M<=�Y�;h��.�=):�<ր�<��9=|������q�&=�ñ�Ce:p&���q���̼F�n��:��[�:(+ּ����<�O�;�Ӽ����_*=���'��p0<�"6��'��ͮ<Uf�;=��<��P;ҠQ<���<�|\=�>j��,ۼ��O��;��uL���m��d=�̨<P'�Z�k��5��@P=cx�%�=-΍<�@=_�:�c ��y�<4�;��zm<�m/���d�Q����@<�R=Y�'�/���ѡN=�d=���;A�Ǽ�	�<��.�7���F�W=4U<��=/%�;L[=�by�.a<�9=�OC��ǋ;ç<v b����]��<;�G=�e��6�:=kÅ:О=OQ<4�J=����ħ;k}8=�<Q-��eW�<��Y<��^�]. ��B<����e9=��;%��<H��)[�R��;���<,e���P�/�ɼ�'��*����C�#DżF�vl��鼿�<�ђ?<����A�~'��J
=k3�<+�q=��[�c�<��
Ç<Y4���n=��n<�=T��ZN��,yQ=��Y�)�<N��|YF=ב�<`Ź��j��ʗ�3�»X�2��vh=i���=O�C�+j�Wx`�*�"��&�<��j=���<���A�]�T�tн<D]����N=,�<=bI��m='�˙f=�m�<1�L=�=�L�@=��;C�=��?&��~�5�<� D��-A=�-J�������]��5�;��H���2¼�^<�A?<v<���<
"=S�%��8��=� =�:��S�b��Wi���<��<
����=7=fW<��\<ʵ�;��:=$q�d�<4S��r=�� =إ�<�/3=�=�E=�X���}6;L^'==�R��T6T=�u,�|,��[��<ol�,���-����)��<�/��%.�U�T;�8j<��<^��ㅽ��F��,=y�2�Qnܺ�˻��<�\��C=�b4<���;"%p=$�$���e=�!I<��S=�<1=��x�k� �H�[��)�9�==��Z<nwG��Y�K4<]�=K�:A8���A<��w<ڑJ=\G�8X��<�|j�[m�<8|żҟ_=Y���A=��-��=���f E��q�{-;
k��cŮ<o+��ɝ;��M�X��<mE=�T�:�6=��:"۸<�)��O��(,��Gc3<c~�Ĳ�n@]��x8<ӻ�	T��\Z<�>��kL��j`=�%p�؊=�e"�B�	��Լ�=�W���%ü�^=J<��߼Z|�'�-=��=	=�<ҡ<��[B+�aA ����iL�*�p=��O;b�h<�1=�)�<�%�;�3?��#<�ݺ\�`��s=��f<ݟ��e�R�%:Ϻ�ϼ`�H=�q�:^Z�<k���_���l�; �.=��{=��/=�"����m��D�F�S�;��=F=�'O�ɵ�!�<��'�ްh�G#���<��4k���#=9v��U�<
�=h�2=q�s��=�s�<�(����<z��ˆ;�	�<�+%=�
�_���<���<�������# �\7=5}=������R��9�y�;=V<�7�`�)�""=�p������)2<��I�V��l=���<U��<|_�<8u#�8�r��=���;�?��~!=��{�9��<�>�<CVj������'���<(�j=I�;�@.=h�����p���<��Y=3�]=�<��3=ꢷ��,��%��9�/�٫c=6e�<<�<�Ë<��1=Eո�&P�:����wO��{T<P�.�%�j=�f=N��9-(P��$�-HR=M⋺ȼ/�`#�;�W=��� ݳ<}��<``̼K�;{o�<����,Z=��<M�=�i�<Lc=u��<Gc�I�`��Ȝ<9�&=�$���!��)�ya;�~�<�d�^�2�ޚ5�#G����t<NT�<F<�ŀ=��+<�꘻�@����N=�[����<j~5��:�<�>��Lr*�ib�����ݒc=1ZW=�H@<3K(��qH=8��<EE=O�'�9��<|/c�9g�(��<�<'��z���6��w�Q���	o�0B�� ==�����H��`%�<7�X=��=�I�{6`���.=Wz�<W�h<x�3�O�R=u�<��l���0=��׺��=�4R���/��/O=622<���<R=o�-=�ɔ<�p�j�=vB�<R4_<}�9�*��<�ő<~�;ppT<d�K=�5<5ԕ��)N�a�]��G!�ހ(=�?=�s�=�0�<h�m�=�<d�9�v����Ȼ�����2=�4���U=Sa[�Lq=�o��(Ѽ��-9�F<���=��[��G=b:�<<N<������V�%=�K��'��Q-<��`<L�+=dR9�$��<A�;$K��蚼�#=��@=�F��#h=)��<Fż�ޒ��ú�$�<q�';>󟼨��<�h�p!��|�����\�*⠽K�:��D=+nS��f��#�����<*��q�N��u��a���sی<��C���˼�P��D=�};=�X)���$="Y��x=<��;����ͼ�s���B��i]=���Ls���>=RR�<��<�<�u!�e>=��l;�r����5*t��>=�μ)�<X�;Y=�=k�1=rF��vI����#��T6=|��Aj<Wb0���<&�J;���<_f=k�׼e�U�w�ۼ��O��	b=� <�,���-�[
s���=$�<��X=�-=#�w=��p=L/%���<Lޭ<<_=Z�2����(�?�-���0=�0��:�;��FP�tE=��0=a6<�
h�г8��V�՝���7=�eb=i�9=�CQ�O_��[`S=~$�����<�g>=�=��׼��.<	���?{k����<�]Ƽ{j��S��Sy;�'=Fg����D=uS<���;�_e=hR�9���<!6=�$=��2��=I`���Z���R���<h�)=Z��<|N=2lU<}o��Jh�<M�N�5P=Q1:̩�<@G=��=s!���B=�y���S{�<�u<�P�Kz��:�;�a&�ZRL�u���L��;��B���8����<C�;+�=@�fS�< ��k=�T`;�!<��ܼ�%@=���	%��;�L��l�<)m<o�M= �|��3¼b�^�:j4�ƚ3�J):;I=�%(��=�y���ʼ�z��m	�;��0<_��;*={��/�x<��(���{=W�!;&�(��j=r=R=�e�Ę�y���'�=�y���;��8<)������I�<������T�pƮ;G��;����D¨<���;/��<l�	=$��n�&���:M�<s� ��q���O,=�c���<�zg<����̷=�t�W=@"�0�<ȿ�] @�M�X�+<=��%�ۏ���E�E��=I<S<f1Ƽn��<?�5;�L�~F�:՝)�0�b=�O�);�T���j?=�R+=������< N��3����^=>��6:��=]��;l*=f^$=gqd<B������;0l���6�);� =}ZD=�c=�~޼�� �5���HG�B��v�2=#�*=�&I�6��;K��Eρ�O�i=9=���<�W��=���B�L��k�i���ݼ��B�48 =��;��[�ѥ�vz=_( ��f4�)e/=*=�z=���V��zgx�f@9=P�;9&&�RR����?=kx~���»-�;�����"ȼ6��&=ݶV=�,���/=p�e��GX=����fv�H�<��v=�(=sEH�K�=&���Z{��� :��<Y%{<�劽-�=� ?$��fY=��T=�U#�O�żq;=�Y�ׇ����ԼhQ[��40=O�.�N-�Y�&=�Wi�- =1:;�C���+�,����]������{<��S��C{��<�"xt��D���\��=���x|���J={H�ٜ�<�wQ=�?O���=�ǻ?�+=y�Ҽ�z�<��k;��<�A�<7�#=��=��S�TB<?᧼�T$=i�;?6E�R(<�݀�*���<ޛ���x�<�_<�k)�#V�L�A=p�2�},L<&�;���<�-=�;��2���Z��?���Y�#�Qv����Ƽ�=��;v��<�Zt<Wq��L~=�^N=�<�<=��#����<�� ��1����<�)=���<�;��*�l�E�,͹�Q|<�+��'c<��<je��=�<+��_zo���<�%�<��h=����s<#Mp���U=Ң��ݻ<�X���[����<E�w:�=k�K=I=�R�<��m<��/��g�Gb�<���񝪼GG9��Q=�eܼ�����2=j�
<Mg=�2W���Q=htK��nD��g��І]�T�]�8OE��D�������)<(�X<���G=R�<�S�cQ=��'� )c�|���I9<q�@��L=BM἗=O�]���<e,C=_~����!�6�;��%=̱,=PD�<��J��*����<@b�#ʢ<�Ŷ��c=�,\���=�X=�1���,�ϋ:9o^w<�I=����xa�b�<�Y�%R�ƣ�<8 �<�q����7�7
e�ڼ��mB�<|�o<�.c�� R<��<t�{�Z/=���>P��D��IN�����ͼ׮�3�Ҽw"u='�V=V�+�ʯL="Ģ<��:-;O���%�3<�DV=Ų�;
O��������<�
5���<�% = �
�~D����G�QJ�<�!=�=Ȥ��X�	������ǆ;���:�/��O�8�g�n|�<�J$�c�2=��+��9ݺߋ>=�ȇ������,��w�<�#�T!E=�<q<a�<�+u=}o���ꃽO��<l�<�Y��_3�);�Ϛ;=�	E=xD��Zh=:��H�;=|'������8=�#�P�=�_<���<j��<R@=��=�S=Y�\�x�ټ �r<6���=E=7�V9T�o���g�Qq.=X����\5=2$N=ߓN=��2;�ţK�+��j�ͼ`7=�s<�AP<QIp=@hC��Xa���<QF=�1?�lqK�쟨�����,f�`�c<�!=�><� =>HO�����XH�=طȺ��:=����s�AR���k�<�ټh4&<R?ʻ�w�JrM��.�9�ü�*Z="y<���<vX��<'l��y��!¼<�;m<�/<��&=2dO=j:�h�=�m�<�/�#H��H�9<>.=��9{�m���j�蜭���<|C׼�yY��kQ�:��<�Q<��G<�P�;�\=6g=��J=4&�:���<`"[�uUX<%� �o��<��ݼ�$�{����=�H�<M۲<an��X �p�{�ؓ��!h�<X�d=�bo�k�^�J<َ�<=�[����|�<��<ډL�·W<Q$Ѽ���wc�9Y���]��������㈼ ��u.b�a�6��Q���QK=��O�4�S=�,<1j�<�F��`=�q����}<f����<���<��,=�Vx<�6������<r6�=r����T��A�<b"=�P�vH�;7#;��k��z�=2I���2=�H=��<w��<e�j=�{���7�h,��;1<�j'���<�[�ݷ�;��ؼ�Et<�[�;��=,�/��NZ����<�R�<�:t�<�r���;��'!�2�{<��x=�O[���5=���<����K=Q}<b]�;�}U=�fo=Y�.=@o>�36=n��<4�3<�)���ܻ�^0=�a���<-�c�}9�<D:�%Kq=D�'=�V�lQ<��\#=�b���rL��K=���j��<��&;0]3�*LB�K��o7��#�<V�:�[=zU=�sh�,z�<��<F�#=��1�N��<v�&<k�<{�C���5=�B"�y@�<������>=�95=� ߺ,�?=;�.<`Sk�^�N=�(�ü�2�����f�P�~<��p�$=���<N�O�8�B=�{ڼ����R��I;�y-�У;d��<U�W���׼[HK=���p��X�~��<rM;��G=���<�b�Ť�<d=�.�<�@�|녻��ּ�<��<�Q�V���4=�(��=5�C<`r���"=[��=5�$<��3<dj*=:@�R�=��	=�+=��b��{ =���R'��A=,=�U=�焻�
�<ue=�_=M�Lro��ב;58��(ټmJ=��� <dwH�m=�F���:��P�:/[�=���A	7����<ݳֻ��Y�	�]�����?=�-@=��>=�ӂ=���<K�X=ʙK���ټӼy�����K��:�<�ϼ
��=Z�U��#=�f=HB=��H=uyl����<׊=��ּ�l�<�^=c^@�7�;Q����,K<C���;4<`wB��:<�cG�joȼ�r2=�=H�5=�=�f�<;`�<�����g��o���b=�S=׆���j=�U?�nȚ��W=�\�q=��w��"O���b��#���=�R<� [�ׁ�<��'��M.���=�=�3n=ۄ�;�t(=1�h<W%b��M���f9���m��>'=s̼u�8�95��;��=��O=�S=؉���n�PpD�Y�� O��<�a=��?�?!�<h��<S�;m_�O����s�<�p�<ɰr���ڼ��);�4��a]=ޙ�~z�=Q����N��]<N%h��5=�'K=��ټ�~c<K=d1=ğ6�]\�<�'�H�y��<���;��<�߀��	}�y@&�˿=)#=��T=�7=j� <��j���D=�S=�Y�<�==(���5��6g%� �0����<o9O=��<�����굼��<�S�O6�+��<�		<`�N=�A&��{?��q�<C*��,=��	=���9Z��;��<x��@2={���a�I�;���Q��;���7F��ּ�Sg=��1=7�#���<yV�<}n^�
�A=�{㼜�'���=�^=�=��`;�'\<!M��`�<ٗ�<�E=y^�/@o=5�D=�D<�:G=�F�<�$��׋8=΍�<�[�h��<�Ѽ��=�� ��=��.��_O����5����'=n"X=:�b�/�T�o=Fv<&3��p�#�����==��;�3��L'=��e=�o�����X�=|��T];f=
��Շ�(h�;n`N���:�����<0�X�Q%ͻ��<	�|�/6ۼ�c�<×B={"�ld��.�����3䁼���=q=�9<�,=��]��,�<��Z=�o�<j���J�;Ȼ�0�<{ę;�w<�ȵ��F=*(K="��<@9=���x�F=%DV���O�Y	=�}�<�/�<��#=���;c\3�$J�<�����;�e:�i��B�<6�4�I�5:�~=@�:���<9?=���^.=��<Ľڼ�Kg=i�"=���wF��<�^=�:l=����{���:�2<vas<�\=�o<Z�>�S;=�A=�r�ȃ��/N=ms��@V=�I�L��� μ`4<,��<��<�3f���>��㜼�@=9�-�qs,<>���eC=l�:�BaP=�0�<m^���b�;�<ZuԼJ�r=1�t9����<�>�<��=ʳ@=+�7��c�<gt���>u�׉t�.t���q����<nq�W�P�j�^��<�b��Xܼ�V���@=�6�;�O�q�ɼ�=ָ�<�=|�
���b<�܅���=�K����Ҽ��0b���yҼ"��<b��:	�%=��{�*��G�<æ�ٺ�����<�$�;y"=>�<	5	��ϼ��<��Ŗ�	@=��޻��Y�@�3=�_<|�ڼ)��<�U�<i���(H����$=��<�3*=0��<��Z��F]�;�I���=�!�<1_W�L���
�<*Z����<	l�<�E�<��<7k"=,8.<�~1�`'=&Nû���<�;�F9=";=F���=H=�p=��= �<$�#��=��%���,�][�<�~�-4C�dN<ܶ���C=Y���F���,=�f5=�G-=�ݼ�@�=�-�<�=�E_=�Z��?�W=��yR�<-�_=�[�q��<ῼa?�;��=�3��/�H=��3:������=?.K���[=�,=@PX<:�޼.�k<<�\�K�<A�'�̋�<D��<l+���<���<6|��><�꼂�~=��;��=%}'�~lH���T�K=�uK=�� ��!4���x���(��4�S2���E�<�C=�� ��y�%�컠"�;���;p�c���Tx���?=�R\��X0��tW�a:6���c<�,�<T�y�m�)=Z}<E}T���ڼ}�@��&*���^���<=o�἟F�;@��H�&��Z=�t:
{*��K
�&39=��|!K���=��:��V���#=��w;j����h��=?_�</[�<��Ƽ�^��==�	6<��Z=HZ�<���<ғ<+u�<:���F���4e�6��<*ļ:���m�ǵ=�Y =�c�<R��<D���D�6=w}]<\ Q:�U�c�!��|S=�f��U	=%^=�<쭷�!ꤼ�yy��[=�t&��4=�S=C5���ɼk�g�8S���#L��z'=��<�[�<��D�j�F=�u�aP<=���<�?"� �'��\=��&�4�(=}A��r!����;�8�G�<�T�y��MI=<�.=!,6�=�,=�7�<�b]���7<��<��=z�h��F<�s��|;=�F��uͼ����wX��۟<����1��;�ޝ:yѻ���S���ü/m�/l%=�wE��v/��e=�/�Ŵl<�(��q��	6;���.���=Fn$�ɬu�>@3=%�=���2��9�̹(+v��g:�O-�<q=]v	�R�<!ͨ<�w'<<�b=�м�<�bw�*���؀<�%�<Y"K�����%�*�<Gs����/���<�7=��=D1'��0=�BZ���=v6)=� ú�U��<2<���{���f�<��<T�o=YH����=޽&;4܁=��o=��=Z�u<x� ��{=�#��5>=�ȍ=��꼔T��ɛ��@_��y���.V=��<��.<v?.=6c�=	]g=5�=�h��J��n���p�<_LO=3=��V=顼<����Aiq�a�����<5�w���A�\ :��4=Yf���><T��;Q��q�p]s�&��<͵��1<j8ļB<G$�����;�_l�d�Ҽ��<�"=��G=UH=%�<��M�q�<��X;�<>=b�N�Rj<>� �����(�����+�|D���m�E�bOM���=B�=I�<@���GXJ=Qf�<tkK�i�=��;.P�<$�M<=<�;�k����<�׼�.�Ǧ���<��ϼ�\��2O=4B�iN�<v�ջq�Z=�:�]����m<����h�!=|�~;�� �^���
8=��:�]�j��^�;��<��a;V9�:J=�b�i��<� �<JƱ<ժ��=��;y�<��)�;��<���#I�?\�98W=R'-;����a=4��e=�v�<��d�N����<�*��)�Q�)�:<gUc=�8��~K<�?�Z�S=��(�n�:�Gx=N9��$�=��+<AW��k=��Z�V��;:�<��S���1���=�������;f�]=�$,<2B�<���;<"	=q=����u=��k�������˻F�+=��=�-
=��ż���<�o<	�T��
�<7k��<�<S֍=���Cq�耣�#ǯ���h��(]<�T��+Aټ�`��Mׯ�JS��P�[<���<�i�<_��j�=7�==a��=`�	=�W�<81�<�g�XA��켳iH=������=�A�<���I=H�'=LcT�POJ=��G�	��:��񼄥�<+Z ����F�:Úv�3:=.�<��<̤�<*��_�_<Ed�;´<΢_�q�L��=A�=x�,=l5&=����N|=��<ׂ�<1�Ǽ���<�Z=&Ӷ���u=(�<�q����	A;����#�;����Լ�P�<O�d=�(=}\8���<�B�<���<~(=NN=}(�=8�c=� i�OM���_��a�:KhI=^;~=�'2�Y"�����jû�Cm���<��ƺg)�;5KּL�g=򺟱Ӽ-v���TU���s=n ��Ue=��=���5����<��ȼjI*���<%S<�h6=媙;�m�iC���ļ�η��*Ẇ�C<��g��o�<�G��2V�.�������X��W=��I=?��<+�K:ИO��Uk�Se`=Mܵ<�=��%����<�I=��<��
=9�����<	�8=�����vw=f+����<L�<܋B=���<22�C��Cc�<m=Ϲ���:��_=���<Rփ;�o�9ݼ�*�J=	q)���=�i>��������<�lR=�@��8��\��l"i<A>���������i���;��<�y��?��<h�m=Bȼk�@=X�X=0.w<qt׹RT�:t�/�=�����Ͻ�<��;��<�n=�(�;&���0�v�i�e�9=�=�N=pNX���R���f=�e��=v�ʼ��v�.��j=�i&=I���|������D,=�M=m��� R���I=���
)<��<�����F�e�D��sG�K�k=��;��r=PrO=K�x�
�<>=0=�<��I;%�2=y�
=��9��.���v	��y<D����:�m=��Ż�f��>S=��m=?Or��=�������+�W4W�2�=������b<=:o&=!�*����<��T�A��<�et�� :�8Z��O�;K=��~<��A���,<��	�א(<��<aUJ��/=[���	�v;}"k�����e����q�<0ܻP�A��Gp�h3�U�J=r2�#b�<��a=H�G=�<�݁�
�����0� R����ܼA(���i�<��.��A�5�=U�C�q7;��O�8�-ܼ?}�<�#;�����e��}*�ٓj=(��; �<���<9��<-��; <8�����e���8���<�g��i,=n��<�Ӽ��=f2���F=���;�
y<Fa�)�c������mg=%M:� �<�oI=�H�<�I5=�_=?�O�k��=��
��j< 3=g�D=폥<þ�[v=ip�<�j[=Lk=��=��-=�ޣ<�.!<�jW��wx; ئ:��Z�]�]Ѹ<��<7%�;%
����<�U[=�>��!(���e2=�GX=HX�38��b�<#���2�a�8�<��< �;<.Z�w���4�ۍY��k���Լ��q�{�c螻��S�s�d=�aҼ�R0���ּ��<J?�<���ʻU��\o�G�<E6C��>����s���?�<�I���i=X��:Me=;`�<�{V<��!�.憽購¡�߾��E_[<�}�	u���<+�*<�h[�{Ԣ�? *������O=mY��8��<�,ɼ��T=�r����<y�<e�U<��t�����-fx<l�=��;���i�<=��a=�=���<�c���54����#}'��\��<�-�������� ��.�$=�v/����<�h=r�;$����+=�mZ�����������<'=�|¼ZSN���;�8���h'�����/`���ּ��3�O�v;��	��؟����<����bBg���_���<��\��e<kl������P�%S�<<'�0]4�P�G=r��<�+�<�(����b=�[,=��>��8G���6�)Xܼ�C%<�
ļ��G<^��<�&��������<tA	;p���q9�<��i=⣗���`���j �<5HG��d���z�jT˼�
r=؄c<'��;�Fn�h�=ý�ۼ�����;�9º����\�=K����w:=è=1�=��=��<u(���d==q��ͦ��{�O<)0=W(e=�ؼ��<��޼	6N=��~8c��Ɓ�v��Z�<ӌy<�k=˕�=���z"=G�V=M�;+��=a�:=�Ǳ:�?׻{�R�L@˼ݬw�<\]���:³H=�͍<xZ=t�Ѽ�Y=<�<��뼗b���ځ����T��=o�H<-������4*�<����==km/<��v��YR�)�ϼ�s�<���<���<���<-���uG��Z���ʍ�\�̺��<VB�=��Y<�B=�F��� �<"p�_cS��¾;��#�f�!=� m=���<�?�m�>�h�=��K�@_�<�x�<�Q�;-J5������Y=��Z=GUG=��=}o�d	��!�ܩ�<2�⼭��<�R�<P�=��=&Q=�x<�5=9�����"�ZX;Y�U�� =�\���<TS2��85;�s��n=W�q�}����j-��y�����<��K<�5�<	��Oj>��5���k漰��i,�d�����z���T=|�׼5�����<
�S��>�=b�=de��\=*���T�<-�n�H�;�[�F�<��	�!�7�vؼ@���`�^/g�0瑽]j�+I�+>=q �<��<u����w�����=v��+h��
��<h������V�6=��������	缬�5=iKB<�A���=п�;\ފ<i'k=�-'��D=}A�T��;�#3�*!��6�8��*O�W����A���<��6�}j�>�:�!=S����y��=bK��[�<u��O��ûI��<���7�eM=�G�;�o���˼jz�K&=V�=}�<o��!Զ�95=�����ƍ<�#��+���-g��d/=a�C��*�6���xow=B=��<wk�<��{i=2[�}��М���p�<��6�����W���=����9�d;>ܓ�߿��m�]����<�~:5�5���D'D=.�<r�<�	�J�&Bu=ZļH�����g<�ly<{J����2�1�<{^!=:%��	�ɼ���F��lO���&���9��8�Fg�<E�.=�A�<��=��d���<Y�<�U����輾 Z�T�V=8\�`_=z�g=�l��8��<1g���6\=-�׼%�3��}=�Y+���R='�<���;0��<c�b���<]�ûiEz�=*R;�Oa=�]��t��<�A��ح��xJh���=��;�&<Z��;��Z;����׸�<L�<؜����=����T�F;��@�Lx;`����PM=�xf=P6���<�E=�O�b��0A=l�����
�?;H�<E�ȼO����<����4"/�o`='߸�ãH��ڛ<�Ui=8%<s�@�C�<�h_���3�4)]�0h��,9�<�.R�+�(=i�%=$����K8=g�K�8i=-x;��<��
�83��8<��=���,_�;l�r;�0#=��I���o�� Q=vY�:=;�;�C�e2=�U =��D�J�M��<��Z=P��;=�x����� u��d�t������p� =bes=��6��S0=mB,=�
�y8��O��l�y�J=�yf=M���m�	����7�k;��<���;5=}d|���@��I�yMȼ���FӃ<Cg�<LR%=����Zi�<t(�<��μ�E[�=�� <��<�x<���9~�I=`&��5=�c��)�<���9ɺ:*���s���j	�s쁼t�r�<0�n=����z5���˼~�R�~�5���;�wG�<�K��yB&=���;��< x==؜�<[ϼ<F<��N=)Ob�����b����]����G�<v��Q�]���z�֤�+� �bG�<��=j��5���뭼">=��%�+�v���d=�0Z��.��`l=,��;�ɼ�!��oJ���Ǽ��	���=�i�;#$���<��i��(1=~�<Y�&=��=��P<Q<�<���<�|%=�"���7�ׄ7�}g�}�L���<��3=$=���'9������f��=�k;�7�;M���&w� �<5)Z=�5�T�;������:j�<�SG���Uɼ*3]=7��8�q=�Z.�������<k�-���<rK�i>^=�t�<�6d=�����Mf�����DID=o�����:�y��ы�<�������D�5�TI"=��z=���a���g�?�鼞ޭ���(=vG�;��<eB�Ռ���k0�=W)���T�<В���P�<[�ݼX����q=>*=��]���b<���:��4:S =�i{�����`
�<��o;�)S�Ⱦ�<MM��Cu��!W<-L�<x�=��y<�e=H�_��  <d`���d=��]=9�?=�zͼ���Ap���_��=9�(G�� �3�K�`=����ּ��h<���1��<�2'=�Sμ~�꼇�<��z�<LQ���R�<�,�r��;p�0����;6�8��j}=\�<u��<��]=Lw<��Ì�93=����c��5^���=�$�<��3��� ��
�;��<�W�<M�)=x ����#�n�d=�s��?u���\���=}I>��H�5$��K�=��<X7=�����Z��|=�����:=[KE=�Z�jq�<�����_<�`P���;�9��mD=$6.���(=���N�4=-�׼t�6;����ϼ�����<pR�;�|�_A4<��3<�����2�|#�<A�ܩq���ۼ��k=�@���j�V�����=2��#L9�z�������1=����f�<? ����:(��<��`*�<S,ͼA�/=h5=�w�<�܃=vz�$��:�K��u4���J<&�V��s�U�i������X����=��-=��x����.-=J38=$�=�D�<k�@�����ڼ&L�=A��<�L=���:�=��(��F�;�$=��8=(�)<>�=��<�J��D��<�8=�͆=JKJ=�D�+y�<qH�;��x<Ufh��Y�<���<~�G���
��罼	�<��7���<1�yk=�UWh<������1=�.%���e�Jw�<���<*��Iּ���0ob��k�<���q���|<�*=�������<α�ZE��@=�K4= �D�8=>��<YC�����`p<jJ�M(�=�"��7("�<;ѼJ4�<R������ϼ��ּxpV=�1�Is�<��<�A<��";�=�T�K�e<_�={����}��?y<�SN=���c_=
:C=��;�w���<q>��X��p�<v�V���$=w�^�<�H��~=T.=6�G��S%�U=����=J�=�<��8<��;=��A=*�<Cd��۷���b=/4(���2<;�<~�9=�(i<�P�<"��<j�1�mVM��6=$*=6�U�h�����<��'=��n���=i��(#�<؄-=\�=܀�����6I��[c��zݼ������P���ޭ��`c=�8���Ҽ	�r�Z�_=�(�h=�n�$�X�;�1Y=�������.����T��Q!��P}<O�W=^�����^=����|�K����<kƚ� �=�zG=��e=ބ�<�Q=��C:��7�	�=����qx���}���x=q�9���.�� �<<��=����ޡA=:<%���<1 M��<K=���<d8�y?�{m��X�_cA�nD�V �<w\����e���1��1=��Q=��R�Z�<�6�<��d��<�Y=�/<�C&���;��!.�~�(=���;�V=�*	=�j=[�=bs7=޺�eHG��X���%�3�7�YBJ��t+�e��_�9=;��]���5�,=_(��&�y̼��� ��<�ո���b3�<���J~�Y�Y=��< Y2�QF=cH��o!;��3���<W2�u�=��X[��MS��\=5�b�CO]�?	�ۀ/�O�<�|B�C��� �ޘ\=*8=��V=�-�{�|�O9.�f�;0�V�TR)�К+=錟��u�<��<�X�M<h�<J =`O�"�1=����G�:=�[�<)��;�Bt=:? =:�ػwfD�4�����O=n�[�x}��CT�<m�v=E��A�̼[�G�u�5��	`���8=��|=[�$;�s�<��ͼV�ż��8=P�?��7X=$m<b��id���=q����R�i+��Du^=������3=�K#;���O!Z�A���b#=��X<�~�<&_=D�=�齼�����#c<i$o;<L�<r�<�����ھ<�T���/=h�:FE�[��=5?�=8o�5'V=���䯷<}Ќ;
����"=+�5$����<�V�<�g���h�?>"=�#���@��$=���;Ֆ=;�N==O�z�
=�弳,]�I���\���:Fj��l��yU�<?`=P�u��S=��*=������{=�@r����D޼ՓT��t��<��$�=<8 =�ln��>;��A=;�8=��<�ҷ<{�5=<�U=����Af�!0�<�����L<��o<��:)�T=v���xO���6�Ws
=7�=�5r=�tD=��L�J_=n���<=<�&�`L=�J*��X�ľV;2���;!�"q�&{��#�.=m�[�N�]�+�j��F=솽bꅼ�S��7�sA�;��+;�b�A�=�=s��tg=�~�<���jg��Q*��36=9?=;�'<>��Q_���D��Gz�<�ż?:<߻���=.� =Y��G�"��E�����:�<X�=N_��-5��z>��v�<|j6�������<#4��,K<�Չ�l� �8ڂ����9O
��as��Q�X�4�y�u=R��<�Ɓ��br=��<�#�8�<l?�9 9��gM=f/<����<�	�=�W���I9=��M�>���ؼ�����	��=Bn�k;�bU=�=�=4Z=����M�z���Y���ɺ˦�G=�>���#׎������N+���=�� =�H��<�<�u��=��;@��<��p�i�%=A��;Q�Y<2I�<��/<GL׼\�����=[K����*==���0)��,>�Ԩ�<���<�38��ݕ<��<��b�ļ ���֪L��<fm;����z5�k�}��\\�:�V�U0%<��6=��"<4L:=SQ:��@4=P�H=Y�s<'&;�x<���<�@��O� �~=Y�4�]�[<p�=�׼���Q�^���;*�(=�m��8��b�;�a�<<G��v��<�0���\I��n;=�|
���j=	����g=|i=�==��b;�?m��?$<��	��8�<[_=ʠ>�&og;+�����E=�,S=��*��G=�rE= �%�[�<��<���V==�J< ��<=�TF=C��<�	�����	�<����u�N=+jW<�\�
�:��ż�6=f��<B�+=8Fs��=��g<��<�;8=*�,�b��<��%=���Qf��4��W螼�c=h�"=�����ۼDR)=����6�::{��=w�͸}�`��qc�^bk�;L�<��=��˻��=�O-=Z߯;������<��<�
��/=��<=�-�f (=]3~�P���j�\)Q����;���<��ϼK&N��l���F� �x�Sh1��`뻍j=��+=`Y=��=b,�<%��x�F=��\<*�A=K��<�ҫ<& =K��	1=y��;�y=��!]=(�<�=ȼ&�����(���0='�p<~8=V��@��$�<Qϓ;�D��y׼%����l;�Ő<�wZ�(h�;�U=�`W=&�<ԭH�ƅ7=H��:�:��=e�)�^ X����<�nP�}3���{¼Ƅ�0�4��;� E�j�[�;�e���ȼ0�T=�<Y+�]�Լq/j=c� =�Ԥ�e3�<!=x�0='�b�!��9X䭻]�܃�<�
D�J��:�2i<�=����v<��w=��\��Ax=n뼙c��~*D�pݼ��+=���:.��x
c�uq�<���vO=��=g�ͼ��h��T��0h�;x'�<.
�<�ɲ��TѺZ(�_#Z=��&=�����V=�����!=�	�<~�~���;��<'3�<K�*=��J< �:-4ļ��=�-�����.����ü�
!=dQc��)z=�;�<�5 =�/j=�0N����<~�:��9��$=QxY���v=�o"�6sS=bn�:��G����	�B�/�<���:m$F�����Y*�<.�Q=�v�<�<i��<��~��@=p=(�󼖆�(���ƻ�4��
r=[,=�9R��E$=�D��[�<뼍R�o����`ɻd�K=�;=����+H����=�p����A���r��|��l��;㫎������<�=�k��6<2z�<RZG���������#<N��� �!�)=�M= ���49v�ǼC�F;�.�;�4A=�O<=���;��,�)�Z=N����=\:�R=��?=����H=<�S���\��3=�F����<p (=;�mo<כ���]�=��n=�ŉ<��<e�=��4������b�<��:�����<� ͼ{�� ���x�;X�$=��a�5�
�k�;�Z�<�1�]$=g�����:>!м�(I�m����Y�����E����-�,����<x��=0�C��"
=u�=M�<�<���W�\ݖ<�%==��+<��-=��<��Sm=hɺ�=�G%��b�=',����
�ꤑ<�t�������܅<`�*��U�<�u�=��S���f�����deϼ��=��p������<@S�<�����ջ�IT<���<zA�a�E����<�z���B���2=�ԅ<
=�8���=��<�r�<�Հ;фG��5=��=y���X�iN=y#�b�"�*��<� =��1<���q�<�Y�m<G@�%Z��Fv���<˲�<�=c=w���B�x�]='Z�(2�<�9��>p���G����<�r�;�=�&��u�W��[o��?#= ZS�`�<l����A=*輆@漉m�����kؼ�C�<9�	=���v� =�4<=�T="Q�;�Dn=�dX�#)�<f�8<\�Xh�gZR�!P5�|%=��=NU=�9���q<a9��?��L=8m���=�ra�}e�=+�g�+�<�<�Z9K=��E=���:��ż��<�.�<��=�?<Vs><��I;e�)��h=|K;,��<�)=6����B=��<1}S;`ϼ�)�;��E�8����ռ� ����<+R�</1��4<.H=b
[����P6�h��)�<cE.=�#J=�?�����;siF�������MM����;+T��L=��ռ-��<�`�m�<�A����"�����4-@=����he<I6=�K������<��p�H�=*�0=^j>=�}^=9殼�ڔ<C��$MU���=�&S��Do<��B�
�8���ZU#��?����v���")�t�5�L�<��"=	��;s�/�D��<s���p-=�Z�;�~�<��P=�EL�i�=8 d�Ar���꼇¦;��=�i��p=�M�<��B=�\�<�H����<���D^D���[���@�YN=L��<��1<�sf<r����e����j��͸="�?=�!����b�<P9���k�:�3=t�-��V<��@޼cQ*��{�<a�`�b{����9lP<ˋ�D{7=��K�H���X=j�<QRݼ:��<$�=?~�l�(�F�n=�F�<P�2<P�Ҽ���<aU�����B|;\o���<��j;����#=��H��U���P=J�>��� <'�m<�<T�ι9<�B�:��1����<��=<�â��=��*a���'��:�����JT=<S@5<N�<f��;+$�<�E2=�+�:��&<Z�g�(�4��h�w����- =\u��+ͪ�*���l�=��%��<!��p��<�=�ٻټ� ���+K����n<�[�<�;��/�=�;ro6���<,'6=5?<���Ѽ6C=s����ρ��8t�_u�L��"ԏ<���f�:��J�Ȁ����w=9�j���<������=�b�C"$=ښ>������{�I�"=O�D=�L��(z0��56�R��;=a�)[=�����<��<}�&<#�>���&���h��q�|���sRC;��j�����=����V=0�=Yh=3�r;z.�<K	�����Z����xR=�-=c�0�g��;j��<lq6=9zM=��c���I�H�<A̼M�<�P�:ߣD;��Y=�U��a����C=c<�@�<�g=�,���ki=��<�3h���-=f��;#����=+O�=��<y>k�}�L<�5�<l��;,Ȼ��)=�Pv��=o��<rw���-<��]<ť��%\���D�CuB�?9��ʢ<X����b�9���<wE�<��W�EE���y�+=#�D��k����N?�<���<X�&;��F�����i���<�c��?���[����;L����C=I�@���2�L첼}g=G�ἅ�
=A�&�����͈#=�X<������=4���H�+=��.ձ:��9�0�$��<6���Y�� ��<�Eϼ�#��Hu���P�x9<�c����<�n&=�Q><��@=#M�8�0<4�@=��[��$u=�t�6�k��o�;�>�g�?��j��!����Լp;��B�	�(=!=�	��6�<Ӑ;�k$�pt<~q�<;��s!�*!���1=-}�<ģ�<^��<�R<�O|���ͻm��<1b���H&=��;��њ=Yr��z�<��f=U�<��j=^�T�Ʌ;����;j�7�(Ҽv� =��<�sl�ͷ=�m��L�"�Y=�[<m��;�(��S�ڲT���<fT��զr�[=�����'��g���K��<Z+�<�L1�Q=�䂼�Q�LV����;}�1=*�<;�B<��8�{R�<��_��=�8��ء�lO �-�f���%<}?=ʨg<��ϻF!�;*Y=�+M=%Ҝ�x{4=_�;��\=�t˼i�<Zn�^��Ś<i�%�w(༳&\��Q�<��8���<P��;fפ;�<��(=|�h����*+��K@�5��<���.�D=T��;�&�7R�L��<=��<O��<{�w<M�+=/6<g��*>Q�.�ڻ�m�<��<��-=�C$���
=�Z<r/Ƽ�<�+*��[=s�����4=f�(=N驼��h<	[�;6pd��7:<h*=��v;�'�݅<w�U=U<��%���H=�jм^T;���7��2�7׼�X�<]����<F�<�}�;�==?`;Y!w=Idj=�0����<8����Sf��2=�6f<5�B<zX=C����I���I�C���c�a���=9��<ĥ��FL=�y�<Q��&��z��"��</y�<��<�z4:�w=�w������>4�ا�D0O�W�����S(G:�����4=.��; ��<�O�-�Y�VV��od��7��U�#�G=~��9�g����/��u�\?����������TȜ<�B��$6��5���E�;?����<KH�6�=���<�Q�<9),��1]�Z�D�>):���X�D����=�q��U��<IJg�5�%�����V�;;*=�E����;>d;|p	�پ2����<ӆ�:I�R< � =.��N�=�>�<��4=�X1���:\z��(��� <f=��B�<��Gj<�=��=R��<�n;���x<�<�9=pE=i��<L�#=�S=� F<F�C=�� =S�=�ۛw���byl���=��|<��<m/�<��<��=�G=n�z�������<�SX�ў|��. <��=⑟<�ֈ;ēڼS����V�M�<�dʼ�G=rɈ<�߼�p���I����@2���.� ����s�,=oK���:�CY��l�t=��#���<7�K<����H�=����u�_�A;�a��E�=�D�<s�G�9��<�D����J;ġ���k=<c=�/����1�m4�<*�`���U�=Z:%�� �P�e=!��<^�<R�i�ɮ��d�q�0=u�b�!Z�/�=��I���i=��=��r[=��;�!e��s+=��*��o.=<b�=�X��۹޼�82���a;j&��lC�K��;j��Ƽ��f�@����N��H����<�m<Qo =�4	=�A�<�6T=5�<��伉���N=��8=�z=G�<5� =���=,=o=��9=�`�F��;��¼^m:u�� �<�%��m������<M�$�:[=<A^=�q��IO$����<�9�;�d���<mC��䓼���<xV<��點`2����;!��0��0^=��<w ����ܼ��*<T<����� �:�����G�;��Y��*��ޝ2�:��7%=�Id��6r<s&=��H=��'�;�n�M={뷻����������s�sP=�?l=�2=0#��l��b=�K/��H<�u���.��b�ܔļ-"<����"Q=��=X}>��[���M<��=,2�<ǳT��X=�y�<8T,:�U[=��<�N ��=`�%<%5����<G�=q�(�۰1��w�<T�e=�`=1V�;���gP��_*=��R=\����P<Sz{:ٻA=Y�)�A��<W�<	�?<4-<��Q=�If=����u<���(Ʃ�8X<��`��D=�޺����|�L����	�=u��8���p�ڻ���/.ȼ n=��R<?~5�W&��A伊��-�<GG�n�λ��=տ��YD=>�����<�h�<h��>t<E?�`�J��${�sP�<K�`�͹@������H=-�����<��c�j����sg�^����8��>W"=�x-=��ϼUV=��S=L7=�bQ=~���K�=�N���Ļq|!�އe<-�U<`��<�9��ܫj=�@n��~C=ek�����'=:5����N��@@�܂�<�c�;��X��-p��B�<��i�Hn;�E��B�(���98���d�<|�;�@�<��8=f#=.�b���{�k���k=��#<C�!���Y���:_�����2�=�0:�<}��;_U����2��=�uE��`�����{�A?�;S���Qr���J�N�S�T�=��<%�9=᭝�����YD����<7Z�;1��<\~U=d.$=BPd�wz9�@���z�rP�l��70�<�4<�E<��
�<�ʒ�s�=�>��;*��<^3A���ټY �~w(;�w�<�Q��<��=��$=R�ռ��Y=�<�(��2� 9�D��%���VR,=;��TKZ;8����=ǀ=�+�U���X��>@)=q�L=��g��H�<4Y�� �b=�H�~c=<�;|=���=�"=�ż��ļ��L�g���R�I�����7=��{=�����[=A�@q=�����<:���x<��:�*=��>��iZ=�h)�������?���-�!=�s<��=�~���=�<7 �d^�:8��'=pQ�=��R=��ۺU�;���<��c������W����1�'�1O�<�[�<��n=G�<s��:��K�q�F��S�"iK=���<�)=���<�ͼ�==Pۭ��D/��ݥ<�1H���!=�;|��<���ZY���=]���"=�����n?=�'	=�<`�5�B?�<�6=x�<7J%=s�<� �=�؟</]��l2�<��;p�Լh<\J=�����E=��͹g��w�݂y����<~�=����<&�Ӻw�C=*oM��5R�s�����;Dn�<W�-=�5=P�;'2���1�.��0�;R�	=r�@;�D=CK��ͼ#�3�l�ۼK�<��<�p����Ӽuп<� =�~��M=�K=���;�[2���F�O�g<_�I���N=)
��<�<�YE:�f�;{R'���/=��<%�\=,�V=��F���3<���#�F<�Ff��K=�e =��<Z`":ȼ�� :<�K=đ^���������<�l<[�P��m���|K=�97��\=�,��g<)c��|׼0�Q�wK=�P<z<��5<%�[��X=`j%�R*�<�m��**��A� 6����<�4=�	;�X��ھ�<��#=�?\;��a��d�<�9Y�r+%�ٕ�<>0�N�6=A�
=,�»"o���+��Qq��Y����߼`wX�n������;]G=_M���f�sc<D=#��)=K[Y�Cқ��3J�:��q�5^H=��G��\��7�<�ʼp�!�W��<�=�=g�:=hr�K�E=����E¼���<�a8��I%�x�y=��Ƽ�/��� �禼��<P{���<Wm=!Tἑu[�);Լ{`�K�V=Y=���D<�A=P�˼"��<=�<��#�A�lZ=�	<�py�z"C=�	=�_<H�!�2dB=ɭ�<ᚖ<�t���<%4<�_��(=�ͺ<��@��;=?+��N��^H =|	5<�лg�<�Q/�h
��Z:�m�	<N�;9�<��<&L$=�N�<fZ�k5V�����k�������;��O=�Y�<5���A�<��\<zE��-@ʼq���
=S\=2.=��Y=p==E��<��8�x���
E6=�w"<��{	�C4�넽[+��N%=��<��!=��c:ǜV��6=���;�n<װ�h0i<�g$=�t�;۳�< ��Ue����^=��Լ�5����=��~��Lp�^G�ϼ�;������I�(�сü���<u�"�#�a�A�h�+]<Y�=��>=�h=x����2<�.=����C�::A���z)�̿�;���ws;=^�_��sc=}�w��l&=r�������x=v����m��c��*:���^K����<�B�<�P�|O�o�<����i�<����F<|��<�6���嶼[�7=b+V=Mu=Q��[�<8��<�I����=�
�<�;�^׼%vX�y��S��<�'=�@Y��=0<Շ[=\d=�ڼ2�<�ͼL_���
�;˪2�Ǥ�;�Hy�֨����P�H�=�V2�<|��C?�<��X<D3�a���f%=��<�>�=������`��в<����^=��.=ȳ+=�^���=<z�=�I<$���K�ܐ��lU��L7=��Рv:��<���g�#= �=�u��)IN�G���dJ�	�U�������<;HC� ����*���4�� c���<$��<�<�>��$�;Q�9��Ϡ<�L<BcK=US=�v�<��'��X�<��;梃����e��u�;�K��,ڂ<��g�΢�;�Ѽ�_d=�d<�aY��:Ļ	����I������]���A�O(.�cb=,C��I����NG#���T;���H�X<�Č<.&��"+=�b�r���� �&x-=sN�<$c�^<Y�2��<pR���_����<��=J<1�Ż��e=��z<�Q1=�N�:�|b��.=�����
���z<!��<�:
:j�w=�K=�=A�����e=���Y�<�I�<��輪�<V绻0w#=q�\=/���=��I����)�<61�Y��
�;��e=�}��S��唼��<6;��	�<�g�=	�	<
��<z:�<s� <��*�I��C�<8X��3�_�vlt��"<�Z�<��<HK��	��;{�P��]`�ΐ=�P:<4Dd=u@�<�?������4=������x=���<�R�<��ʼ>g��3=g�+�ɏJ=S�ü�Oȼ�^'9̮��JJ=\h��\P=��J=KHy<G
%�rл��;��W+=�X6=@s��s`=e��;�dt<��Ӽ�O�<X�M���=��b=bBe=@0:=22��#c���;X���`K=<�Ƽ%���� /�S� ��f�r*%=�,<�1A=�������<8y%�\��b��=�$=o�k��mo=�Pn=e�P=fj=��=��A=����<XZ#=���<����:?.�����Gb=Z6�<�Nf�
�D=u�v�H�V���=7�M��M�tݹ��\�<Z��*�i.[��
8��>�ƣ=1���r<��];p-h���<ɥ���C�<;s���μ��<����2=�6���;���d�|BN<�e��\�D����<`�;�Y�F_$�E'Q;4Ys<��@���<��G<lKj<�hv�2�R=�����^e��[�<����Ӽ�(���B <'���K�ܼ[�����<��<�'=�� ��
<^ȼ�z�b��:�	���ޘ��m�;��"<Y��=�s=�̼5�=v�?=T��<@�L�ԧ�=��;�׏<ǆ=J�*=��=�,<p�"=�O2��B7K�^��e�;��<�7M�\:9���=βa���;���=�3�인<T�ʼ�<��<��;�ހ�jO'�����J<�3Լu��N(��@õ�U��<ȉ��~R�=u��<n��c��i�I�=��)�a�Tj)���<��<`�<�F �8��2IB=x���@2��+�<P�= ���
P�o�=w0�<�5��~�Jn'��g0<�@�<jڂ���3�8�<��U<����F̚������j���)��V;D�/=��<}�I�
�컜�=��|<)�Y;�8<52_�>�s<F�'\a=I��<Є��9�����o{��<o�I���q<'�<�'"=�m �2�=�B�;qT5=�"h=��0��?�<d9�A����[Y9-G�A�r=j�>=�L����3=�˕�_��=�p�<3�\��]=�,�ٜ�<Q��<>�@��	^����<��<�����y=6�<��S=G	Ǽ/X���O"<h�û��;Wx�e�ʼ��ɼ-�Y;j�N=T��U��<���<��<�x���-���<�k���=�YU=��<d��<F\��3U��<��<F�V�V��j�`M��3��/=r-�<�պ�f��<L���3�'������2��Z��F�Y�ȼk������l��2�ߎ�<�=(=���<2u/=95<S�;�C89�͆���G�4&�<
_=q�==f�+��P(=�2=�4=(�!=D
i��	�ឧ:�{=��V�Yϝ<TX=O�<���<{��ؙ��� ��ހ;��<�\����8��sݼ_���q ��ǭ;X̻C^�<U�;�!��0�<�᫼��	=qB<�-���\����<��Ӽ�*6�;�����;�(��T��2�;|����%<�/=�<V9μ��'=\ߊ��l��u�
��a����P=�$<�)j��O-=!�=o�|<�� =�0�C� �I�I�ߝ������~zS=S�O=J��:.�{���u�;��<�:���"���(=F�8=�Y=-$o�~�����=��3=8�<�P>��S0;��S=7]=��<2�Ѽ~�ɼ��A;Y�G����;�𓼹q����>�qA=�u3=�7���;������P�d��:���<�����<R�����0=�L%�Ȋ����PWT<�[���u���/�ş�<A��=��@=�a=�}��+�;=p�W=c9��Ö<Ak���W�㻏L=�`����,<]�<1�S����<V�<�*u=b��<ټz��$=����p=֞<��ݼ����x���V��)q"=��=��<��N=f�P���ԣv�_��6��P��o���iM��Y�<�-<�I��|������#���G�D]�<0F��`�<_c��"��;�=5�/=��2�b<�"�V�=��z�:�0<����o�=�tt<��<2=Q����=%�����H=G�4<�-�<�<=Xh<ė/��(��ju=��<���<Z���J�l:4:2���;��.=��)b=��;#�ż���<q�U;,Qx��uS�T"<��<��<I����9����;{���U=���j=~�|��%U=t5=�u���< gո#=S�p�;
м��D�C%=���X==>=v����m�;���;�x���I��6ۼR���1�p�=��<=V~=���<T���
��z�<th����<��8=¼T�B���<�E��;ND]�	�4=�o+=_��<hH/=x��<L�4��ў��1=�^O� Tb���<믂���D=�SD�%!<����v�<*Y<Χ'=��+x6=إ1=�\=T}=
���&�����<��k�;*�+�ڻ��z���:���=��<��ݼb�]��+=}�=="�=�u=M�<�?�<Ɤ=s���^`=ډ6�g8,<�6< �+��-��=�=x�<�&��<6 �<Π�=�
#<�� =7O?���;��v������<�*=�|�<��=!�>=�C<8v<�A��
�˫׼�A��J�R+=�r=U�8=H��$�};�g��E=/3D��=��u�dLA=!�\w�!G��F�|��=5�{=nBӼ5�K��#<h������� ��l<����+�z=%"+=�o��M<0�=�#a:yA���1��&�d�C�n�V=[8=�3�;��缡�3=ZQ
=�#<�9]=����k0=D�]��n��N=�$ټ���<)�&�6�!�D��:1al<U�<��E�Q����Gⶼ�{|<�	��y�<�
=��*���W/9<�����N=����ǾQ=8�¼/(=���<h:�<vv <9�̻�}�y��<�#�;���;��s=���<�\'�Cֵ<"=�;c�C;8l���]�<�e=�Ǜ<N!=E/��<��hD�<�ɔ<Zq�ͧ�"�ּ��<��=�/�H�sPV�� =K�&��P�<#9���7<�~*�|��r-[=|�W=j�&=�>���+=X�9�JZT��J;<�X󼊔��GI>�%����&���2��Z8�wUr��������R��0=��U�[_;��%�B/=��3=�<>=�9=�'5=]_)=�@�pH�<��<su&����<���<r�'=�yq��7μ���������`<,��b =,=8?7<�=rg_=�,�?�=�'���
��BI��<=��<�R���a=�U�ow
�����<��[�=������c#���� ���=$9^���ԖH�Z����<4�;6�A=}A#��6��N<�u=���)��:s��<4�x�8# �����C�o���=�V��b/u<����GY�dd0=X�<���<[�=� ���;	7ļKuU�������{�㔂=P~=��9�}0�;��B��z{b;f������g��j�B.x��@&=μ���}�WJ�<�c�O���7;���<�(������b��< F�<>��M@d=�����!���.��f=��X��3�.Z���O��0����:���{H��l=s��<�n��Ђ��2�<���;�iX�p����k�����.=��,=?����'=�,��<A@92�\=L|O=�=88R=��f��)���ie=���<6�^:���<H��<w=�����"�=;�<q�Q�C�s<�z��Ö��f�a�`���7]=6-���=�`A=�n��b���tc|=�w�<��3=Q�d��s�9Tls=�)=`�(:��a��F��́��pڻ��I��=[K�֐O=�;D�r�p=���<���<R����&<�Pk��u<~P˼�M/=ee=�+�����|/=BR>=���E�%=�_���r=�j�<��q� �3=vwƼt^ּ�z�`�"��	`=s*=��a;�ώ��4�<fP=%�ƴ\=�8-<B�=�� ={�;���ڼ,JZ�|�A:δ:�O��	���aH;���Cɖ<|Bm<9�<h˼v�<wj�J �X�U=O�E=1K[�E[;��(=����KI=얏=r��5�ʺ�g<	��p�<��<~��<��:�!�<\B�7�=�k�*�<�,���j���Pj��n<�e�C*��=�=�<Hz�;F�������hB=esi� ��:]�~<�p���'=q�Z<��g�f��<������!=u&����<5\�<��<��=�P���&����9�S�D)���n��#Ik�$|L�,l�2���K4=��5�/�X<��Q�A��J�=$od��9y�T�=�ۡ��A�8{�_<��$�����Fm�o�;���<M�D�b-=4!�:1:���S��9�����<�B<��1�/�R��Ѽоp8J7?�l<���</�ȼg샼������l;k��M�=h�ּa�y<�j����Q*X�"�;f�=��A���
=U������:F+=D�\=@�F��pf=Н8��Y��A��K��C��<&����<um��ӕ;�o�<���ָ��ji�+1=
�Q='	R��H��ze�鸰��X<X�7����&��<�&�<�x����k�:�W=�j������;�b̼��<5�=Fh��b-$=HՉ<��?=A��]�n=��H=��S=/�<��I��N�Un�d``�ٴ��FTX�� ��XC��@�>��<�
���l�Q���.7�ˁ@�<�*��h�L�ͼ�1�:q�:[�*;��;𝷼���<�Pn�DF�2��Ûع�A�<��=�(<L��<DY"=�SG�;�g=Z,��� � 1�0.<���<�D=۠<��T��X�/�;��E��T�=� ����"*�]�h��ZI<�籼mB=Iq=�K���G=~$=`���������<6�t����<��}��m:�[+�0He����<�1<�H����x�Ƽ!;�<����I =�U ����<�';���q�I=����=0;u=�m׼ FK=�s<c�g=t�F�.V=Zؗ<�P<+�]�H��<)�K���<q��<<�|<G�K���<�2;�iD<9��d��b��l=�J���|�<���<N�n=�l�<�%<���;�j\=�Y=�M�<}����<=�8��Ƨ�=�<uC+=v�U���5=x�+��(=�!�f�Q=.Xn=A\==�\���Q�SZ=���_���;`�B�8�_���>� M�Q!g���1�>�]=�{w=�n�io���<�|<���<ʉ�<'#���N(���=��<�dW�.�̼�	=��t�;n;�0Q<i�<�߼��#�-=��>=ޒ	���Լ1��:4t�<@�G;��=�Z��u�}B�<�����=��t�&λ}ּ�Vw<�? �d��<�M輯()��Z=�`�<'���8���$W�8M1��U2=��ܻ�2�<`��BM��t�"}�<�j=�����<��e=J=��<&pr�K��ǖ�<�A��}Ȼ�^:=��8<%]�;���<��V=&OO=�<@=뾻��𚼧�F��R)�BC�<cM�<��༧2j=`Fd��AP������Nu=�J<�v(=6,=�8%�>����<�r1<�|�<�~ü�A=^�h=7#]�Y���Y�<\�����{���G�Vȴ<�0�K��57=��޼V���
�c=Cּ�F/=��E�B3�#�=b��Y�[=���;G��t�N�"�|����<
�<J�X��=�=����p<�̵9�q˼,Ɉ=�����<��o;����p2q<pv<��&=���=w�U=�?�<���؁V=�k���꺈zg<L�Y;�4=J{Ӽ����s�;�<��=�ܶ<�l#=��<&��9b�`��7W�V��<J�X�"։<��<��;w7�<��$�*� =y=��b(=	���t2�r�B�J1=G��f�s�N_�9so��� �1�v<�*?=�Y=^�ἓ�<&�=�^�_;�C�<�`E=�0��$5�<�̒�ma��;�鿺|c��&�z=�&T<"_�<
U�����<�����b�r=��<���p=��[=�=<�>3<ɉ�̳���s�����%μ��*=ў`=S^=��V:_�����<�	Ļ��;�Qb<l�<��;�"	�BG켶��w�7=M𺃲 �^�g<��<;�=q����<'G=��==��S=�Qʻ|'��pvZ:��,=%k,=�<��R�G�<��;�?);����B��'=��.=ax<V��<V�=e��<c<=X�Q<�ü(\��4����:��/�o����<r/c���?��]��0��i�O�/.>�WRü��޼�q)=8�+�2�<����<bO�<d'={&<3�������=�A=���;��W=&�I���=Hdռn��<�� �=&P=	�ü��"=	N��4Ѽ�n[�@�����'�B��=�E�X�p=�$,�U�p<�7��D8-���k�!��e��'a=�Q����"<�
��+��&�g</�E�������%=�����a=8�e=�`=m��H=BJ(�Y`<l1��p^� ��Ɛ#<D^�4�D�!<��� G=�
-;�ɩ<[7�Џ@=���<_���0<�M4�dx���Ӽ��5���A=ۥ%=M0=�Mܼ({�<�j�<����������ּ;H=��Y=�u=�j=��*=�֏<EC6=��������L似3��A5�:r'G=zB�<��C� DP=��r�G�*��<�@�<j�
��@_=�FK=�NI�\�ؼ���d��<��c�d��9��̻��
�1�'�5CJ=��<���<j�M���o�/d��/=2�=�s\�,H1���#=�˱<(��:�5�<�c���[)=��0�r���<�_���!�������J=�4B=w?ټ�Ǉ�0 꼤3�:I�;�9ؼxZ>���=�J�<w�a<���5Q�<#TH��`�<V��:#�==� Z�rLB=m6�<���Jk�o�U=�s=A�=pY�5���8kQ=��|�2�1�z�%=ڽV=��q���Y�Z�5�Z�8�vU7��G��h$=�T�4Q�\Iz<hf
�Y]��nC�}ܼu�R��@*��c}=�6�<�l�wuc��<�gO<����7��M��T¼߻�m�<ra�[Զ�^�+=!&�<!4<Kz�<��O70�\���϶;����4�4=�$��6<�3�<���;W��<ǑP�\�e=u[>=�En=�ց<��\=���m@/���C�x +�*�	�2��!�r=%��n��(c7=���;��=��<wX=-:&=�2<+��<���:R�d��h=�Z= ���'���*1�~U�<`[5<�܎�A���W	S��D��ñ[=���<E"ݼ�T���������<�f��w?��LJ=�>�<�
�;}�
=|��;�y^�7�.=K'==�\<#��<b���&[�a
��7� pἜ�R���n��g�<i���]�n���)=<)=Cض< h�<���ޠ��v�o���G=��7=�Ճ<]ǧ��1�=�!���3=���<q�<M�7=~a=N=\����;=�a��C�Q=̹�m�����<z/�����;2	;i*P=�[ҼD<�5>�j׻��h����^���.��U=�v8���~=��j=���<�>�;Le�<
˄�i��d>����4�0�=�����*�jD^������:��|��3,��ͳK��H=U=x�<��T=\��:�	=x�N�w�M�k?[��<���'�g�#<d#;��ټ�A=lO=��</j�="B =O[�/�<ޓ��~S=�KD�tr���<�F���Ų��<�<�U�����<��7=G�r�z�%< =�� =2�:�R<��J�)��<��<M�E<jL��=N�=U=~�m���7=�	Z<PQ�<�n��8G:;LC��O��3����(S����:y��<�I��1!�B�6�A:̼$J3�tS=L����[;)<e��m�|��]=Jh=)l=��ռ�`6=4�b��I=U���=`�="�K=d�K<�?=Fɒ����<lnW=�7�;��ȼ��?=I
P=�bA� 0g��<(=ˉv=ُ��\Y=�%�<8Z
=ô�<�ݓ��^�<d=�[����<e��<x=�*:��#R=�&8���A�������<��<�v�<&FC=$��_�<O� =HC=0k=g��C�R=�Jp<m�<���(j=�d=�C�=@��;�4Z��3ּ��?=�2=@<N=�����߻E®<�N�^Up=霈<5i�<�XI<F�.�<�`<	W<�G%�;ZK�9��:�,�;(�;�0=64���a�X�R=� ׼M'=���<�ff<���<�;�<k��b�=�j=:���[q=���<��<�}ּ��vI;!�Q�H�6���<�j�</�";r�<pヽu'<��r�R0����a�{�-�i�=�����lj<���<a
<b�<CV�����U�;u�ޑ�>��<Kc�����<��=Z��\�<�!<bA+�kf�<��<� 1�\;q<Ɯ.�h�<>�e=��R�ˉV=�ى<�Q[����<��f���ڼl�B�d���[�<e��<"i~<�L��.���p���*��*+=g'4��)����@�;):6=݆=aSb=��ʼ�M<?�2<���c��7�-;��";=�/3�$�<�-l=8��ټdlt��"���:f5��Ij?=<�c=�G������� 9��?�<�����V7�u/b���V<f��<iS=��=ё�;�� <�<��>�==�4:}:��^�E��
=�?R� s��s�<�u��=YC=�K��QB=��7�.Y��Cc�r�=�zD=ĕ���4?��N����<�5 ��k�Z��ɹ���B8<�/=0��<w''���t�� F���=��F<���
��.��<���;Ú<~;l=��C*<T�=f�-�
v$=��=�d�#=�3�=�\=
�==����%�<В�<�=>f�����<>89���F<F1%����tV3��#A<96�<��e��k��6�;�쀻�6k���༨�@�5�Y����<�f=��8�n�{=�������<�G�=�R\�]$r=�fź�g'=&�W=�"�<����,���/R�[*G<ev�E��겻�s�<�>W=��=��.�S�p�S��M�P=}�e=���G�Y��[�;X��<N�5=C�D�x��XE�<�p�<� �<��<�2'�lU=�H4K��M�<"H�ĸ���v=��+��5��R��<{:9=�J=��1�0�1���V=�ŉA��ڢ�����q��
�:�[g����<�=�<�����6�����<��K�������<7�?���(<g&"��	��W�:�~M�%��X�<�i�<H6(��'�"�U=&�J��ռT�P�}Q�:�l���N�t� =L��<�����1g=�FD=q���%����d�J�s|���;=څ�<��<���z�<�s"�G��q��+�g�<��4<�p<ȱ=ʁ<H�<��I=!�V;@�x=��ļ���<�5=���x���<�}�Ev��ɺ�6<�Xp;�ʴ<t?<7)���8I��u<w�g�O<�^<p��<��1=��<SY����N=�k=��8�A⮼�l:�弰���>Q=�f|=�[4=Ү3=۸(��f=y7�.9��^�=?ð�Hg��n�/=x2�;���<�I��[�!W=�,��*Y���7�$�8�`�:�1<RF=j~.=�E���ռ�H`�xv���+$����l��<�_��+�<0x=[�1�ht<D(<<oH��U�<�.=g��>���Ι�<���<ģ�<�B����SW�;Th��P����oE���N=	7���[��8��<�3=e������\l=�LZ=����}��2�����<�Z<!�O=>�ͻ�k3��x���3_<#Ik�rSf<�[t�~�'��a��B�81��:�?����0U�;JO�<>��������U�ļ���R=h��<��=�p=���|Y�;=Fx=ӶR<��������ˣx�W��<s@=�5�<V�H=v6�ٞ�:xZ'���=�*���o�<�"�X'=D@�EO������x�=(���}=/�:<y-�<��%��N�<~��=iʼ�Q@<�k�7���f��͏<A�<^0"�;�p�N6=y=kk��c�Ǽ#i�<	e���8V<�2#��x���=ۀ7�ʕ���E/=�/;��m=���<�Y��%ռ�0Y=.(��
=��<&
�<@��<h>���>�l�_�M�[=�~J<�s�=�{!=r�3��߼��@.��#��㉀���G�'�м�D)=ty=�Z*�P���=���e8���=��,=����Ĩ�~�};�yͼg:�<�o�ꪻΈR��(l;�σ����<����ٍ��:ļ���lGE��=Sp ��X=�P<��s)=Jv<�@��ȼ�ѕ;�,�9�\=]X4�iA5�����71�������9="�U��<�6)���e�\e�<R�#�q9��<�;Ţ�<w�l�� �Um.=��;{Ŀ<��3yڼ)��<<��;/=�u�?S�=��&=y�B=��p����<4җ<W�����T���μ�˦�+�3=���<�z���1+�;	H��CB:���-��j4=p������<~��<��$;�)m<�T1=�e�<E��<�?]<�:<<�!<�JC�	~�P�˻�^��;[!<�?�=SC;` �<�k�<3V==�F��n89gv���Լ\��<X;�<=*�<4�=[A�<n=f5�'�-=Se���=���=Æ��+=�q �y޼|��{��)%=:�	=�ݟ<K#=L�����?����y�5<�d��D���Q�υt=@�g:���:�Jc=�+p�*ʼ���<=�v<s�$�R����<�C����̦="h@<��E=6�[=`�t<��c��D���?=τ��ڛ�<5�0���8�A����Y�M��<�r��Ɋf�r^.=*�%=*�=ǫC�&zc��<��;O��|:=�JD��S=��?�0���w�;	12����؛���a%<�)��1�<��y��2�gb=Y*�<����v`=/A#<;�=�;�<Q��QM�;>��n=�g�;��G��ü�lT��a���I���B=��'��%<X!�<w�������0�;��p�ZH2�بq=�7�:S0<=*!�u�}����;�A�8Rk:���<)0��Yq���z:.�V���z�]=&�^=�x=�0=�6N=��i�a����<ʛH=�ڜ��y-��І;K0��t�;Yu=�=�k=/��x��;���� �
�i�,��uܻ���q�O=]^�,�U=n�	�RW�F���S�<2p>�xm޻�-O=�xN=���;�L$;c`%�f�:��<l<����*�A�*=��=Y�,<H+{=E�b��`㻃�=��Q�j\��ZBF=�����ż���<�T�<CÐ��k�;�^������=�"u���`�gϱ<��V<C�=�p�NRu�׈,;��R=?����"��a�+�1l�< ��<:��qT�r�/=["��ʭ<w�?=�g"<�3$=� �<!��n�h=YG�b�d<5r�o�y�Ara=�g1���=�3k���=<1=�f�W�3�݃	<4+��	�<��t=�0�'À��Q�<m�"=�w�hu�<��<�i�<W�=����tۼ�b6��}7��>�⼹7=�HE=z:n��%��YjںN���}�-=O�u�O���(��,=Հ|�0�<�1=����[a=V�Q
�<��k=^w�4�<X�`���t=�=h� ���(<Z��<,|�<wDx�pػ� ��cJ�P��<5�<QR�<�����A)��}vK���������������=��L=0Q$=����.~=ut�(����-,=�0<���'J�==����<��h=���l�G<�2��Ta?;S
=�\����E=|?��;ʼ��)�A�;Vń;͒�<s,=f=5=�iջ.p(=��x<Yf�_ ��L��7׼��g����9���<v�&=��<*�8%H=J���^�<�1�<ly�;=>�;MT��~E��f.һ/�>=������©��4=�cG=W+=��=�9�r�˼uqͼ6�=q;xl{�P�޼~z�<�˻Z�j��yH�6	����J�M!<��<�Ȁ�|�=�L;	���j���H=i�<Kg�� R�<�����3<I�\��%Wh<���t]��*f��"�;�%ļÇ"<��<����Y:;^�<0�D��Z<��<��7��Y=�Q
�I�5=	/j����ո�r�h���	�T�<TN=�fE����ż{��;���<G3�;��_����<��<R	 �X�<��-=/?���\ܻ�xM<T��d��9S��pܼz�[��Kf�F�<���;���G a=4�2=��K�nl���9���1żM�ܻ�D ;Ov���'D=BP+�;'(==T»8�<�v��w��<W�=lWa<����-=�e<V�d�I���eM<����!�x��ӣ��C���|<w������<�>�<C(2=���0�R����TJ�/@C�-��P����J���kм!7���==�n�<��D=$�����=�������"�R<ԃS���L=�){�`�,;V�<��z��Q�����nS(��Q;]��{���T�<�����;>���b� =8R@�9[�m�O�cMȼ �<���;���< �>=���]�<�)��=`��|f=������;�;k�
=��F=��d�B�=�e�<�Um<��,=��f� ����<(��[N���臼l�>�Y=��;��u<�+޼OB,�c�;=�xP=��3=��#:��<�/A���W=�?�;.M<�����ɼK��<�`�(�`��������q��i�@;)�=8u�<�<����#<�kݾ<�Y����=�����=�rG�"��;ߚd<�49=�K==���<�6��E�]<�� ����U�:�½V=��<���<����(E�l1S�%�2�C�h�3�c��y��FƼ�'��i~=��+�@�=%=��7��/�F=��*=\b�<��d=��⻮���eE��1<%C�<���<��t���T;�'����&�ؼ5��=�G��.�:֚�D	���/���F=%"2=}�[= �0=txM=Q���}�����K�a=�{)=�1���<�Ғ����=P���{<�A�U��<���=_мm�=�e6���<�U�����=jtf�_�>��!�s�	��p=��Q=N��<�G��y뼗��<�P�A=A�=�ۻ<s[,��|=��	\��t�٨ͼ�V�<�	a�k���@�C:=�9=�/=�4X=0:V<��}=z���@�<)N!�;-��<�l<Yյ<-�D�˳K���<&�R�N�=.��<�h�<�6}<���<�6 =?�=�A��(A=��=��K<���<��ǻA�7=a`=����ޣ;i(��#=;�L=<o<��D�;���<�:�������<��Z<,���4<m=LX<W�;;�~��N�T=6�=��������3W���(Y��Y�<"L�<s�-=���`�/�cc��?����=T^%��۬<��L�*<��$���<�SY9�g<�7:�w�ݼ�������^�%�J����ߤ�r�����<(Mi=	�<�v�<���<܄���������;v绨5/=#�);�����"=�<�qx���S=�Z�<�|1��Ζ<���O [�B�T=p)�gsI=��^<I��<V\=)~]�?� <HY���K�=|`=+�6�P��<�<.����i#���@��i�<m�����:�P=�(���;�/��x7=��M=b�{���47�<Re�ka<�Õf�V�<�˿���<�)����<V=	J[�	߲���Ӽ-.Y�t���;*c�;�s��)��=ݐ�<}�	=QPp��Ƀ=���+<�)��a2<=��-�������U><����f�<t�Q<��=r�<K��'�V�r׏<G=����<��R=�|�xi׼��ۻ�B��RH����H�<�E�;�Zx<N^(<��A=����va4=?�j;���t�x������ӼL�<��<d��=�x%=��}��~^�׍=i	S�^>��㛴<k�<=;�e=i�<@�A��%=�G5�ɧ���W�<�5�qm?��Y�<�qT�Q�d=&X�<3z����7����'�=�N<B�4��#�<���Z+�A��ث%��l=2�Q=z�h<R �9�h���/��RԻ���30C=��P�Wsݼp���ڼ��ʼ������<���.^<+輑��;�݉;�).=��<����6=waX=ގ[�&����B=F&=�Ƞ�Gr��7P<��;��<��D�Hc�<I�]<h0J=b���:����o�<��5=5k�������m�{$�f��<L(=D�޼|x<U��=/]�<��<.�ysj=��w=[r=7�h��<�)�<�9�<���<Qw,����<��>�cX
����<1v��N��;�Q��a=!E�r�b�0��<'_;�P�<�)3��v)���<n� ;��˻��L3�<ڵx<�y�<�#��n+<e�<[���|�"��%�8=�E@=!9<��s<V�O<el<�=m<=��<�%�q�<!�,��O?��x`���һ��<S�z���,���<���;�̼�!j<-1>��Ą<�ۚ<Mrf���(=��(��iI��"=�@@�0�}��!&��/�ܥ�;3_���X�<]�����$=�ʰ�%d�Lf�k�#�� ѻ&YT�!����  ����<��W᤼C����=���<1K��KD<;_�ȭ><�E���/;`d�E�H��BQ���#;��E��[G���W:��<A:P=�g}�I{{����q�ۼu<F=�H=e�	SJ=���[e��}pX���H�<�V=�L�����<A�\=L��<�b��-�)<a�#�>�C�w��;�x=��<^+�"��<�ϼ*GG�oq�<*�м6E���*=V�<KK:�����J꼏�i�M���R�@���D����"=1�<�|<�̰��C�<kF�����U⠼�%�B;=���(U�Ղ<�6z�Hl�k(�:��e؃�ͥ1�k|���&�8A�<%Xz����V j=-�O�k^��y<�� ��I)�B�Y�U1W=���<~�8���ou�Z�Q=0D=dNJ=}�:
����gF�<��x���<�M��,=�'��]�<I��<�H�<�.�<�*���ؼi���H�w<��8��`=8a;���9��� xc;n��<jC��|�<8�=`����b8��4b=s�Z�M魼��^<XR+<v-�:!)Y�k��<oa�5Zu����<u�&<T�"`���z9���C�=H%n=@4�<���qJE<�����7�x��>Z�$��;�(��[=��=�I=rt��	8׼��^<�[��ޚd=|ܡ�#�<�(˼��<.Έ�fJK��O�<�>@=��<�e!=��A޼rl6=^*���vм�����<��l�S�8�N�a纻�E =���r�=�=����R�����<A�:�:;
`�<�U��B=�4�<jL=*�\���%=_,�<>���T=l�9R�O=a�����[=�!�=Jx����i���ɲ=H��1�=: �9mg;PkY=�ݎ��f%=��B��Q9<f�D��j�<����F<��<|Wü�F�:�r=���<=2(�O�g=��<ݡ�;k�K=]�U=ȲM�Yx��W�yh�;��h�Τ<H]ݼw,���<��V���V=#̓8�|*��j=�ް<1p�k��<f6V<!�<��㼴�<"=���<h�l=�X���Zd�˹k��M��G�<;a�ż ��:�#=Af���C=�<\=tY�<�/�<��={P�9A�x��C�<���jļ��-=�c9=͙=�Q���f���k�
�����B�Fy-=�p=^�t<w۱<��)=Z����'X=Q����]��.= �h���=!�R��:X�3/=�����:""=uc�<�:;A<=$߻J�=4�;�{�;S6=��;M$�<��<Ok׼�)�<��:���<5r<fY�<���/�<�Q6��޸��p�ib�<������	<���2�<���?D2=6�$��!� 2=��ż��M��g;=�*o=�/ �k�s�k���1=4J�;�i��Yv<۪� ����T<#�;=�A�H��<[�g��rF=�.w��c�;o_=kn�ނ�;-�-=� 6=&�R�U�;<.�+=��<��'��6=]6X=p��;�V��Z��<���@�D� =n;�}<<g��L�]=�$Q������=�8z��.Q=��_=-��;��a��W��z
>=9g���ˠ;����}�k�1�)�;��U<*P�:8�W=��V�C�����b��:�����?�H5�<# ����t<[�V��<���]O����O/=C^3�9R��5�D=�-����0;T�I����R<��U�օ�T�L�.O��e=���<�qi�#�I��n�<�h=-3�;���-z���wX=���<�� =�Tt;C=�a�_�[<6��;5��<���ji�w��<+��&T�<e��<r��<H�����n�=nO<�L&�_��"=k`�=�\=�#L=�%V�6��~���lQY<�yY��W�<�����L=��=�#=K����ߤ�<�`�;�&3��8x�?� =?#t=�4�8 ϼ���<�8=�d+<s�;�|.=�,b���<�d ���(=&�j=� �;s�>�ۛ$=�b$=�m2=kV=΁<A�������:�V�M��"=�e]=�A��=j�l�x<bu<��t���K���<,|\�
Ku=pB�+=�<����w$<�bW��R�;}�{��<�绻)���]=��.�b�=M��̛)=+�<�Ө�J�~���"����u�(=6�� ��U`x;�?�<AW�<N�ar�<��<��I��E=��<!w)�{�<�򥼇�����l�����e�h=2ᨼB^�R;n�һ�ܻ��%�m��;��=�`�:���R=S~��j�< ����?��Eq<�T;�^A=E|=5	�<�!�<j��<�伵�T�"�-=bu`��ݗ�Ӌ�ѩ`=y������`�?<6=�֣�|ұ�R8<:��<`�8=�:��G儽Cu<�N�b�={��<�)ʼC	=z�=9�<�%`�r��>�<PW����	��	c�rF�<j����;Q<�H=�P��`<
H8�����p���3�;J@W�����a��Fk�<�d�<��\<�1���˼h�u����<�揺���<���<Q�<sm�<T�[=<�:5�\�ڮm=�_X�i��;�k=/=?�T={���W%�<G�;�W��'����<j<<dKW=N7=DT;��<lIk�����O�㼓��=?��=�I�Q4.�Ͱ�9N�A=&�<|K�<S���V�<���<�"�;K��<+�v=냏���滾�Լɚ=i�����f=TD���e?��Z	�V�*=�za��/=�� ���$�Q��<aa<o���٦��ޞ���<��4=�e5� = �;=��}��y��ďW�'ZF=�X�<]rk��Җ�]����ļ��P�	J��a�<�I9=�a:���D=��;�ga<�|#=4ܕ<b�1=Ӗ~=M�����;rB<U�s=�=��D=II��e=J�E�^FU��0==�w.��C1=,z�:̘D=�8=)us=K筻�58�ak:��$<,��A�v�z�Ѽ�*�=�-��,��<*2=��<��̼�bܻ�=�1=�����C�;�`G��a�<N�=�#��c�8n���Ƨr=�a;�q �����<��%=l+H=���;Ҳa=�)s���K<�$=H������mD=��\�3_<�y}ϼu|�	u����{�E;�\��#<��W=�80���<@|Z�T�&=i{���<K�<��:�s��SX	=�J<%@�#�<�nE�_����=��R�\���
/z�1v�'�<y"��2J=a�^��e�l�>�b=���"=���<`Ğ�֗�+8=���<��<L�<���L��<Zd=����=�켿1�K��<(�E=��.��=K�K��ط���3��뒻#':�CIi�[�=�ϩ<�Վ�R;�;��.<;Vż��)=��}g����漳O�yg���.Y=_:���<��<4l�;����F�<�e�<��[J�u�p<��H���=�2]=�=�r
��u�BX�<	 =�<�j=s��<?�%=򬆼��e=�=��]<L��<3�<�V;��xH=]��<���<̔m�1�"�b@=�3��5�	=�:=���<��g=���<G��ߜ�<	h~<�	����<���<�7�:ks&=��Q������;�;jd"�eܡ�Ĳ���PJ<��:@a�<�^μX=��i5��'m<�X;�C�<��6=��;
�<I�'=M< �%��ij�k�ػ>�=$�<�?c���=�]�����77=�&����<�s�K�<<0����<Eư<��\��*G=��D<(IM�
�Y��IX=$}L�+�)=�R=	�p��P=���b�:m�=]4<=�Mj;�e���3�;f�=���/�#A;��8��oy<p岼�tk��<Џ=M<ʼ��U�V���"�+K\=u\E<�(,=��f�A=?��O�	;��N�bļQ�;n�bf#=n�ּ'���!���a��b=��D����3�<���<S�x���X=��Ļk�w���)��l=���#h4<�FZ=�d=�2=hsN��򼊑�=���1��ZR��O���� �V���z�;R���uT=�ډ;G�,<���<�46=�Y=�Y!�S������;�U=?��<���<1ˮ<Y���8�<�N<MjC�����\=�q&=U����<�,�;�8$�~z��-�J�,{@=������ak�<��D�T�$�X&0���n<�L�@�ҼQB"=�K�<�yq=�$��nI���D�/=l;u���Z�;��<q�<��6�vh_�F2^<�K~�d�^�p��<���;r���(��p�;8�3�G���_
\���S<_?���U��!w���ݼ�A8�����j�s=�ر�}��˼��b�o���b<���;�ԅ;>�t����(��l�a�)��:*�G<y`��/^����<y��ƥ9�`�ټ��0�b���t��]@<��;!��5�+:/í�Z�=V�N�9h5=1T!=4x�~�|�I�b�� �$º`Ѩ<��a=��^�ı=Q��<Ţ	��H�<Sw=t��<��D�	A;=�h��R<�X=G��;�;���a]�$q���<����t��~�K�S��V:=���#�f��9=��u<Iԅ;���<� ��Y&=�⵻�"��ߙN<r�#<3;���=#�޼�EL=��Q�q��J=8�a=|��:E�r=AE�z ��'�<C�+�Q˘�r�<�Ƽ*=� =����u�",�c*㻪z=�j�|�������.Y�JW��r}(=�
;��#o����X��;|ݼ�Iλ�nN=#�X=%k@=��<)�:=F��u�95~ڻK��<���"a�<�|�<�1��s�<=>=��缌��<M�6��,,�����P�<q;<���l�E=�r=\�;�g��*W=�7<���:�j�<�W��7:����ߞ���J�7*%<R�d�ၢ<�"=}a=ʎ�<u1a<���3�4�rn=�$=)�J=�Mp������u`�U\Y�	��w��<U+9�m��<�CG=�f/��發	��<ђƼ��,��P��N�0�Pl��L�ߺx�H�f9�����a�;��*����<��!�6�<h2v���v�R9�B�<U<��PB.=k=6=d(}=�><�î�ԕ)=�L|�u�n<t��<�hҼ��H�=�������8��q�<5W�<�ph�!��<d��;sW���˼�~�<��<`�}�L�� A�<5�y=l������<��W��،<����$=�Rϼ}(�<h9=(f�<��K���8�e���d&���J�
�(p=~����仩{Y=8)=�˟�.��<�)��޻oЖ<J<�H����~�����<�F9;'@3�L�����g<�\�:�	�;_��Ej��������<�e=��ϻp����!�<�WN<���hE�<W�	�G���v=����I=�K�<|=��!=��Q�pm��Y���F��gc��& �V��P�̻�P���ļ�g�;fg=;�;<�GD�J��<���;�?��z�<��;�95<]^=c���!1S��%^���<��;��g�ʕ&�nko=��<���X��<;�Ҽf�9��-w��c���+��*t��N���"=�E@�q�!�J{�<��:d:�=��A�������<�-=3�-���R=Oi�����<�Z�<F<�����<QУ��bf�x1h��T�<�a?���Ի�6:�<�;'b?=	�D=!0D����;h�7=7�<��<�����%V=�#=�=yl�<��U=l�P<4��R肽b]��/���D=��=��/��^��+�`}�N�4=�S=� W����<�c8�_�=�󑼣gO�n*(=v<D�'<9�� �5=d�;:�=��?��y:`W�<ͨf:�l}�A6��]��;�y-���<�M=�?���uI;���#�;ݹ=��%�0�����=�c=E��<��=Ԥ#��.o;@;��H��U9f=r��<NR��t�p��<�59�b���� ��F�3�\���=�o�<�9=�\M=;2���]`<�w&=I�m���9���=����=d��8l޼$�;gbO=piS��6�<Y��y6<���=Kl=�n+�sOU:V�;(���-��<�r���!�_jX��4��ZJ���;��)=����N�O=y3= �=� �G���0u=�5f�8�G���������<�&���o/<��j�1*�<0={ǻT&=	�<G2�=�c=��H����<���`���Z�K�=�,�<�\�<�1t���5���+�؊6=�H��8�=��d���<��{;5<��"�����6��&�<�5T=3x#���Q=λ��7<����m�=-A}����<��l;�Ǧ_��G��<1.�<���<Ҩ;�Z��<��n=�=/�}</yȼ\S����xM<<�<���<�-m=(��<Z0N=3;G��~�괼3$;���8��;��9��S�*�K:��O��jj=�������<h�x<��|�xXS��2�� R�OS�#�y�^J=Nmm=��a=>e<�es�; =���<G�+=#Z�0&���p�����������;=���T����=\i��
=`Ⱦ���B=�@�<Q��<�Q/�D;�t�<@;�͜:<0��a3�*�<��Z�I3����<�a=��=�ns;* =7:��+K���<�=�uM��g_=�$1=\%��l�<�#���~�LP^=x��<Cg�<��<���K��<?�G=6&�<=�%=9ϼ~VN=If[���~�/ �v��Ž!���=���;�(Ѽ����:� ��5��W��Բq��=�w�5��~��f"d=�@ =w�K<!�;=�<�~���o<�MJ��H��B8��\N=�鋼e�����:)*=�	9=\<�:�����=ZK=�#�<?�<X�Y�[�<Ā�;ҫ�<�߼��9�*�9)�<S���z�=�y�<H�#��kA=�<[����X=�,��o ���'e=snF�F:��;���N=�Y�<��<H:=��:� ���<��O<|xf��=E��;Dz�EgD=��'="d��]=�,��(�͂�� 7=\\=��{=dy{=gO�<��=z2<J��;�7�<�u�<�Dl=A0�����=;�Ҽ�)��Y$��|<�""=ӟn<��=�U2=��|��ŧ����;EK<��; $�,W����J=�J�W�-߃�q���j�'=�5=!�x=�m�%�=�?��+=��޼����L������ܞD����Z=E�=�a=���cd��~N��?��K�％~�<A)ּ'�<����;�ݼHFǻ�A={K��1��<0Q\�~�K=�:�2�m�e�0=��)=	��e=-����=�`V=�Շ���=��N�:�J=���M<y➺�@#<�`#�8a�����9�J=@PL���=��W�s��rߗ;�ў�����;�<�.=��=i��<���<�OC�4����B=+k�����ڻoS����<������ż6Q��P�����<!�z��值��5�G����<�@=Вa����<�:�<�=c�U���L�9��M�=��=0���:���ܳ��ME�<4G��y*;�o=5Q�M�?�㋆=���J�<^�	�����@#�Y�$<��J=&b��Ar�����ic<^p=�C���;���<ѓ-<�����l=�1%�ݶ��pԻ{q	<P2b�	Pɻ�2L��=��#=H��)�Y;�ͼ٩<q�;�o=<k= Č���!���<pgx���;��5=�˼ YT��񼺭�f�]��<��S�0"<��a=$�$=�
�<�f�<���<6���;��G�6w��VP=�N%=�ʨ;�23=~��<A����i=XM�<�c<P��\>�<콛���D��:��A�<u�C=�SW=\��U����`M;ؑ�<A�<ӡ��^�H�(��G%;=C>u=؇=}�@���ݼ��:=��<^ [<�s3=}B=�gU��f��qC��(=߄6��)= P���a�/F�<ڰɼV�Q=���<�R�������G=�]+=��=y&��\���=7qq<�~e=UL.=d�r��=��<	��Cʻu�<6˼�z<�׻�{�g0<y"=�H=��Ż<�<T{=���.�i�q����;����\d=n�}���<P�;��=)����`�.;�#��MO�=v�:�큽��3< ��<ЫY<���</�n�IX�Cr=oEM=�o'=�Q=*�¾�� ߼���<�T�eݼ
�K=O�ݼB"%=)�<Rcƻ�gD<��K=���<��Ӽ��R=�Z ��V=O,�<��;��7�8��<�.[��'-<�&;k��<U�A<�y<�iI��Y=��+�~57=s=(�|�,��<�=�N=_�+���Q��u{�d	8;��H��<pA���r,H��+=3м}��<�z��;0=���;�}�<(��;է�"�ݼ���==��=���<4�ۻ;μ4�<9+����滨�^��ё��<=���zfv�auu��Փ��z��t;�<]U���<Kx���޻`?�G�мx�^;w<��L��<nY���4��&���@�7_,��f�<��F<]�R�#M:v�R��n=-ᄼ�=��F<_�T�G�/�)I=��M;��=�2=����o�=x�/���<kH�<��ϻP\��q����=�8��<�W-=�!Q��%Ӽ|���(<O��<C�q��S�:�Y�<=��<u^�<ː#���c;P���(F��V0=�A����z; ���9�<�=p�8�^(_=k��;�Y�;|�X���<J����$y���&=Y�8="x�<jc=2�P�.9�������^��75:Pf/�6��<�<=+[I�K�"��'�;���I
=����97�K�6=�G޼A^S=�e=�qZ�I}��]�Z�=�yz<�0���h<,7$=JV�3��:Z� <��������+�;{[�j�Q=;ve=f�D=�x��������<t��'^)=����I�+�=
��u�<5��<j8+���)�[�+<$n	=s�]=��P=m�(�Yu�<�>B<;�v<�j`�A[��!҂��kk�"�ڻwZ8��4Լ�.��H<�W$S=�v<1TC=��ɼ�I;�꫼h''��y�;��J�:X�=ש@=#�8=܍��/6�<��g�Ἴ+(;���n+	��@=�]����1<_���[ȃ<2����=�<U�=-7�Zq8��<F�S����s=�� =�8_���:���)=��n�9�}4���;�5K<��Z��ID���&��0���dk=�%H=�DZ�3(=�p����y��=.EQ����?�0���;���<�=Q���<���;R4p<���;��|���F�խ=�"E<@ꔽ~	`�?O��lO�<�K��x�y��,�;��<��Y<�y⼟<��<[�ռLh���$��jG=<��dI=?.=B�%=vX�<�Eo�}�I=f��z/0�Yt:��	����<0�=�8�<�'=�������03H��R���b��=#=a>ǻ\��;*=U�xj=�����;�}�;��<
}6=�h+=8�M=��=��q��K����o�j���,�Q�<�����ּd��s�߻����c>=��m����<b��<�6}<�F=D�=�<�90=�߼�==Y�ͼ��K<�)¼��I�z����V���=�j�N�6<���S׼��;=��=՝m�C;G�9��<5�;���ӛļ}�;C޿�f�H�Ǫ$��(��y��b�l�+�#�(�;����kP��=�-\= W�X��<�-P=�C>�l��{݂<�Z׼2�h�����\;4N��i"=��	�c6�<�q0�k����>Q����<+{:��g=�,�<ǘ(=k�2���=#U� ^;򧼨�d:D�T:A+��=d��r<�A����6=�6=�W����;�U =U��.�A`E=ca�L�@�3�q��7�<]֨<�UC=/�;�\8=��һ7fR=����R�>*ʼr׼��<��-�F��S��➻[��U�<$,�k��$�mM�qg߼^�>���2=�99�>�C<^#=!E޼�B=��/�3��������=!&��!Q�f���=}
,=�UX<2��|n<��E={��;bTQ�8�7=g��<�;���0R=�Lмc�A=y:X=�����-���5���b=��Ѽ�����Ь;�1�����;���<��C�L�=Mn=�Ȋ�
��<W��<4�K�dֶ<^�<��6��̼Fq�<�-Ѽ�˻׮⼖V&<��7=��=��M�y�:����e��<�E:=�R���j7=�qA;�߼@�=ER;�7�����#�4=Um�<�O;(g	��|.=�u=QV}=\�<��P<ߛ��<�
�<F�q�V�ѻ+ {<*FG=��Z��󘹣�����c<�F8��=�R�<���ͼ�E�u�?=�	D=�Vt�p�<!A�;�8;Gem;�
��*�<�:�ʕ*;�cU=9�%=3$=��K=���<�'<���<鿒<�tἮ�o<j�?=V@3�m��<q�F�&�M]=�7&�ilz=���6�H=k�6�+q����<��$�DeW���C=d��<#�^��ʅ�}l~�=H�3)}=��'��w=(*���-�����<Sj��9�<��
�μ�<�� :���y�k��b5���z<���:�����a=��)���ۼh�8��˻��7���<����G=�)X=�A�<?�D��~�<�@V��R|�f�=���;M$=sF'��>�$�R=�DW����<�L$=N����e�<	�<z�;�dT=uP.=���<ɼP��<�F=��<h=	�2�ż����<�Z<�;�<��=���<�H�<y��[TL=l=.<���:=$�"=&��<=f;����=��7="��8���?<ҩ���q��XB���Y��;�x:�!�<
�D���=�d����=x[�P�?�'"&= r�<(�:�<N{=��v;�*x=���<sFa<��?�v=��<�Z�<'�o=�Ӹ�4#;o���?�3���;�d=DH=����h=����ϼ]=n�<=q��<��<^�p�z��<?��1�T�8^�CR��
ؾ��"�<u��;�e�=��:=i�ټw���_=��t=�b=��S��<�R���u�<J�S��΀��Ѽ�<�1C�<��~��<ƈ� �C=+W=�ĥ:���%s��N�=��T�ǿE<n��<Wz�<O�#���=�KP��;=�'�(!�q�����==�ٺ1Y�����<��W����<���+��<��`��Ă��!s:|Y6=�&\=H�4��rj���>���=�H=#4,={������<��=a�:p
�~�=7a�e��<�����1=U�>�� ,��%1�](]=�W�<aU=k�=��F�z
�<�G�<�u3�6+0=�ؔ;��R=n9C<��~����=��!��P�<��;؋����$��@����>� B<L�<��=?�����<#��<Ȥ)�������<g�C=P��ۊ;<.,<\�B�o=�|(=�� ���<�97��G�<��ͼ 8R=������=/�=#g��y!<��X��������.���7�;���<O�<�!����<�?Y�������K�Q�����O�D<�2�n)��R��;f�����ȓ8�~gu=��<`�8=7K8�|��<�	p=�(7<ַ�� �Ƽ��=��R=��=��Ż��V=���aּ29�6Y(��s;BO�<�?�<�?=P��Dv\=�=B�=��<C=$:p����<Go���=�?<_R.�e���K��&K���T�fR�'�]1�<��Z�1����7��b�@G<�/���>=<�
����U���S{l���X=�)�V	Z��wj��;e=v�3=q>����n=uc=���<\?6=�
�</�2=y��<9�=���<�C��dI���5=��=+��jʠ<!���Ǿj<?����}<ȑ�<STX=-�@��p�<�:Z=����D�f�a�:J��`	o=�6�<�s�<��<O��<!��=�?�4���o��<+��<�d�>h��>��`��P��<�����Ҽ�T�<ĕ�n}�<;"=U��YU��e7�m��:��<���mv�<��� ��:64K=���<KV�1Q�;��C��G���?��o=G����,ļ��Z���:���%=�pV=��~�;�w<����4K=�6k=|2S=%<6=prq=(�;�W@��!��ɮ<o���`�;��r=�!)=gR��Q��g�`<�e�<��:Q@'=��S�0B<��2=l��@�=�
=�����<���<�K=�Huj�ix�=�&�W����\=��B�PA<�� <��c�P&�\j`=�!��ݿF�� �:|M��MF=꾛���m<���:�<)�P�rȣ;N��k*\��D����<EG-<VXl<��=�w;�G<}LP<�.=��Y��<~)o��O���&=�<�KB=�J=�1���T�C=� <W��'�E=�M[�I>=�=�Ľ�;��
=w9=4���[=,d ;���<t>=X���I�<7Y�<��j������B=L��<$�M<�N��Vz=�8��m�5=�V*��+@=x?;�M�<n'k��8+<~����R���3��\�-��"f=��=4��N��<�&]�t~V<e|׼�Z=G\"�J.H�+O�~��؂:=`�5�#"U:9�=eZ�.�v���h�fP=��U=\�u=�w�<Q�=���5���4�|�ϻ}׽�v)�F6o<*R)=6"�<a�A���x��7+���M� $-��!);|�2=FP<�_�<FH�U���P�<Օd;�U���=�<�j@��W=�#:.��<i  ����;�)@��Q=s*=�o�G�����t�� 6�<� 6=�ڻ��;�h�J�X���=K*[�w&=�d:<����\=sv"=�+=�B�b߁<g�=���㢼��=4���<����K;=q�=��=�E=�_�����<o�<�n�0�.=՞e���4��k��("=,)���v<����1�Nl�=&�<�`=�,Q�1����F=\D �m9����'=�젹Ta���<�g�;-^=_����=
*=�*=����np<<�!����*㾼{ ��_Q�C��;\&1=�3�<SQ+=��6�A)=��Z=�i�<f 9��͛:�<������<�m�ohE��C= o�>�S< �=�L���@?=e�3=���<] �A0�:bռ��<AR޼�������7�݇A=�K����g;��=��.E�5]=+u:=#�a<c�#=�m�;P�\���;$�7�ܳ��q�N�\�=S ��/XB=�<9ς=�ȗ<�@�;�]���5=�1�:<�.��Vk=�H�;�ٺY��;�T?��a�"T!=�+w=_.���m��Ti��9=����xH�wc��������<�e�֨g���=w- ���;�=����2��x�U�l�:�$�=SqC���\�`�=�$_�\v�p`�Q="Z ����<��]͞�A~�;.:�n�*P�w�м��=��5;�Dj=Crȼa<=�-�����:��2�;��;�2��b��4�;w}ü.g���Y�W=��$=*��<�2���=nݻ
�!��;C�)=��\�;�!=�p7���\=�_�<m�O=���<{T=�D=��+�� �<����l�<�% <0=CO)��:�;�j��tK=풇<}�;�"�	$�;םM:�$'=+���A�~=�����D���������' ����;���6����|�D��۬-�M�����=�U��Kq=��/9�U9��j���u���K=��<�Jn�<��H�S�/=&.���邼�\<�(3�M"�;B_���4�,a;��d�<��\<;�_�@T"=ѢK������Y=��&=� 5=�������<W#@�b�g�4nT���q=�b=��-=>�h����<b6V�6=��<)�q��e)=�0�<�RL<ݧ�<$�<n�L�� i�1�8^4-��v%:�en�ICK��,�=��O=�)l�?l�<��]�Na3<-{V�U��ʡ�;BM�y����`����0�M�������o��:=f�����<*<��.����<�R*=ͤ$=/D�<vH3<�^�</��<N��^�=�J���'fW�5�<JD����5��h~�q�<	�"�Vr��N�Z&���;���^��<��<�O���dP;P6-=�=�<�mQ=C�H�G��<k�U�� ���<=:��<ب�;�8�<��(=��<��L�tƺ<U�J�?�'�<��<Qq���0'=\��`!�<���}��<NP�a�	=�;(�\,�<�J����Z�'��:1lW=R@�H�<0�<�C+�c	��'=��3=zm��Q�<��&;�Ļ� �;b�Q��/0��.=��<D4��	R;��<����lt;1D�7:�<Hkp=.�м9�"=��G�w<�=��3=}'�<h�<<��;3�7=��e��4�=�4A�� �<��<�Q<7�Y;^
���=���o*=��<p�����3<0��&��<��<<k=�>�<�0S�s�j�SW<[n�<6c(<�<&!���p�<��?g@��:9=Yq,��&�;�Z��$)<^����<.[��*Ҽn�B�v%=K�A�c�й#����q!=ʍ��ǩ�܅=��<i�n={���|=��
=�\�<��|�����uPX��3�}�'=�d#=�
={��ydh=\<�uh��28�i��;�L�;�rA=m�4�� 8� ��q�(����A
�<��=7 �<q��Pw<��R=�o�x=iR=� �=��C=��A<Y��<?d�<�4F=�r/=�]<EF�Vh4�>�ݻ� �E�U�>�r=���KҼES6�O���}
�٩��~9��&֧<��:��GA��@b=&�w�N<E<���z��Wm2=��`=��$�k�V�xO��N1=���<Y�ڼ�D�<h <"ր=��	�K,��>i=�	�<FC���u���*?<
�,���)�p�@/���=�=[� 9W�޼�k:=x�)#=��<����(�<��3����R=��d��}���f0�<X�᷒��S¼7��<zt	��+E��r�<6[5=�}5��h_������XǼ��
<łR<2��k� =x�H<�_u<���y���1��!<��m�(,<0_L��E���<��#��=�)=��;��C���J���*<bZ��R��ǤZ���T��9�<�<��;�a�;Z��<c�¼G�U=(�5����<
�<�-����<�a�<��%=bv��ơ ���K��=�*=+�<�!�Q�U<q����$��<�&;b�+=�a�����G==�-(=�zd����;��ռ{#-��yG���<�_=��=�G�=�bq����<ڛ<mI���=@�s<U�~�q'=jY��j�/�{����<�?�r�;�d =#��<�����^��O����%�-��;�..����<�0�Y�<rRd=�(м��Ѽ�=�=�Ws;!ok<�E�q�<��Q����͝��êr�w�>��M＼M4��?�<l�Q�꼰<^�Ǽ�/=�)���r㻧Y+<Z˸�����x�W�O=c�Z�g���:����׼/x=ȼ�6<\=��=��	�m�ռ���;�#=�x缏�=GT=Y	�4��<�M�<2h���<"�<k�8=Y3=�D�<��%�!=FҼ�6	=+�=u��<.V��+�<�X���7="r9;��=��I����;,�'=��ټ��%<����s=�5=i�м�Y.=�&�<�.���<A�T=���=3��z�<�>�<�!:��*���>���:Ҽ�B����⼹/�<�WF�+�%��jV��b<�;��
>(��a�Q=0�L��=u�=��	���I;�2��9�����8۟�FBF<hU�<��=a� ���Q=Ą5=I�W=
M�<�X=�=ƿk�?D�<���;s�*<�<��ؼj��<\,������'�l��+Ӽ&��;��=���_c�<�=i�U?�<�>;�6=u3�<R#��-���s<\�4;&��<��0=1!�;W��P�9ʔL=�]z<#��-s[=��=��
刽�2ڼ���sE�;�6��Z~���B)=���<�U@:;5=x�'=/3(��⏽�<s���
���"=��q�t2:=Ai=G�C=��<��Ǽ^��<�6H�hi=o����ݢ��P�1��<�,�<b@��G�6s`��.�'p����<���S=�\5��ܴ<�<�a���|P<M�O�Q�X��� ��Ƽi�F=B�,��Z=mt�;X�5=��μ��<��=q2=��<T3�k<��7:��d=5�<�W�;�N�V�
=S�<R5<E�<ugR�_�o*N=i�0��<aN*��՗<���<S���F�;��%=���<u=�G�<
�0=?�c�夙���K�3�X�*�gD���׋���S<�#=0=Qj=�*=�t���ϼ��o��ϼs�9=�B=\P�4k(=}�<qv=�� �+O�<��=t|-;��=~�ۼ-�=�=ܤX=
�P��;��:t�<�N+�	E/����О����˼�2G=��H�@kz=~�=={J�<���{E�� ߼
+������`#<ݞ��#
=3�N�W�L=�gK�{>����<�<�kr�g�S<��H=q����@=rb?���<��=�����%�˿�<\�@=N��<�UG:�'=�*&=�K=�l#=S�|��*��z=\�<Y�{��l�%���:�tܻ)�&�=���R�<gbi���<L�^�vJ=xLZ=�Ҽ�"��o�;�	�;e=�i���;�|	=�_\=ps�<��,=r�<�J1�ŕ�<PwN�*��<��l=|GT=��a=���;�'�<�����=�I�<p�-=��<ݱ�<��<=�%o<?6�:V��<��4��� ��<l��<��|eW=�/�<b��<�m��ٍ<�6)�Q�4=[����3B�h��<�M强oC<�G=UҼU*F=�J5=ŕ�<�6�������t����Z>=ҙ��s0=�M�<.6�1}8�8�<=�\h������=�嬼�����i�<<�L���ּ���;�mo�;.��{�^_<.m�<���<k�9�i���]�<�(O<��Ҽ*�V<dT�;Rm*=�&�\֥����y���,/=�)�=w��W�f��c�<���l���=��!���z{=��
=�c=��!�V/���=�<&$=�V���A=��k��\�=�S!=�W�<��;�Ec��@C�
)���N�<։<�;N�Ө��!�+R?=w)D= �*�a:��b��.f�k�?<�#���u�<-��ͫ<��Ѻ�$�<-��x��<�PX<�.G��t�i�?�.]��{,�=�u=�)��$9<��"�;�><�汼J$�<���<8�<��;��b���=���=K��,�P�Y� =|�*"�<	=k�(޲���<���<�,��Y�:�+d=Q�5����<4Aü�=��?�:$C<�|�=�`�4iY���\�����μm��< �ͼŨ1�5<U����-�B=�� �l�0�-�6�����;HlԼT�<q4�i��a����<O�<�D]��ݒ������MZ<��T�]���[@=�R<ET�<�F@�k��ދG�;��"=T,��d��;[�w=�Q껰ݼ�q4��[���Q��)��T�<��e=C��$l<�Q�Y��!/=�^��^�?z�=޻C�2��<yǺL�<����:�;"������ݴ/=��=܁X=/ᙽ�]��� ^��V^��-T�S4g���9]�ڼ�`=Ȉ�,�q=G�K=�2�<�w=���gb= �M�?
=��2=�D��eg��e�?*N=�����=XUM=�0�<t���ٱ/=\�<��g)�R�'!/=zI�����<5�=���%�A<7�D<K`q�֛��h��;�.�\&��K�6=w�C=d��=`�k���@<KE�<�F$��9L��D�;?. =>�9��qV=��v�|�J=���<��#��{>;���;��<p�_�>
���7�F<
8=�zQ=Ƚ�;�f�2!=e��<��A;�`,<�S_<�NE�޼
c.=�}�<� �;WM���ȼ�6#��ā��^R< 'K=G�|<���<��[��K�<AF�<@rS�_D8����9�B6���p�Thq=�"=�X�Q�3=Pc�<1�l����<qg��Q5���`=.T=T,U����<?-}=��!<0R�j2Ǽt��<�M0;ڼi4H��73=A��Q6m�e���M:7�t�����d��9 �"����䙴�8��<��伸ࣻ�V�R�˼�hh<�mG�h�{</�	�H5������5=	O��Y=$R�td^<htV=T�\���n<�?=2�S�q�<-'��(=��v<KHw<�{9=`=�y<�L=���<��;ve=)��<;+5�''=.��~�}=��K=AWy=A6	;�G.=�'���f=B�]���e<�+:<��,=T�2�s��<o��`����{�RO=��ͼ$��W@Z=w�7,�I�)f�DjҼ�&�<�$�<�N=m!R���t<d���Ek�-Ķ<���<H����,�T��I�<�ּm�=X{��%ȼ�5��9.<{���F�'=� ��]&�h.�;[6�� =�6�<"�;p�U;��5�owM;����ǆ<���j����+�<5�߼?l�R&<~���^=hC�<u�<$���v����ݼ}���^���K=b%��{��B�$";��N�;��I���<0|�<�ߘ�^��ql<� G=���=��1=jB���}��&a<Sz@=��c�"�8�<{�y��i=�m��=8E<Z-=�O=�%�<iLs��0����������t
=��1���<��'��<J=F�;��<��<��ú�<��Ӻ�K=oY=���-���S=��=u�g=(�)<��1����<�\X�D<�u<P�&=�Ԇ���<*��;�2'=<�N<�C�<��y����ӊ"�!���p�2�,=1#���9y �O�@=�볼��s�=�9Fլ���C=
Q���$�F�d��g���=�٫<%'X����<� ����<޿S���=Fqu;~��`�<?��<�t���i��%=��1=4Ά=])#=_6:�	�@������ױ�Ϫ*�J= ܨ<��@=Q%S<~�;���bC�tk =E]�9��S������� �o<b=���oT�ö<�Iy��=2��<��5=��f��H���o<p����R���� =y�8��mA� =��_��K��>=�	0�=� =U�¼~�9:��<v�<�6E�!�+<��� '�T�Ƽf�=��=,G2<'z��(=���`=5ꈽ�;�<�u|��bټ`��=�dQ=�#k���<.<��26��Y�}=S�;M������a��2�<T1�<$�;
V�<��D=�+�;d|���G<�{={�i���,�����i���l�;�9��"#=ݚV=��9;7���7W �c�����5�E�<b���|���s��n�̼Θ(���<3�ɻD���0+�2�1�F�~���|>=��-�o�л)�!~=�4�<�yʼ�:E�M��FC=�<��=X��<�1a=��}���L�A=�ؗ<8��<\=�(�<�I�;��<2�=���;�>�<�������=�W0=^3(;�D�<v�>=iU�<h�0=�?=��K�C$,;���b��;(�=��,��\c�lT=��6=���<%����h;����<7��fPS=)<�EQ=MJm=�n7�8��� ��$�B=��l=��d]�<��/=�%M��o'�����$Z��F-�|���s�.���j=u��K[=��s<��ͺ��ѻ��;r��g1�=�@=%�9���=�=Y���2BU=��<�'(I=�?5=w��_�]�X�<J��<�\)�U�����<^B�;��3y/<�$E�[��W�e=pSp=��\=O��X��x�U�����E+�<tV=E����<�;s�l�5=�Fû��hY��S=���<¦�<9o;=�U�~%��',�cC4�k�C=6�g=,Ǽ�w�9M��=��u�p	�<h�X��.�<�Q�,c�k�ʼ��U���M�@-=�U�ruz=�]�^tI=��F�۵V�_���&= g=�>=�D?<.f\<@���ͼ&Gb<ڵ��=?w�<�ќ�&G��*=,��<�
;;��e��#=�=���<�0\=��`��x!�n�h���A=� �<zP�<�"�*�=?�W=$�W��ϼd�#=�u(=��ӻѼ�* �X�=[���"V��0�<�6�V��%�a9=nS<��<I '�B���������(�ǛL=Y���F��<%c�Z�N=QJV=��亂���2<�e��>̼���<��=�.'���ܼ�.=��;��=�u����M<X�<��<<2��<(O=�:����8=W��ľ=+]��Z��扼���q�O�d�D��6=�D=�v��*b�EK=��;���k��<�����;Q�=�
��OR��:G=<�@<����<W�9=]�;�eչg蒼r?=���7=-D�<�Nz;���<r�<p�E��i���iB�#P=�J<Y���A�=�l2?=�Zּ�"��81�;��&�<L���y��M=Q�����R�`]�=ӈ=��'��w�\��<�"�'0����-��*I<�x9��l4=!%<I�c�����̼7�N�O�==D� =���Ak��0l�{�<)8	:��=zK'�Ѱv�/�^����<0�������Y����4��'��=xJ=��������~��H�;.�K<S�<9�I�쑆�_n�z�2=�-E�Pi�9R =�np�[Z =4?�
S�<k���Ќ�� k�����k����üK�Ǽ���q�!�I�*=C~�=�aR��?+=p��/�=;�=�G�]=W+K=� ��b��<�yA=�'�:/�<��8<P]==��;�?�)��,I=SP�
�;��a\�y?ۼ����Ӭf=�ʘ�?V��E ټ^�=0��
�=WU<6�=~��; ��<����eHp<�}���Y�7���w/��*=�=���<R��<��<it�<j�g�� t=�u�(�H=d�,���@=;��<߮Y�ʫ�����<�){������<�>���H<���:M�=���<km1���V=.���A!�<�@< `��Z0�+ Q�	��<�Y⼜�Ի^4@��ML=��E����;�E�l5=�}�|J��&�x��T�}>m�68f=۶	=���<v5h�9�<PA=�V>�M-��������'\"=5��<�M=�A���:�p<|�ؼ�=�R�<vBԼNA�;�f�<��;cݤ�K���\�̡���,�		O�*�μ�a���<uv7�	H�=[(��X����q=�i�=�X�;8v���;��;46=�
(=�	�<�����<&�=��<���[!�<��^=/�A��PR��P=# �R+�<k�o��d����<��g0=�U0=p����=a�,=ڍ0�d맹v`+<�0=O�Z�߆[=]Xw���|��F^= �̼���<}%ļt�s�׼�?6�.x�<U�q��Dv�����M�;.Ci;҉j=�R<Z��і�h�n��⋼�xo;��<�Js�J6T=)<����b=��j�A�=}% �H��<ņ�;E�{�I��<���%�_���!�g�ּ�����0=����^��D�+=���;�-J�{^ <O����r��ᨼ/xD=�i=��d��Pl=?�5=-�=k,ļ��'�\;f<�o�<��ܻ�=Dvo��x���K�?r=/K
�g>��u�<-¼NK��Q�<h=�~ ���E�8��<�+m��>��	�v<tK�<�� �XGN:S4F�O��;H��;2#�<�Sw���3=�q�;���( 0=o[ؼOז<�+=�lp=.�ɼ!����D<�Q����<�j��a����9���<�2�<	�n���ƻ�z5�6�=�,8=`���硞��z���==V��<�½��zX�#<�*�
�6=f��&&k<��Լd�4=�5=�:k$�;N:����<"U�����<z�f=y>��D�o�kH��$<��5�;l%=�
��F��K�[ <�c�589��(=xD=�q-=8´<�9�xZ�<�9���$� �����<_i	���:���V�M������P�f<YL=4���4�����<�)��ɛ�=���<JX��eL���6{�<��<��j<�[=̌i�#�=>f�E�"<C��<v�c��E=$��=����_n<��[��"<�" �@���;f�;�~(<S��ER��ZP<�F=��r=r��:�!=C�7=f� ��)A�r�J�sGX=��=���?,=F�]<�伦I7���!�䛞<=<�\y<��;����Ky�=T�=L�Z=6 E<k�ż�,�:� �ƌM�}	A=D�b=�jt=��s;`ټ��<���<$��<\�-$��$R=���TF�<��"<4��<���<��H=hՙ�B,C�9@L=�;����N�N�]�J�<2�s�ú�|&��<@ξ�n��7A��t�<�="֙<��Ⱥ�Һ\,�9*/�;u�2�颢<��ӻIg�<g�h<�:=R=�ǻ{Ļ�}�%�K6�fg:��n}=*Y7�(x�<�v,�v�	�e����<s�'<˫G���U����O:`<�=C��]����;}��#|v=�=	��e��o�==GH�(�v<(�<��ѻ�8-�� B<�Y��ܯ���>�@<-�<�MЕ��\���.;X:)=��r<qt�<5�X�;��R�<-�<����ȼ�7;��5���?����.��<-=~�s��|b=S�6=�����N0<���L���;=z>��>���V�;@_=�<==�y�)z��8��U���}�����;;t3=�Q�<d������u���-=�2�<�b��Q�<���;`��˕�<f���q\=���B߼!�$��5=�� ���7�T@�<НѼ��9=3�H�>;;�Ӌ��Y�<������];=��<~Vw=��o�Zӹ<(S=�)=aZ��k����%=z\�<�
��G�2�Ii�<�fۼ��2�h��<�==H���&J<$��aO��% U����<�_G�d������� {=�:=��9�!�<�Hλ��D=� �;�H;��N=yQp���I=v;F��p���H=��m�͙e�H��</$�<�==�yU���/=�F���<6(<��Y"=U�R=q�;=��
�n�9��8���<��<���;iJ=�A�����t�C<��l=Kg=�68��M�_9�<�
�Z���n�=,^�<���O����!�<�C뼣��6��������j=�W<�"༑�<��=��=��X=�u���L�@�<�(���hC�Y	���Y�H�7��o��h9�m�< Zo���=��ػ�()=*���'��=�<�3��Y��:�BC���ļM���b�$=r�=3�6��~K��Ą��0��V=R�E<��]���B=��;�1�\	=�g�+D1�k�(=�Jü�<M5����g=��>�� 3�@db��*ܼ`�E���N���F=�»;�;�:�����^<��7�8d�v�J�H�&=���<|��a��<{�^��2.=�,�<M�Y��eP�G>��$�<Ţ:x�;�j���`�<��C��JF��#�)�l�Y �&J%=��>=����)
�_��=�<E*=B$��>¼0��;�M⻻�m<�\�s+�<(VQ�Ѭ�<��=����<���<cּ�������p�b�;=XkF����׶H=?�A=h1�<3��<����=c�:&��E�/�7��<��x=�4R�N��<��<�W�=ߘ���5=��*�����A;�=b`��]8���#;'�ۼ�o�<�$����ۼ�v���<�����(==6}%��)[=(9�D<=�<[��1��n���պԼ�1�3S�;����%<�M=͓D=��<�w�<>H�<��<�}�<� ��]u�Ŕ����<�(.=e%#=v_;Э~=�Ŕ���=�|�`����/=<$T=erd��,=vu��:�i�������<�E��`�=�<$=q�[�ǐ5=S��="ï���=�>�]�"��������[��d��<MU�;�	F�~X��e�U�|�<&��9a"�F~\<��6=��`���*<�|=�@�<G�C=<�m����<��'<�μ���;�����8�j==mߔ=ͻ <aa�O��H40=��<?��=7~g<[Z=>9=��E=FL�<)�i�BUA=X��<�C7��_= �S=!�Y�Hh^�w�!=�����U��<?���.p��༘=�<��N�5��<������=�Sؼ$,k����<ߥ<�,�;��R��J;�#��c�!��Gܼ�C�:��P��\=�g��o=I9=f�=)60;���<3�ݺW�<����w�c�-�"����<<����(�;��5=A�m��hF��U=P;�����
Ѽ��T��0��ѼfC�<%�;���׹�;)� ����xy=߾7�
t�5�M=*ؿ�	�p<�M�k��<x���$��)�<=�Ȯ:��E�%=4��1p�E��<�F�$�м�<]N�����-=SA� ��<@M);��P=܅ܼ��K�r�	�G=A��[��cּ�y����<�`��<4�z�K�9����<hɉ�5$�{�u<�XH�=��<�n[<R��?��܊=m�=�E�=3�==��<$�c���\<��=�[�;���;��8=T=҂���(�W�r<{|�;��H=t�<���=��v�\)=��ռt���x'n�����m=x�<�q	=�����I�`,=���<��R=�y���-�h8��]J�0/�;%����0=Q�F=N��.B�~ل���U�1O������뽼D'	�t[�Y�=_G5�Q�`;��)�Z:�䊻(�=�����<���>�e�d��[/��D�=�4�<EG�<sRX��:J�*���{��K������ �=�#��c�<1���M<�lZ������<��G��/��;=N�N$#��O,��JB���<�\�;��<5��;]õ�Q�A=KKI�S¾��J<�r;<�m�;x��<� =����(��<��
=��$<�f:�׺<ҕ=���<�)D�2�r��6���Y��Z꼆��;�9�<��)���b��^�]����-#f��#�;����䬼r��:��{�9��+~C=~V9���O����<�ᐼ�W�=3P"=``�=�̒<�+=#3l�U/O��r&=*O;>�g֒< 5󼪺ͻ�u�<�b;28r=�:=�C=�b<i������l�]�U�ϸ��F�¬�<n���}�<2O=������<�J�ǐӼ��H<)�7=��<eN�4|=��\����|=�]E�_ ���<���<"�/���v��=��B<l6���Q��Fe����:�K��_/=zZ#�<��<
�<٭ûS_���[!=N�Ϻ�%S�<Y�9�? ==#�:��� \�,AϼŤ�<��}����"�O</��<|�<�Ԙ��X����&�|�m=|�e:o�Z=�Wf�5�=�.:<Ţ������U=/�=�.������d�<��k�Z�y<�@	���<h�5=&���GH�Y�6=���<:�=����g��� ~��R(�ʞ=�k<͑X��=*=Oy;?��;p��<�<^@A��/=t?��&���u5���a��ش���<S18<�5�%=~�'����<ê3=['ۻіD=�f޻]�E�èM=d�H=G�^���}=�Pz=7	\�%x�<)lR�� �L$?������L1=�Ѽ���<,R�<�:����h<�H��[�8;=�h�<J"=�R�<u0'�;�ʼ��U=��=�F�Q�B���=UP�K�<��<0�`��D=���<�O�;�F=1s?��ޣ;ϫ����Y=��A=[lo�����O���I=>
=�W=����<N�	<�}D���3=/��q���M�<�<���^ @�2%;-\=��<xg�x!ل<?-�w�[=w�=�E���5��6=F�,=��z={�/�@�<�9�<�9=���*��}���<C����N���~���=0{;�q���ܑ��ĻaBl=57���<y�;��L��=s�(���n�ռ��:�):�)��
c�<,�ϻ�:���*<8�=��=��t=/8,<�φ<ԈQ�ј��eL�M&��堼�sG=Q8���eҺ�Gּ8��y�O��^�<)/�;�����m��y��<��<!"W<А�	=k��;܆L=���ҷ;L�h��C@=�'�<}TW=�in�Ke������=%�<�ܥ< �T�&��<P�=��=K/\=-��<�J�
�!���=��f����<�W�N��<�'=}:=R�T�-)���a>����<˩>�/y�<4�K=���>]@<��<^9ӻ�+Ǽ�iļײ����)�?�;V95��).=d�ȧ�;<�^�LC=�H6��~�:,引v5=L�:��9=�6G�r{<!\3���K����qI���ͼ0?4��^�<��=�2��<�g깅�B�G�u�L�ݼr#]�3��<�b�</V�<
$\��e=^}w��)���٫�o���j�`=TBh<��6���ϼ�B��+�<�)y�y�d��ܹ��X�X�:��pM=Ł=a�Ҽ�<��4��<%=�:�g�ﻇ��<�R4���k<t�><$��;��N��K�<�BA�G8=p���[@�:>� ���̻�o�<�
�=�%�v�I=%'�f�<���;v�%=ߩ#=+�A==�5P��yM<��b�זw=��c�^$�;��H���;;�x�<��0=397����<���<xCD���r���<�����=d��<�����<Vs==�6ɼ"�&=�)=�=�=4X.=*0�;�<���=q ?��lB��:=Z�8�h;G��i~��_��Aۼ���_��C	�<�ڭ<�ԅ�`�]��?/�@o��LRἯ�]��qϼۡX=2h<��5�C<����oC=�|�<x�=�:#���%=�xw���.<@���3 ��j^��^����'=/=ڟ2=�DJ���=��&=�c/=�K<=��r��3=�]V=]9<1��<хE<�F�هP��bL=+Yj<^�0��=r�)���=U�=�p~;�Ļ�})=@P=�4�/+�x����=����^R=Q�=�T���V|���.��-�<�*ɻ��@��l=�!��z=�r=K��������V��c9=^�!�tG\�b/l=�K=,wR�H�ļ�<�Z��_d����;=ޥ�w�=d�;�F�;6\@��^=�<������ɛ��ݻ>��L6�<����:�V=a`�;�'=�_ػ:GлoE���=,Z=_Fʻ�1�<��^�(��<j�k<�j=a9�<�	�<>�=�Ĩ;4Y���[<su�<��6��5*=h�$��=�1x��"[=�b��-aY=uAἘe�<�/����<��;���<՛<nt3���C=f��>�<̝@���t�`/��k�<�@<�7�<��8�>�,;%h���U�K�E�n7�<�6c=�1<F�4<g�!���5�m; ;ʫ*={�]�ۼp��2F� �_�B=c���'�����H����;�ڠ��\=�S�U�� F�nQ=Rm��t����Ti�΍���?�<�|��:���Q��cN=��#=��μ���<��߼+<�X!=*=|�&=v �=& *=Dt�<����v=ig	=E�.=g�r=�'P=�\<��ɼ*�K<�4<)D�����K=�獻��=~p�,��WV=�lJ=e-���2
^=�3<l=�9��R��3���HP�tV<<��"~��,����<;����ߘ�<L=[k�=���<O+���D=:?�S�b=T=�(�<��;'��!Ui=5�8�B�b�3�ؼ]W<5����D=o=�Xg�^A�9B��FF����<x�o�UP(�
;z-C�h��<Ŵ=�/�[=������Kf�s��B��@����L��s�ռ){�\�;�y@�mf=;l��Y:��UM��Oܼ )�� �<��<�N�;��<�]=Nh���t�_۔�ݮW��9F�*m&��O��+*=N�C�q��<e�\=�^�=H�.���!=��x���N�F=�!�7u{��l���C�x�p�z�V�<�)<о����;=�w�<�Ao;�h��*:��n��Ү�;�U�;���E��<k1�k�!���j�el¼��h=*�ry���=�p�s�7=��^=��<E�d��5C<`I��W�<a'=S=�i�K���Ԭ>��������<���=I1Ǽ�l��[��������<	8[�pfֻM�1=4�� L�<�[��N�U����>&�(�h=��<�ɠ=�Cb��I�D�+������+X=��5<���;�F\��Bļ3r�L�`=Ӌ=�?��;�<���<Xû;nn�������;P��<-�߼��H�=����;�,�=���\CS������Q=�]5;��R<mM5=M�*�%R�;Ш���;�_KR;3��<��|�4sl=�U=:���W=
�O<�ϥ<�g=���l�M=܋���&�I"�;#�ּV���q'G�0�@���%�d�+�p�-<�=���0k��Q=��%�&�NkM<��,��=s<��^�;�C�<�J<��s=��q��<�����\<��l�+�y�n�<o1��q�=o�<p�U=��v<>{4��眼�7e=�|�<���}|�<D.x:�ȼ��B����%=� ��Z�'�8�:{<���<;����>=$�=������'�<P��<�l"�kA�<��^�w��g'#=��7y���}=@qq�W�=N�=P����.<O��<�C\��1X=7��<Wq#���=��<=�܁;o�f=?(��H�:k�%��=$��<8d�J*M�I"=W8(��=�-�<�aM�8�j��<�6H��

=Q�����<��?�N����;����:-=���&��鮍;�p�<��ļ�D���f!=U�U=�,S=�g<������<5��/q$�ltA������8=Щ��^��<,d��8�B�V�I<�y���<#�D�ۮ�<^1c=)�8:f8ܼ1��r�<�s=��d�����@�8��=�N[=��bռ֪6�xʼ�m#=?�����<��-<-�`=��������5�==����<Y=�D����=C��(�
��2�3�F��+*<�i�-�=vq���_�)�R�������K�5��{�<G�z���(c(=�o=��<M7�<j��;w<ڃ=�়�=�si=䣼^C<��)��Z��j]='g^����
l6����J=d�==]\
���K������F=�a3��oO;0c�< �����<�t<"��<�<��	��	ݼ��.�k�=��O=�qI=��N=�,O�%D=v��;�k���<��0=Vy<���)ߌ=8H����;c�S=��=�j켻4=4��<F(�<,o�M�N�l+=f2�G<=<@�=�6,=�^��1��p����;��
ּS�1��8<6����s<^�	�"�<-�;"��\,E=c��|�6=��;�ݼo�Z=S'z��=x=q=X����P�8��<�;��#�u�P=���;��;��}�4ѻVԨ<f�"<�Ỵj+�Np1=�g1=SƼ}���73�<H^�<_��il�IyM=ˊ<�m0�<_Ϸ�ޥ�<'[��0˻�yd<*��O/>��뎻���<��<7"�;���Y=A7���Ҽfi@=�}�<Vg=�����j���=�I=< �<���{E=��W=�e=R�F��g=I�F=rT<�C��"�<q^=g��<��޼��w<E�<:�߻w�E=�.C�>W�HE���rM��_�<�DW=��A=;�=����L=�G�=(�<�<��=c<���*��Z�8�W�3;#<��&=p#��b�P=��k;K;=��H(��^=����dZ=B��b�=u��:\��<�[=UAK=��X�s���l�5=��<r�ܻ
#s=��^���S��;�:�[@�L���F;�K�H=�����r=MwW��A�Q�]<� :=�8� 4S=3�l=��*=S�`��)=�J�������=&=9�.�$�=�Z0=FKo=
�v�=#	;<��<��p=>��;�ă<�o�;�=�B����#��<�[Ҽ0S�<ip=�Ϳ�������ʼYG��ؼ�S�|��;��=�ˁ��t���;=t�/���=*_$��mݼ��0��R=���<���~:.=�܄�]�=
(�<m"�<���<��+�#�ڻE�b=�}y<L� �r�K����S� w=�M6�	A��H�*FJ=d�D����:Ei�<]�<p����1�;�v"=�9=_V���$,���7��޼�漧=�?4=$����	�<<�<j`=9�9��\��u=s�T=Y���ƺɨ[�{�ɼS?C<�������G����2A輓�/=������<�}j����<e�h=Ow;�@����2:���V���-:��i�:H��� B��;<Hh�<h=��;wd<�~4�(Z�~9w<��K���/̞;�̳�K��\�C=�KW;�Z���=�g�<��{=�,<"������F����=B�<{t�C�ڼKm"��db��7��k1=+q�<s��gG�<a6��̜2�r�;�v_==E�<4��{�μ�Z0�������P�v���e#¼'��Y�W��K<is=������<R�8�)9A�"NP=�cż��9�լ��м�=Um
�Oi�k�<1l�;1�=���)=!g�!�z���=ɍ=�bM=�u���N=0�ڼr(<=`I�:�PD[;�lP<��G=�f�<âF=�=*=�f=�=.���<4>�<�=�sK�`�=1��s2���'>=��0�*=�xN��帼�d5=-���=r��<S�=]k��G=]s<�9=L��<�qU�(��:�V=�� ���������a=y�0���,=�{=�6��ݢ}=W+�b_=�`:��3=R�>�8�o=��<ܾ)�+K��G�U=Ԥ<�3=�'�<m����<C^=8�����/�L=�?�<7(f��== �<<�����4<w%'���0=�s�<��b<kQ'�k=��^=G7��:����	�>0�<	��:G<%=�+@=�a�<2g����5=Rxm��J!�~�<K�d<�D��x6C��JȻyI��TR;?�_�ϊ<RGP<2�,=���<Fpa=)Ǽ_�ڼnN?��V�c'/���l��=
#�^�=���<t��<?cR=h��;[��<:���[���ϭ�&����P��`�?��,λ��[�Y�&�F=L$�����~:�!�VJR=���<7�=��K�}�h�=&��;Ax��q�ʼF�=�D�<=='��<mY����O�=ňe;�0�<�=[C#=H�ż�HA�FŜ<��D�wiZ=���o;�R����<?�^<G�ļ=L7=)��;σ=�����k��1�<,Nk;��(=F���`t�<��j�L��;t�@=!=��!��2=�8<�N�<�� <�uC��ȹ�UW= � <��0=�&<�d1=��a����<+Z޼�GU=��=�;���İ�+2���o,=SB����=��»\A�<�y[��~=FL=po�<�j-��	��M�s}G<�����r߼B�1=k��%� �L>:=;�<�ԁS=���GZ=�+!�EhB�L1�<�ﴻ��r=l�<'�L�ؖ�6�<{�s����<�0�u�<�^�o)��da=�(�V=+T�gFp<aW=qU��X����_�\�v�A�%[�˧`<L�<%�=B�=�;�>����AU<s�<e��<@p`=���<�D�QH<��<�Fռ�,��B<ܾ�����<:N=,��G�.�,��7=�1i=�k�<��K=j5�<fu0<�^���� ���z=!'7=s����D�<y˸��sH< U�6D�Ƞ<_r��*=&�s��9U�,���`�S�[g�<I�e�_�?���8��.�>j<H�9=-��<�-E=��<��<=�N=���<�z>=6�c����<�^;Ԭ�<��"=|i��pʟ�Ik<���<��J�m{@��X#���A=��T<���U��h�H����Ҿ��_��<�։;��-����<�/=K��<ǿW�V!a<莄�j8�2�	���<�R�d���7�A=l ��V�7��"y<�=�j�<V\�<�mp�X+X=�4=<��G�Q=sv�:Ø�<�)�=�*�B�'�k;��=1^��^��AF=�뻵�<��;��<r� =��E���n3����Xh���<k��<�SY=�f��c=P�$�S8�<`���!8=f��v�=)�=~j<P��l�U=C�G�D�����<��C=T�<H�|}��'��9:���A�w��<.��C�M����<�1�<��Q��H=@lӼ���b�7�=��<E|=T�3���;UR=�?���W�"gc�Z��<D~)=�M�{e=7I�y�?=V�<�⚼��=��]<,�9��z7=���<�S�<Ӽ�<ڿ@��7$��#=����
"�b�;�i=<��>�<?F=�Y�<"m�Be���=�c9=:* ��2F<���<�2^����<���:��O=�>��gU�<S5��/�#�� <�TJ=�:};��������E0��\=�+v=�}�'m�;ʋ��&��3E=m���査9�O3�(�e�A|�<�,=l��<p�鼪68���l�/=���<T3%���=z����M�CF�<�)k�=�S���J;9	I=�� =@7�QL<T�3�A=���_��:#��o>=a!���;�J\=�+)�R�'=�Z�x�ź���<&�'=�@=��@�>��<��<��0=9λ��߻�c;���<�9<����*�2��~=>kT;l����㼆�=2��<K;S=��;=��D=�	=K3�<X���*�x�m�<��*���=��=��3<3Z�<��%��ϧ<<=�²=�'}:PR�/�x=%�R��Sk=oN���ֹ<x|N�xT^=d�=iG�<��4=�f=���=�<��༕� <�*� ����0�T�����K�܃d��������P=b��Rpy<&핼
�����
<���y�λֿ��9R=OI�,�R��]�<Ԣ�<.�޻J6��
�=Y�<�ϼF�D=&ͼ�\�rH�t�H��T!��qM==؋<Ԣ~<�H97:���=��X=�-�qZ����;�5��+����E%s��:�<�K�<g	�t����:<�jl�
M8=i8���.�D���?��<�Ū<����?�<��[<�o<wz�M���e�h��
1��D����<��=E�໸���dP.=�B<$=��`=y��<��T9����ao��OR"��p�#�lbX�{L�<&3���ہ���g=2�b<ظ�:�2�<ϧ����<諥<ꗸ;�t&�怽N�d=£e���P:֋�B��aD?���һ��[=E�&����nYi���
=d�~�@7=���K@&���B=��7�yU<Q==�o��Bx<D96��P�;H���c�<�@<僊<o�C�L��)j������Ζ=<�M8M �:G�<\�\������s<j���P=.E�����R��D)��w�z��;�ً;�v���k���P*�h�B��Z.=�Q=4��;M(c;jV���Ŏ<62�=���<�S~��V+=Y��<eX]=�8O�x��j9=R����<��<{jN;��=��P��wҼ�)������]=,�B=Z:�<�����?���/=��=�:��<W�r���]=y=Ka�< (f=Ov?��� ��v]=V�+��|��"�ܼD�.����{�E=�$��83�  2<�� ��<��-=��b<a�;�5��K�=���<w;!=� =k9�<^�:�L�=��o<E3=~=�����F=��'=_Ҷ8��,�Q*'<�Ȓ<�c#��p�<ϟ�<�	=s�=L�ۼ"�ڼE�Y�WT=�񞼌k��v�V=M\Z��<�0Va=u\=�$�7Z�<w	�F��<d�<���<�2�������rxo<v\K=[!�C<�''=�_q=K������<�G9<>��<�}\��V*�e�뼭�;�r�
��T�;�J=EϬ��𡼶_�<���<��>�u��9��#=B( ���<rl¼ܖ�<�}g��<L:�<ٌ<i
(� ���4ɼ+�;=h�k�V��:�=@�[��i�=� {�"�R���Yt���-:�Hֳ<D�<�"|=��̼�e;T����`�=�<��J=�1޼܄�<yv��y�/���(� �H�\}Z=�rt:EF��ْ�L�<�y9���^<{�t=�0���]��JؼV/�<��:cw=_ᑼ̷��P��<��x&y=I�e3;���;�FG�{��^�7�d�s�����g�<u�<�O�,�<	��<��=��=MPٻ��E{������l<v���B�=5W���K< =�=e�{<��P=�e�<jd��f��G�<�ܼ��x��.P<��E<�_2�iXS������u��}��x��I˼`Qf<��<?�����R�K�<��=	R�����<�J�;�n=;��V�0=�� =WQq<T[b�T'˼�=����,�%q<_4B�a�S����g���;��;��4=���&�< Լ�=z� <�Wn�W3� ߼��^<S��Y�v*=��<j�8�5�%t_�V��<Bj?;����?k�{A'�oj\=� ��\S!�t(޼8[���W�<� Z��d��܃=o��<F���P=ptu:��:ʍY��;=FO� ��8Fz�E=�[�<���X=�K	���%��R_�=)@�=�H=�a<�fT=���n�=����!=��*�A�;�K�E��w_=��;YNF=5��:�,(=��U�'�=g<r��<�A=S�|�竮�p-=�1�a�P=��(<��<��C?=y2����.}E<�,��x7��(5=w�<!�_=ƽ-�űϼp�K=.BB�0e�<��b=�(��]���R=�D�;1¼�׻�L�<s�o��n&�k���Xc<�L�(2�3=G��<��|<P�V�y�;"*���^=�2=O&���P=���<��<�sl�^�ݼG;/=�=���<�BR<�D޼ziܻ���0<�A�=>t=�漒�P�O_̼�\���-=�:�"4a<Q�b��6�����D)=s=�:,�=��=M^�ON==<�q=?h�<�-��G�<�x;6|"�EI������0K<f���� =� �<w (���#<T4=i#=Cu�<	�j��	M=�(�=�XT����TU��=��H=��4�KH9��?�Bؓ=����q"���I;�t;���=bq<ja`��}{�1=l�?<lׁ���"���G=F��;M�=~�-��+��ͪ��[�	�"�f�=��!�p�Y=8|;���<ź+�`&��&4=�=�<z� ��a=��!=��9L[<-e��a���mm�<ԉ�<R��<��;=k������\P�2wF��R�z�»4 ��W�=����k��pz�"�;��n<�ʻ�#@���;��5</&9<�L���i=^.ẟ�<��=ܹ]�R��<VG��-vV=��B<�]�<?���3�<=�/��u��zt\���>��t<�,�<�m=��=�ň���=�+a=�r�;�36����<��8;3����<,ػ�]h=���<3��<�*F����<�������"\��C�)��<V�a���<S�~:�+�;�J� ��<�C����<B�E=�60<��X��T_<�t���cB�3�h=�J@=m៼I[s�G)󼝗K=�n:�ƻ�I�.q=�
������'%�;7$d��V�<�/����T���^�$��<.�3=�6<~2[<I�=H����<��n=<s�����<`5�G( =���G-=�\��%��;�~M��p���ռo,���=�3���<�z�������s��;�%A���+=m{�<��Ѻ�}�IW�;Z���<w|\��;��
��o$�}��=�٧��C=������j;�˼��L=2$�<G-l=�=��p��{R�j�9H�:��<�M=���<l�U������t=�|"=qֻ�
��[��j�<`3Y��I=�4�<w!��y��eF;�@�<������&��ֱ<��T��1��<���<��5<�{O=��U<�q�ӗZ<�Z�<=_0�i=���;8=��q��8��,b���=� ��{'��.�<�AƼE~D�<y��\t=~�;w$;��=��<�W8�LdX�������Y=w+=�Q������ne=���U.b=P=�%T�q���Zڻ_NZ=P�x����6=/뼰����
:���<��Ã=uyM�K�<(_:=��f;m p�%�g=�3����<o�=�����<2D��'��C�+=�� =��>=��$=ݧB���)=t�<�3L�ߵ'=�:���+=b
=���</�:��/=6ky��e�<�A�<'�a�`=<=�O���q=}��<�&=�* =�~��.Qe=ߋ=_,�<�v�<��`��S�=�p:��9���&=����:�<�Q1;�����;=�Y=�D�4�(=��=� =>�;�u�;�U=�d=<�����p��|ˎ;�s=�#<=�d��Ջ��cS ���'��l<#�d<��=��ϻ�\q��̠�tʮ<�=Ju�<�o=x����=��<e@%���F<��f=}^k�<�==�L�<�=/�~��=�ئ�u~;�'Ӽ��<q���I:��z�=T�n�M,�<�;���];]nB�]I�d�+��p*�X!�G=�������3�<�n��ț��`�<�_E=��a=��`�sd�<���ӠN<)�p�r?$��)���B=x�M<oS<��7��O�|��<e*!=gl*<N��੣���B=+�)<�!������t:�Ы<��<�%�E��<
H/=fo= �=n�y=D.�@9=Λ=�	S=��o�\��I7�X�g<���<@L���r=��d��mR�)���f�$���G=�C9�ds=��������3� �<=���;)�lQ�;��ż/f�H
5=r;-����Dh;1��<��ü�yj<=�;�8^l��JC�`	�<pfj�2��<$9�KA�<k� =��-=i�8����<�3=�� =Aw=;�=!�=/չ<��R=�H=���<��w��`B=��0���<�Ͼ<��'=%I��K���!=��=��M=�c�����}�-U�;�=r���<�<�%<9��+��<�oj=M/	=�c|=�+��	��K=��G=~C<�a8���<38"��%�<����k�=����N7�t�[��c�ͯ��@�Y�qZH�zJL�߭H���==�
�nxA=}d:��H
�����5�=��ú�����G=�E<	|H���<��`���$=�,D����<�-�=���<���=��a=vQ����-��W=	��*4=mԧ<2����<b+�:Q$���rA;�=�< D�<�'�:���<d{�<>$ϼ��H)�=F v�t�<��ػ��Z��tz�nl�:Z�B���ּ9�z �<p=���<i4�A2A<�E=:�E�#�s=��޼)<�v�<�=V>,��F���>��E���������1�@����& ��<i#�<ӂ=R�F�ʢ�<4�<G�=J9n�X�3#=���<%X)=��>=�=gx��}��7�<�60�?=U�)=���<��r=�G�<D=$o=��N���)�dA�<��t�#=M=	��<��B��@=��=\G7=h��<��N�G�M0������<P���=��7��.
�q�$=�M<xS�-�(�K==���;��<ٓG=Eoe=�M��������;f<���<�^��F���=��$�������*{�i#=��뼭w�b��<�<�ā;/����O<$=���D?-����;�և=��,�#���nn�m'�">���Լ�j�<�.&�Y�~�5�����Ǻ�:���u�?! =�"=�YG���<������Y��6C=�L=a ƻ�]��=���;����=��8<w��<DJ��-������7���?=V�<Ǫؼ`�=�Jan����<�(��[=��O=�sh��t�^lR�Ҏ=Zb=�K=��л�]��-'���:v��<�c?��Ŀ��f��Y�4wi����<qJԼ^/=lz�;��q=ޘs;� �Hb<��u=�0$��o��C/<	��<,��qB��a=-�I<%�V�������<�9*=N��<!�;ן@=-;s=�.�<j@���a=`�ջZ>�ɲ�3׹ ><6��=��e�q���6���;UE�)�<N��;�o=r'=É�g[�=խ;<�b��"���=?�ϻ�P:A�y-I=0��<�z�TB���<�kq�IG=�=x3~=�c,=~/�"���H6=��m;Wc����<�ۙ<�^;=�Ҽ��ż�*.=��W5�� �4=2�(���'�ɏټu%�<_�)<
�Y-=ǯ<<N�>���x;�q�P�K��{:�F�\=�?�^k��I�<�2p�(aO�ࣶ<��-=~0��U)�!dy< ��d�	�NeW��w&=�R�=���<�c�zP/<�+���v<1G�<��;C�*={X�;A�<�Z=���|��<�N����==�n���,=�#s<�}��9=���<�^+:��7�e�/=��%��<�L�~	��]:4=�D#�Ħ�Pa�FYe��ڼ��b�uؼ�;����*��V=R�G�&={�˻�Z=�úD�=��<`��<	O �K�������DG=pͼ�%�E=bSW<c3=�7y��=ʔZ=�'*=��޼��t�}�H�`�̻G<=�J����<�Q��Bq=���9���\��]r`=�l����<{�кh@M��T��^`z=�B=#!=5G=�E�M��<��=��)�ƶ�:Wc��2��;A�μSM=l��;L���W�:=
j�<>N��t��1qu�8�<)U����+=�ȍ;wz�< pۼ�����;��X<���=6��| =m��Ú.�2j<x��cp����+\���,�=�9�p�L=�MR�pD=c)ͼ��p�`�=n�]�j9l�ɼw)+<�m;�r;=Bi&=:�¼�:���<��Z��5.=���<�i=��;p~�<D'��?��5�<�g=��#�<���c�f�ۛ��:��K=�K
=KS�4�ۼD
ػ�*^=84=������<�m<�yQ���W���6=�G�<?���84��L={�<<�E;�b�<�oj=+�=���<�v��7�=���%SO=�Z�<��a<Sy�<�U��L�
=���<%t��Ȣ��HɼrW�� ʼ�d=���o	�M����r8<V,*����ё�<���<q�A=�&�hi5=��<	�=�M�f K�� ���	=��=~=���<�Y�=��;�>�|�;pj�<4Q�B$`���=�-
��4��O��.aݼ][�:�7^<V;G=�:*=� ȼ�^����<������=(}߼]�=X@H=d99�����񇼜"T�����M=���<�}L=���7�L=�mѼYw�a
=�
��|Lt�C���a=���;jzF��1=��5=H�ϼU���	䊼2�K��_-��#�G
��_n=��[�Mj��,=�}<�����ڇ=�����a.�ga=�m��oZ������"=��9�!��������!?��Vٻ4\0=�C2��l���X�Aa=�S�뛽��q�<H3R�&�R=�̼�0���<A=+�<X�<�M=�	�<R�#�6�L=���u��y=��&�{�����;ᬕ<S �<pA޼RC7=��w<O��;��5�<MLr;�<���l=�(W�&�)�k[<w�7�H�t��мF�^�3u(�T�^=�ú�`��<�qR=��:�8q=�v<��<'l񼀫�)�%=Ղ=��<=N�"�G�N���V<��<\oU����;^^�=��$=�j̹kT���)�k�<Wcd����;>/_�[�J=��8=�G4=�����Ed�M�V�O=hM<\��>b=H�|�Z6��Y�a=��>����<�|�gUN��(����`�4��;eB�<U�)�N#=L�<�6=���=$%�B�����ct�=��(=n*��i��<e�Y=*t���̻y�=]�=E=L��Z֖�6.���f=��	=Kh�5�=�Lܼؓ���#=��5��$=-��<HJZ<G|빭�=`�=�7]��"�<�+��0���f�<'�3<U"�<�.@=�y\=�r=ݬ=�`�K�(6�ہ)���4�|�,�V�d��������q~$=]=;��y���
�	�b_7=[S�A�_=`yZ�����=b�F<L�E=֚�<pg=�:<�<��h��󇼋U��y><`N׻�6�=��b=.�9=z�=�"g����ж�<��<�g=O�=��0�!��A=���z���?���Q=6�`�D�C<]��<���<� �M֚<�<>E�����h�;#=���;~Ӏ��o�����%=Cϼ`Ņ;���R����/=�W�8X�=�K����; y<uq����껯�����(��<�bs�a�_<Iϩ��M =V�-=��M�|��<�<C����b;)�<t�;D-G<���<2�Q<+N8=x���,=Ǣ�<jy��3=�<��'=�o=A=�=T�%��܃=3�M<���+�tD=��+~���=��<[]<�@I��Y0���M�oü�|���]2=6K2���&=�˼*�F�)��T�D��g�<3���#a����)=;2=�)=6�-��8=��D���<����k��7Y=�&=n��<'��e,��ÛF=H)M<��2�c4�(pX;@�=���vp��Mh���<���-�`=����)��(h=��9=�\j����<K#��]6=ޢ��ֲ=�#�<��<�|�mV;w�w��V<t=��<�'8�S� <WwZ�W*���5;�D�;�t!={��<�T�;~�K�L�Z=�=��с<�[X�q]���>=O��<vAq=bC���,��r���n����<D
	��!����<�n7��Ь<e{<䲩�E��)sB<��%�D]�Y:�<�\ƻ�C��^;Zt ����:g%&�.v=�p=�;:(<2�z=m�=9O�:`ѻ<�9C��N���1^=���<�((�k���c�Ή���1=>$=<����V�"œ�Î �m�V= ���v�;�0<c�ȼ�j�<a��D4=�(Ի�=���F��m������JX��t1;�d=#R|�w�żX3b<�oռMg2�c�м��G=j	�dĞ���<�<#�N=��7��
QT:���;�5t<�� ��C��ܢ����;�w�^E8=�7;��|���;��O�:�+�Ƥ>���4�J\��s���>=Qs�;Dz��QYa;$� <���<�N�dh�<#����,J������D�<YǼ6�A��<!��A=��<Ă���b�<p�#�͆���-B<qb�RM<����� $=�|X�\�*�����x�_��<"@�W/=���<ɓ^=������7����<�Oe=�
D���� !��t��"���0]�q�);����7~�"�	=���<z��<�n���,�k{�<�9���<=Z:��D;xF�4� =B�޼v`=	<c�� �<�� ��o��nZ�</d�;��5=}�2���<]�׼a6��$UB<N�*�`�V��+�<f@'=�� �GEW<�1���[1�T�޼�:=�R=���<rr+�`/���)=��X=jԽ<�� ;��ݻ�<lo�;<���4���/=�!��f�;�wh=���;~��^���;�<��:7�<=��;�<��<(r�;@�����: ����N�y/�iG<�ؓ:.�3��=�T=��S�Y]=!I��Cf<��,���^�:g=��r��>�~��%�;�F�;�E�8U�O��9�4���<1ca=���e~��
����<=�+��G���+����<�$ټM�Ҽ�Z�����9]=��l��z5���g<�tX�)ժ��K=*:��92;L���9< �<�hK�=�N�Fg =^�G=56=�0<o�!���<]�f��k\=N�1=��!�Y�&��0
��� �Tx/��f>���e=W�<� ��PH�+�G���d=ޓc=��#�=�%=�h�<�.�:K=�=]\:��l<��ϻ� e<$�R;	=3<�x��Κ��n���5���x����8�Z�ռ���������B�?Lż�ߐ���d��K���I<c���[�<T�����м4_ż�%�<�c�;��Z=' ��}�q<,;H!=$�a<�*���F�s\�;%w�<�:�D�<c>�<�@9:k����#5=r+j=ֳ�;A�/�tɔ<���<�}�<N.߼'-�[Gm��6�=6��z=˞�<_�t����.x^=������<otV=Q�
�NAH�fi=+*�<��+�`�.���;r� ��?�f�l�L�=�M
<�$= ��B]=>3�����<@+>���	=t�I=� i��?���.=�m�;��b�f�o�����<�脼c�A=\�<�gH=r/�P;Y�ڇg=��=e8R=�?=��xм;����R���������[�H�R=?�='�&�i�M@Z�H�@d�<��<�S�;�I����:Z�z�訾�'=����r�<�=�=��=*===�=�HT�b�v=B�޼�+;� (Y��r�%N�<�4+=To"�X�T=�[�;g�L��=����<�	@<��<b{=�;ֻ:pF��n��L�<y�ۼ��ۼ��ֻ��9�=:T�\��<����Ƀ��2��	8�ٝ���q=ݤc=��L<��D=T�)=ʛ�� ��e<��ļ��<�۟%��߼��=�z*����<#�<�=,-ݼ�b�<;��<	���@���=�,"��G�<���;LR5=��W��-��ķ���P�*y��>R�ឤ;�|s��`�<����׈<P�_���<���<4k\�����&��8=�7=!sZ=�����]��d�a u=�s"��"=�^�;�Σ�7輑7b�t=���p�B�i.=�`U=�h�=�cM��k�<�F��0���\�e���h=T�P=�_N=�ҿ<�d3<�F�rL�zR�;��<��I=:T=}b�<�$r�#��sB�;��q�+Z�<>�ϻ����� �Ci-�Ӆ��$��4�׼�v2=���)��;�w�<J	D=<�<5��6�K��6��,-=gw�<�q<=�;(<���1�$��PA=h�t=1�.��<�FO==���M�n�H�	���$��(��y�=���;e��<�l��b»��!�⨸<=���~G��<e���<�m�<R=�����	z�ƃ��MԼ�s�3Y=:����4=�~^=�VS=��8=JOݼ��E�*��~�<��D�Ig<�^��'M��k�<��2��31���Y=1�h�x�� ��צ�;/�&<�H<=��(�=*Ѽ�,�����"�z��=�'i=�U=�f�T`ߺ͏R�"I��\=xj<Ti�<�9x��4�<s�0���1=�A��*h�<3�=;�����;>?\=�\¼h�<n(=�(T�ݱ,�Yم;�K�g�+�F�a;{�*=\��;�>=�k���<.�4�ޅ=��R��s6��\%�Nl�<1a��I.�?�B���?�t��)/k���<�e��˃[<��@��T<=8sE����;�+r=
@X������&���!=Ag��U=�a�<��1;m�<R�μ�VB=�Y�<S{��Y���b�<z��<PhY���];p�/��@�:[��6�H\�߇R� ݣ�e��</��;h�P�[B�P�`��J���S�h&|=_�W!=_� = (�<�*;���D���<������`=pWǻн���\!�^�¼�
�5��tC���=�5R��6ּ��u�C�<��9=/o�l�%=�d%=��,��Q��<����c���@;Ѳ=�?�3V�<�(��B�<"�弈�<g��<�=*�%<>�>=g{5=r�!=(͂�U��`5=�U=X ��@�U<��~�'\<X'=O����;&h=/ܱ�*�6<�8��ʼ{���V<�O<�=�Z:��R�_�8��N8=_=�9<�&p��&r=SYh���#�gJ��B=���<�}<oʆ�pD�"�1=�y���U='��r3Ǽv�+=e�=��;��0�B�պ����%�7��<ޡ9�z���N=�[s=�<!Z$�0�P=CGT�+���=z�+�b<��<������u0�+(n=qǂ<�/=	0<p�O�� ^<"`��4���P��3P�;W_��󼇉ƻ�<y�6<'�,=V1='}�<��F��J�<��:�eN<}�97(�<Y��<Ji����<�e�< �U��	��Ǽ�:�&�<%���;�W�)#�"�;��'�JC��R=�d��+=b�ȼ;D'�
���!��V8 =&6�;r�ڼ==��!�sU=�8��鈼i�����A�n��@�9<c��;�R�<�	�������*<Ɣf:"q=�'�R8�����Rbj��Nۼ���Bc=5�;�F���Q��������i=h=#����@��<�8�<J;���<5�<S�'�fVL=��R�<���ۢ���� ��m�<W&��/�����<���<(~��<Y�=D�e�d�=�]p������"=W��q� =�M]=���8%��X��#����<[P��;�y�>=����#1�J�V=2=��+=�t�<�k�=��"=����L��E=���r�I�t��<�e=�K�A}�m���(z�;X�-=J��� �2.��d޼I ����L=���<a�e���]<jY=N��<�1�<��>���4����;��պ<j8����<+p.=���hѼ=UZ=�Y����*=4�=-w�3���>=��0�����g�<=d���0�9r�<��F��|3<8�ڼF:�<�Vw�͵s<I�'<Y8d�@�����-���<�/=]���}Z=B����-g<��;g(ݻ0Ҝ�GJ�XE]=�7=w�=�{���/_���=��1��!�����8���?�	�۟7=0�)�<+�<�b;<�oK�Qd���ڼʃ�<qBg=.���B4=�r�;�ʼ$�X=YA|���X�c�m��̻��d=�m=H0x=��=�_%;��2=ΫB�v�=^�S=U��<�6I�ϖv<�o&��w˼�;ؼ��]<`��;��x<oq;���;$=�C=��8=s�V���{�b=����>�<�m.=M�����VJX=�U�pW=w��<��8��0W=���3˺�����|��fW�	2=Z�<%��<�⑼D���	;���<�H<��������f�&Y=��)g����<����k;���<W�N�uT���*;���fۭ�S����ΰ�s�i=D&B�n
Z=��<������Ǒ�<%:3�h�/��!m���y<�N)�8�� w<��h=�C1�ΉR=�5m�ι%�)��<-t��=h =�UWv<3�<<:;scE=߉p=��=��.=
�e�S��;��;��L=������:�b�3<�K���1=^^�eq�b���t�O��X4 =Dr=uۼU�̼�*=P�%��Z<<�=�LP�l����R��	tؼ�aּ�M��Wi<k*<�r#��� �ˢ��s��<��3:��V�L_׼�><<O�������黣���t�H<O�Ӽ`}���wK;��<6C�[��;0�t<�Xe��`R�����4��}��<��C�n!�r��<@�'��oD=v��D+=I�F=ļ�;�ݻA?<!��;���<����0��?��&z9$_,=�e��F=�^=�m�<��缜J�<�q,;z�=r
��v;�����=ӂ�=�w(�Z�}��g����;K�4=�[����<r�I=��d�Q�N�[���h��I���������<Au���N=e�
�zw��I=$޼�Ȑ���<J�/��؇�؞M��]Ǽ�L=��=��=$�� VE���<��3=��3�t3�����P���Ozq=*U =,
���3���̼9=�<[��<>[�<TV=f(<��y� �<���*Ȼ=��<�}��Np=��<��=kL�<NqM��r�:��(��	<Y&\=��
�5=�iP=�h<�Z����<ȟ�<9��b/=��Z=.y�0=Yb<M=�(}��x[��/��G��.�<�>I=I�r<��;<�Ы�g�=��=A(�4?ڼwI<�b�6?V�F"<=3=�C$�{΀�����v=J)����ڼ��̻N��qS=\3=��Ѽ�,w�� =�,��<E꼬g����<
���F�ͼ�=ѻj?(�(���PO/=�]:̆#;��g=g�<x9���7<������:�=$���0^=p4=~�=�@!=�=�bW=5�:�Y=;�o��=�o=��t;=�+�w�3=������B��9=�g��pp=qt<ӕw��<7���/@=g4B��@B�Q�0<��F=��=���L��X�F-=#��@˻�X���4=ٸ�<����=�����b=�=b�q�^w=��:N�0=וk���X�kJ��$�<�T���y=b�g�/5t�)��=*�»�y3<C���T;�M=<|��;�r����2�(B(�Fd=�匼8��$��?{�=�с<Q&�K$>=�<t�O=��L=�{�7Ϲ<G�K=�<|<�fZ=�Ƹ�;[]���;i�R���=Յ$<�j�<x�<{����pe�~�C��ą�E�H�È�������K=�L=V���fA��,�;�2м�_:�P:�1J�[�=�9� K�;�&L=��g={��:��N���<�!��"��[�?���?��f�=�I=u�^QD�q9P;+\=d�;�Щ<P&�<E�&=&��<�W��7d=����<g�;�|K=���s��`<b���<��+�ς/=H����H���qo���(�j��<��]=��;u ��=����a��<`��<�B��B׻����HҼ^��<�0�<�TȺ�� =�-<0� =�![�ߠ�;ꍎ�Q1M=���<Gэ<<;=(�=E)=�.�<�'�<����}=�ρ�����P=�B�<Կg�7�*=�B4���%=�^�<�ں۰����=x���xKм��F;sJ=d�<?%=k�E=-BA<���<w �<]J5<�W^=���G����b=�mo=�ֽ<�G=��0=7�<k+���c�����<ů6=�=2E�_��]0����Q�1�x`=<�Y�b�A���=EjF����E�=��5=r�<c�O��JL=	�/=��ʻMHt�lL�;�9B<�0#=V=�=���;�\��q��<��y�zI;�R ��e$=s7:=1�;�O��\/���O�\JѼ6�Z�r_=9�?�׆h��=��`���4��@���RA=��_=hF<x��<�����?|;z�<ip���⍼4��<�O��݋:w!=�w%=m��W{�<EC�<-i�<"��:�<:��<��=;9����c���<��s��pE:�1�<_AY;���w<���A$���>=�!<̎A���A=ދ
=j�<j !=ec�<��=Y
������,��Z���do<�Zڼ'�Ӽ�#U<�y����Լ���<���<���<�˜��_:�3=�v��Oe<wg=�%<g�G�k�y�8���c=d�:V�Z��7���Dq=Xa�F���Ϥ���ڼN�<��<�,=��N=�!�<�%��s=I,�Gg@�:��D=�t'<��B=��ټ'Z���x��@���$�ۃ�[B��"�m;�<�:�V���׼���<q�F=��>=$�<�&(�_�3=�!�<�?��h��M�<�5��n�<��<��(�F�}=ؼ���<GC	�t�<�ڟ��%F�J��<x�=���ҙϼɅ����w�U��H�4	
=��5=VG=��	=��Y�t6W�z&�G"�<�em���7��
��;�a��a�=�^I=Nb�<��s=�6��S=�
Ѻ�fG0=���<�f���q��Z=��<�u5=(�H=2Y����<��+<Z
�<���=SN�ӳw=�fg<<'	���<8]?;�*����12�큽��W=��6�ғ<����<��;=��<�s*���g<V��<?��-�"=T�Bn�t��<#�1=�x�;>y;Qsi��yۻ�YӼ!�=^�͹��A�+y���{;(
==OJ���@��o=G�<�&J�w>��%���0�.<�,=�_l<&��Tm=Ī<>�q�m�M=�P�<�P����<X��=�2<���;l���1�����K<�h+�B^��0C���)��=�s�<�C��|�I����=�v�\��|�<n�^�*���K�<+�w= �G��6���(=���>Q���N�<�`=5:<�9�ZxO=�3d�'��<f�$���<��=H��:�X���rＤt>�/�>=�it���;,��<��<���	�;o����=��8=j['�� ��>6�LI��������ا�< �+=�Z��==DmU��,����<�����n��F<��4=g��S�f��P���G�%z�<0��=A�=;/������=!�Q;�s_=�6�<�N���N=��<N��<s�7=�{|;�N��x�`� 6<�6<�l;��A�{�<�u�<���}PM�2N��B:=D.<]��;i�j=��=�Ή�x�b<�J���Y��߼"�}�4�üڰ��H�1<O)��@a<r�&�?��g��;�,N=���&qY;J�1�3���Qy�a/f=t�B=#�ü(�!��	><��a<(@�<��<�=s�E=�]��K-�F4��LV�:�&$=x�=o=��6�7�����T�d��;˫�<B�6=.=�H+=��[����;�UP�.������{��P�=�z�<~Z�;�M�<� =C��V��kӔ��=0�-�HR��L<�K�.��<6U*��@=�p��T/Z<�v�<&�VJӻ�Tx��̊<�Sp<��2;�,<��<�19=��缊6���\8���Q�I>=z ����s���@=�x3=�	���x�@꼍M����,<L�}=�Y<��� J=���;�X�.�=EY��"�c�`n4��ӓ<땼�ռv�w����;om�<|�x��AL�FG�;���K�='@R�����Q�<ܨ�<V ;<I<��<��<r>���ػ��;?"���P=�Ի��}��-�;ٱ(=�}����ȼ]߷;:��<;���~U���U=/3���#=ThC=�G=�&�<�,�߳)=�����߻ Ʉ�S�K��)�:e�^+�<W�
=�t��u�;ϨҼ�:<=��,=a�<UaE=<Z�<�o�<V.'=��N=�'E='�Ѽ�n=�4������l��i��#ǻXl��V=�Յ�衼)� ��Ň�:���[<��=a��<��k�gM���`���=	�QΜ�OW�*��\�2���˻��;���;ͅ�(�;�kh��쐽ס<[�?��B=\W�:С<���<7=�Lc<�{[:��R0]��)i�{X0=� �}��<k�꼐�h=��u=Kq@���I�_1�;,�<F,�;�"�<z�<|4+���<��n<�B=�䍼��?���{���������"�=��=a�k=e��<�;��������a����R��<| 4=J�E=��V=c�9��=�%W���|ټ�;�H=��6��<�
}���S���#�����a=!N9;wk��.�<�.P���<�澺g�N  ��'μ�����u"��J󻛅E=�pd=/�m=:���;��?=�2�=�YѼ�e�<�KT=~��B-	��*�<!���J����J�<�����=���;��-=f��;��Kc���<}�ڤ���M=+��#�1=��/=/'��Q;�A� ��<��e����$��=��V���ȼ���9`�=^��;H"<s��;AC�o�������=M\T����v�5=�D'<>�^�O3P<{�<a��U6]=�==�<}��9k�;%��h`ͺy,~=Q ;Tve���������.=z<W�׼�3=Τ{=��<+n]=�=<��<ء�<kR(;]K�jhb�9�<B�#���p����:����Y=,�>�&���_f
��l����<Ī=��.��H=�}0�Y�Ļ4I��p�&=�Q�l�c=hB��uT=y�EgμA��	��=N�5=O�&=���9\�<$N<�.�N�"�GPɼ�C=��&���>���M���i=��<ث)�jvJ���0=��J=N(�<��޼0�V<��<���<�7=�0���ּ��=y����O="-�<+q�<Z=�(=�r��	=�N�<���<�
+=_μ�qZ��r=��)�`at=���d�<֒�<8�h;+Q�[Ai<c�<��˼ʅº�������<S>���ټ�d�<�<�#�ѥ=[|v��>ʼ8`=8�d��S����ż�oؼ��<�^W=H3��"��B�����.Z�N�P�y�����<�S��Dv=�I����<y��<�B��{�=��A�D2�<�(^<�e�<��<�ڽ;p�������S�"h�<�]D=� =S9=���g=S��m�L=�e+=��=F�f<���<k-�<~��=�0�C�=$D=�u9=�n�<�+������Z�=F�L���O�=�U���<U����\��\���߼��<�m=v�=�޼�
缠3R=���<O`��0�����B=�l��U�<�=[_����ּ���<+��;;�=��
�
v<��;ҡ�<�=�A�@^�=��<Ū�<�n�<��<�2��`c�^��<m�<�<�?��JL��T;�s��=�=P*�$�������v�<~�P���;e�W��٦<_==$ '<#cY=�r��Pd<�O=r!���y�:(�w=e|�c��9`���sI�<51=��=-�K=�I2��:`�Z(μ����1z�ps���Dһ%�R=���&��]��3��-f.=%#���<���<��R��S���P%�����g������6�<����И��.�<�|<<�b4�
�^�iW��yj�:��;��<�rf���<�`&=��E��%S�"�ٻ = X9���缾\�<�5�<	lA������X_���)=�Y=�L:��6<��><af�<1��;�!��!DE�q?�PW{<��x���P=G��� �Y於ds��q)=�t缧�e����o�9.����Q=�M�<�8=w�e<���<D��"�=�R�<�_���N=��%<(���,<,*�7��<���s���Lc�0C��X���I�W�k�;q�7=�N=��+=QP�=�	��?��=�9W=U�<FI�ubG��CN=콶;�rT=,�`:��$=�(~�����o�qE��Շ<�K����<�=T^��aC=�M��ˣ?��k��r��<�~w���:��ּŜ"���B�͢�<)�;�zj=H3�M6�S)T=t�I�Y�:<8l�<�Z��J�9��$=��U�77���6�V�R�����A=��<R��K�=M0�G�Ҽϡ�Ϙ� �D=�g�<N���� =!.�<��3=�xX�#S<�x&.��#��{_=���<�¼��1� ��$��&�H���<�<z�;��/(�IYg=��y�eb�<�f�=�4	�4�b=�~;4C���fז��ZJ=������B��9��<��F=� ����/;Oe	=���<���f�;	ړ;��6�뮓<��<��N<i]p�.{=�s�=�$m<��m�	���<�R=�tK=RQp9��.<��N=�u=�;�s�<�K�$�	=2 R=S􅽂�!�Ft=	-:�o�h=��z='7�Y1���k��1=(L�D�$��##=$<`�C=V�R|��lg���A�J�;���<�l��B!=����B�N=�B=�)!<Nk@�
Y<�>D��3>=��J=6�L�ü.��<��;_��</L�:+��<�B�<t�w=������>��"=?�>==�ܼ��L=ߊ=!��`[����<�� =Y�=e��<�hX=4v�<��0��/�<s�W=FQS�V����i�;
�I<��o<�H<���k� =�HC����G�<�wD��#=�����L=�R=�!<���<gC�H�<�#L=�T=X�<���DP:�[:B=��<󨆼v�=�'��ۍ�A�=�缇�L=�s�,$=�b�<��f�gi=�.Y=����]��;����;U�9NW=�kܼ�}S����*C=��6���!���y<�t��7�<\X��=݋�<�:�"ǻǄ���j%=��=�-p�]y�:�dn<�"�<Y�0��p=p*=���<��������%��i(�����0㚼G<���=%�==��淍��r:=�R�<ͥa��Dy�Q;����<�ˋ����B��
j��D�!<:<�W=[��]�Q=I�(��II.����q�9���$��� =��f��|�4L=S.��!c��a<h4=1�F�9�=*�<mӼc��b��Z���=�޻|,x��'��v�>:�!�<I/���H�&�:��=爫�F
�<� �<��4��W~�'��<�S�;����<�<2M'=Y����Z�=KM�<�<t+=3�=c><��,�=y�\;��p=�Y�@O=e�<ދ�������<�� ���h���M;d�.=��Լ�=���ɼ]"B<�$'<נ=���i8='����	�eE�q<@����,�����$[=m��:$�V��1g��R-=�6��=����\d�K�B=
-#=5!!<��Z�����.���e=#��Z==�L<��ϻ_\=Wd=��<=���<%A��vʼ�_�;���;���<�F�<�S=��;�~��~=���<��&<�2�/߼~��0��4[=P�:9=�}O��Cq=�D��.S=?�'�ň��|��C��;�T��N�O=#���1�� *���<����t_<�_����PC����<�H;��<�A���+�طN���^��c�+E��7����&:��mC=oD�P	�?�S�xBQ<��==2㷼m֢���l;��=X�=D9���C=l:=8"!<'?��:��n?���Ii!�uF�;]�~�W�;��=k�df�"69=�\]=)��<x��I#�<9T=ci�(혼tH=49�ol����`;���<��#;h����;��<T��<�g<m�'���.<�!F=�1=C�1=cKļ�N ��h=X2����q<e1"9��;"�`=F3=��;=��=�i���8G�kR�=��<yb-=I���j<}�\=T�x=ti��@��&�y<'���މ>��4Y���<��d=kd�<4k��*��<Rws���K��? =�V=��û�;9<~Z��k�a�=�j?=%[��\<���= �=�%A:�#=���<�!�<>> < =S E��a¼5�a=�߆=�><Y���K~��]� =Z-�Z��<��%=��=$P3=����.=�}��>�<����I2��]�<�<���=>�<h���RcO=�.;䤑�B$ <s`'<�^���<�0&�냼�7�<�;�R���s�\��5gK�;���7=���<�G+=�=k)m=��T�����-.=�<,<��<{��8<:�:� R�\$�<�Q=�Q��ǿ��9� =g�����'*�����<鞲<�=�"�#Y�<�~1��="�g<+����<�o�;�]�^R5�$�<>=�ڲ��7���;<���$�=�t=��="͏=���;f�ͼ������h$]�:�s<�8ۼ����H_7=�!=S�0=��$��3�<����e���t5�9�D=F�D=�Ү�x�h<�22���	<�'���=��J�*h'���<�=�Ҽ�E�<ϡ]��p�</EX�~�:���;6Ҳ�t�O=	�����d��*�L�w=��C=�.=�-@�J���[ƻ�*�<=�м.<=��</��<r� �g�i=���<F��<Z�����P��w/�S���;��e�V�� ����:S�G=M�I��JE���l�2�q�~���4;��8�#0;�&�7�Ҽ�z8����<!~�9�[�<䲆���<L���=u��<�E=����1��߼E}���V=��h<�/=�=Ё����wļkϛ�g���D�_=GĦ�uqX��=����
���g����:�j��u�=;�<<Z)�ؔ=�X�K��;��6��
/��6�:���=��<p@-= �<�E=Ll�Qu;��\���J=N�:k�u��=Z��1=�`@���м��߻7��Z<!ʃ�F�<��ѼQ�;�μ�E!����$X<�Q��#�~<&=䶥<%쌽�����hI=[��;���t��<!G�<KQ=~����<� ����<�7�H�N��ޕ�q����T=|5�<�f�<���<"�:��^�:E�q<�K=��T<��U�[�<߃���>a�<陻��$<|��=jS˼�vM���7� <)k�s !=,K=��%=�p����]��<z�\�w��;�2�;�$=�;�=��D=��A������Hk)=�ڭ�Y���hs&=��<����3�1� �_�]�-0�<@��<]`�/V<u���RY=>*��s��V�{������Xi����<�"�:͂�<�P�f"��f!�#o@=j�<�ȼ;�f<�p8��D�<�k�=m��VY�<�/_�o����c�-�?<��)���'=��r���l��x�<'r�<���<����;d=�&�^C�<�r=F�=+��<�J�;	w7=O�ܼ�y���s������z�;NA���ʼ��Z=ýϼ ~B=�����<���<�����}$��~d���;z����<�
e<!iʼOۙ�%%�qTѻQ��<#�	=o:>=�6��&���+�ƷV��Qr=C=�I=��=���#�א,=ވ��ـ��֨�=F�Z��}h����;��u�]>�}{<=IT=E㲼�=
=Z����'=�8
<���'P<��e;)���� yu�* !=��t��O�b}h���<�pR���0���ucV=/i]=�+=˱��TN=�=F=%^z;yن��yK���.�<}F��Z�<�DC��3d�W�g%�u�^�l �<���<#�<4�{:9)=O*���}ꬻ��w=����-}�0����^=(�z�N�
��LV��j#=��q�-�<]�T<H�⻴�ݼ�V��.���O=Ne@��u$��f$��QB��y"=W�0=��غ��>= g����Q�<��=j��;Īl� %=1��<@�i�02��G�\<	@=�)<�/g=�M����6=0�F���
=�N�:T{�j<�.�J=�h�<�`���;�<]�E�gc.<����Sd<8��<�L>=� %=��=�~3=S]=x+*=k�c��a�h��?��?=�l��Y���N*�������8=[%�<V_�M{�<��=<2�
<�쉺9��<+�7=��'��P�;x�<l�<ᆇ=�J�<�Xc��=/�N=@5=��$��u���o�7a==�_����C=�;2x�<�IG=<� =n!=5�.<���9�r8��:��Z���j<�!�<�ꂼu�{���1�>=N��.*=f݃����<�=L��:ǪG��a(=,
=`��<���y F< Y2�*���Z�r<�����>�?��<�^=�U�<
}*���g=2"��Y�<Y�<�:a�<��K�f< L?=��)��� =W�-:+5���EP��i =�4���� =/!<�P���7=?=��t�<*�@���=��2�RE9��oo�Ay�s=����@�1�~w�=�q_=�2��S�!�`<<�4�J�<��߿��#t�(����[ü�P~��O�Z�i��;�<`x��(Sg�۳<���%>=��L�v���|A�<�x�������Ꮌ��,�_�3���x9 =m�C=�bI�lS���;�\ҼP�=�Ϟ;�〽�Iz=�?6���$��:=�#N=�,ϼ?�D;[N=W]=^ڰ;/K�+{�<�c�<%:p=�oC����;؍��  ��:=k;;6�O=�B���g<��=U�=�1#�럇�E?���d�Qrݼ�_U=@�Ƽ/�=�9�<���<NF.�A9=D~��
�;=��(:�m<�����Ǽa��<��1=�D京�N��؃�O�=�D��c�<���< R=���Q<�����tq=���;�&T=")������,=�5L<S�a;6�<��ռ��<\���1��0/=N�=z�g�G�$�E8�c=<xʼ���<�&�B����9<H�?����<�t�QLͻ��#<��1=���e|c<�I�*T��L�<���C�s=�=dMG=�m�����<��"<P�_�u<���<}�c��1�G�����@�=�5��K�;�qx<J���B=PET�m�<�:=�^�:Sy�<.ρ<H=����YR�<p��8�=K�i�Ī�<���l�<B�=�}���<�Ur�ɾ��"��<�Ml�I�Q=�� �.�v��(��V4����<������+л�'X���&�3��<7���j�;��<�����U���<G�a�<-Ul�n�ټD�=��<t�b;(�<e�@��=�b�ⴸ<Z�v=#ǡ<��<ߛ�;�n^��,�<�u��2.�#�	��F��Ü4='����C��j���n�;�B�<�&�������Q=�H����1;	=h�<����B,��n��M�û0�H=�Yr�����J=j�W�=�.� ��<�q˻�Yi=c�4��<z&7<}��=fg=6S^��v<kԛ;J�=����uq��SD<,�L�=02_���=!��<���<�<(=���ѯ�ǰ/��#{��z=V�!�ƃ�"��<�����?��E���9��gQ!�MZ#=(�R=�M=�=j��:�|<��;j��[ռ��
=
b�<�ʱ<�+j<7��<=�p�ȕ=[�l=���<�5���<ʭK�Ӎ=�#��¡;��H=GL
��)=V%N=uD�<)o.=���;���9I�j=��I=1.�3�v�j�����<�Q@�Ļ=�3R��>5=}�;����-s<�e�<��$=��!=[�A�o=mp=��<�/�U��K=o��;v��<�S��U�5OF=&b����<�<p�V�P�I= X==Ż��;VC=�[��V����˼/q;�j��Y�:o%=+hw< ��<�mh���3C�J��;�m�<}�j����<�-E�?
G=hy;+��<EBt�� P��a�<o�:�P伛�L�	�3�`��<%�=1�<��¼6��9���?<�Q�<�d�xJ�:���Wk�'Ny<<B<}�`���缽�R�_�{=��.��<�żAY=d�-�Ә���2\=$��<2��]�W=�M�j"Q=l�ż[dڼ΃��=h�^��?��d�>>�r
<��� �=�Q=0r<�����t���E����<^������<��3=�>�<e�-�?�<�6=�gQ=*��<�ka=l�W=��h=�d=x�
=��2�����LQ��fF=���<u����x�5CU={�9��=�t|�_𻱋d=i��<�Q�;N�<=�n�:*5�;)������Z$=c�Թy2\�\8����N�
;:7�<�K�<t��<��g����Rd�[�%m���!<�Q�`�7�D�鼁=Q�w�]}ԼƟ`�(� =��0=x"�<�]I=d�=~�<󊎻]� =ݤ��za�;�,v����<�0˼�JD��y�:�u=�%=� =_غ��M��$�;�o�<��K=�b&=�Ѽ���U��� �;	�?=�EJ<(M$�4�U=�)i���~�K$+� y=�U�Ӎȼ�ʃ���Z�HRE=��5< ��<�(=�&=�ݠ<d
���/����^�Q�ܻ�;<R;4=9�3=A]��_�}=�ە<�"�Ψ�;��ۼ�2�<�_��
�\!=Q�=RJD���I���<{�R=Q�,c�<��Z<{|T�N�j�������t��'��b�;�=���<�"� �2=I�;��XY=7NK=�/Z=ƀ���'=�k���o����=j�=�@Q;	�$=X�=er�S'��6��6�<]dc<>��<,��i�<��C=�7=�G ��)C=�A#<��^<�B��9��Mu�;�i=�?���ewp���μn��<��8=[-��}���=��<��{�<���3�;�F�9���w=����V���Aj=�ȳ��뼆l<a[�<q�<�z�<�@5<�m��v ��UL=��8��G������D��Y"���R��W�<��)��I��Q=w�S�2"=�K�<�<��'B<u�<D���a��߳�;� �2��D�;�bS=C7=�2����d2<���@n<�����߼�֍=�H�7F�́C<I�$=�%<�\��LN4=�0���ME=���A���a��<��c��֖�I�R�1L6:�-�<E�P=^��Adۼ,^=4��<W� =;�}�Ĕ�<#�W�D��<�j��)=�����Le���)�,��<צ_<h�J<M;�cԼ�=���Z�4�f��Hn=Н'��`�S�L�j\�M=�eɼ���:3�Y���8<R�c��E =/�:�/=�v�<G�P<c!�Qͼ���GG켨@��^A��=ԨT�q ἕ_�=�!�<�K%=��1�2�J=�'ü�{$=�wQ�ts=�7�<'�\�4n����<���b�<��<�v��%	�:��<\����c�v*=Io�<R�N=�Ϻq��;�],=�d=�ӆ�OhX�N&+�]����c�=�;n<Xe�<����<g<v��RN��-;�w׼[�$���ռ��`�t�<0����ͼ�G��V�;o�<5�<��ɼ�0�K1=-=���;�6=o�������L�=F��C\��;��'�F�<1u*���]�ag
�߫��տ�di���<�N=-�)=�2<=n�E��<��'<:C
<�a1���=���A�"o=��b���<��=7H=�X&���W=��:<�2W�z��7KN<צ?��`��%ח<�`b=s�)=G95=2ʉ�.&=^��;L��<�� (�t޼Zv�#�f=��e�r��<�K*��+%��K�Ć@<ml���/��J	=n=s�M��a���&<g�;۴����\��;�4=�ؼ^X�<J�1=$َ<�Q=vp1���=Cל<X��7��&v=$P��5n<MM�� =��0=�.��x�<��-=f�N=#�R�b�;��uJ���J=���*X*�-j=5�y=�\=��<s�Q��e�<�����R ��l;�o4=V�;*T==oI<E<�;=B�S<d��;ߞ_=Wa$�#��뾴���S�u4�<�~A=��¼��Ӽ �<���Y=��ټT�;k�;��==�
��am=T/`=�~<�UW=%gU=������:�\; �O���=�ꗼ`{Q=�I�;i���+S=�.�S���.���2����<��Ӻ�<���<>$����<!1�kFM���j9<�]:�_�B=w+�<W�c�o�%=���<�:�r+�: V=�9�:�d=ԥ�5�w<��<�R�`M,<W�˼���<X$�<�%< 
*�A@K=܄;+~Y�oF�<8R����<RX=}]^�B��W�=�X��(U<�}<	 &=a���5Gq��=B�d����<d0<��I������3<Q�v�A����;=Y�<w?=kf=rF7��~���%=���v�|�b5��E�<�ܮ�T:E�&^̻12����;�m������7�n����<��ż�ya<�]J���,=�(V���^d&��K=d廨�Q=������><��g=�� ����[�<�F�jq�O�7��l�<)=42�\�4#e��=��1=:Ï<#ƌ���(<����c4�ȷ=������x;u=�nụ�><w��$d�<�N_=.�>�̒ռ������iH=x�#�6s���:b��q�s��R3��v<�\�ݞ�Q�7�V
�;mm=M�A=Ԝr��y+�H��I�;Ù�<p�<��"��>x=j-���=�#�A��e\:���>�)��r�C�
�<���<��<�-|<U
�y�$=���<r..�5�;�*��;��<��-<�{��ۦ���\��X=/4]�/0��<d��;��=3d;a훼��7:�"�;��»4��źx���=<��o<��澀�;C�����K�<�_8<�����<�z��h��;�<�U��!�:E�<�p<7KN�l�9= �,=�%���B��:TP�<��#��(>=��7�|+��9�x���=?7?=��d<�a'��g ��Ѷ:P^�?�(��M.=o\�<)s����O=�|��΀C=?,=��g={x��#�M�J=�� =��Y�e����󍼃�L=�0ջl6<=_w�T n=�ld=�°;�!>=�T>�$ȼ3
˻�0��6��F���"�^�I=�wh<�#=��ݼq�]<��*�%�޻I������ۚ�����Ȳ�<l�>J=��<�鼀����<�N-�n����~l=���xu�<F��8�p=	ܯ<}&�<����i=��V���=�j=]�D��2*:j'ػ��<��=��/=������<7	A=�{���K�<��?=&���!��<ƅ�ej:=(��5{=��Rh;zr�－Xv�\z��A"$����;���<Y��<.�=A0=�-I=�B6=��n�N�+�D�V�њ��ݵ<}� �'1=�/=~1f=�#n=���;�ʴ:�����q;٩мQŋ<N���ڼ��=a@=T�����<���;Qʝ�Ϊ�<�I;���:U�k�n=y�=;����==j�=�	=s����ڻ�)�=� 1��)s<�\�[1�����;]�<hzc=��Q=<�d��=%����Ylf;��!�1=�`�<ՁN�+gD=�=�#='�ʼ�+�<R�=��ټ�"O���>�� �P|*�ϴ;���Gܜ��-f���<(��p���� ������㊼	����q�8=}4�<v-@��E�<p̻��Q=:*�7����.�;Q�F=l�V=�+<��t�:h�{�Z�*==Ѿ�Y=����h�:��<-��<���:f �<�ڍ<6n�<��^�a�/�6r��r:�����<�E����6�ߺ�-���`�Ʀ�⍃<�q�<fiB=��J����;�����߼���;w�n<�ބ<�k�=���<��׼�<�=T}��y�<,�����	<T���G�<-���\S=�{M���<k*;��3ɼ�샼zF��{���cA�
��<i��<��=�sI;K�<�\=�|���+s����e+��:=Gg����<����Y[=ŧ��o=��/�[=%N�~.w=U��vi =>�]��Ѹ<t���B =舌=�机�����=G�Y=2����<���<mڴ<��<������<���<�s9<��{������A=uk*=�$��-d�]�?���;�|�<r�g�#Ż�6��Է�<9�<���b Y<�6�:����<���eI�<��&�;��<�����Uo�<�<<;�B��\���G#=z���"=]`=�H�<
��[=m�w�m��:��yz���-�K!���(=�5=[�}��=GK4=�=ǎ�<W<��D=�F��c��<,:�$���;�n���=�X�<օ�k-`<v�<Z5�i��S=yO=
�Z�����Vf�^.&�G�K���|���}=�༼��B�{Dռ�W����\��qQ�7G�m(#��<��<JRA=�=�`��d�KZ=��Ul�өǼD��.�=���<�=��j=뚨���<Lh;�*RR;�*���ɜ�����d�!=�%;�uA=�;��^=w =l$�� �=�e�9�<c=����;]���k$@���ڼA��Ӿ�<�Z!=��<ȟy�Aqv���t��	�d�
����<ҟA��H��I��Us����<<����i�w��	�gT;�`�;It=е=�=�"��m�<,?<!��<�.=��n=a�"=�c��h<��=r3�$�;�G<
;<��>޼��<�B����=�F�G�9�v����<�v�'�`섻��1<��f���|����<���<dl�]��;(��F=9��<�;_�8Ǖ��<=�:a<���Wa<��W=v�4�8�Ӽ`�(=b0�<辖��S��"�;88O;+��;�O!��4
< 7=�S*�I�h<9a=h�=�wػ0"��tnԼg�a�]��<򑢻�>�<�H��}2=%��<3ў�Ӯ<L��<v�7=˥=�
G����<�V1=t�Q�?�(=,:�:��M���h�1�*��z�UK�:'�_=��<o�c=ǐ[;������
̼IYȼ�a��pX0��f�<�����=U�+��I��F��;�ɋ��&�;o���vr<J?���ۼ�};^?=(or=���F�O<Q��@�]=�fs=����;=M��;�S<r�=[r<	׼�瀖��#=:ʹ;�"Ƽ�Z<!F\;J�=��;������ ��^�c�g�l�R��;��Z�;��e=�Z�<�r����s���F���<��C�&ѕ<�ˋ�!T;�&?=�󼹀&��rD���)=/)=�m1=�(=�-=�pڼo����Ի�6�蝩�X�<$�=�ļ<��O�غ��o��ѿT<P�T<_���w5��+\����<4w׼���@������b!��/�<𐵻�j4=��	<���8��=��:�:8��}��m���U�;ex(��6�<�NC=���S���^�<B�=�A?<��#�:Y=��;�y�<�d�m��;�~����2�/�=B��귦<��$���p�d>�<h����<�蹼9f�<��<�?����<�!L�9��={�\�.�<�a =���;�䋼�S*�p@M=�����v�<�,����<��6�ߛ�Z��<}�1=Ƥ;�����y=���B���b�<�Sk0<��B<9x�	\���&������l�<���<���� =e��<&ԯ<�[/=�q�<�;|5*=g㘼�=T0ϼ��\��'�;8j�;T��;)v���B�<���yR=��=x�����(����;�]{���<pX�f�;���<68�#]=ٯ =)-5=u<=���;l���h諼m=(!=Z����3����;;xA=GRE�;�1��>[;e�q��b=qWw���4=��*<�a��T��=8 =V)�<4�j=&<7�\/=-y�<x�<�������-J�m���7�;q~�<+�U
���P=C���s7=�ϼ-P(=~A�=��<{H���;��=TU=��H<VT��ڼK����!<��r�����OY�ngҼ�� ���ͼP���f�
=c2�Yi=�0=��Ի/F��)7���ּ�K���H<�C=|�:䭺�!���v;�$E=�n�<_�:���F=a�<V�=5�y;��	��/�Ϭ%=��C�u�3�� V=�v9=VF�;�Ǘ�Z�~�(��<�+='�μ�wy=56>;j��:��:=ED��F�;�Ο��޴���v񆽽�û^��e���I���<�
J�K�<��3�_yc=�����B�-8�<v��պ�� <
_j=?=��/=-؅<�t�<2���#2��'���^=�������8��K�<Nf¼����[�=��a=�ҷ��]�<˳<%�C��p����%A���A>�<�&Z=�[.���f<�g<
�X<C�y=�+��D'=}	v�W�t�4�Q=&�<�Γ�z��j$X�mGA���(=����+༫]���Q��U��<�#.�Ƈ=K&X=���<m�=G;=b�=��Z8C�\<j=���W=v�)=�H���A=.E^�� �vE8=']P���Ȼ�W�yf=��<oD�=�|"= ��<xu��G==��)�K�=;v����4����<��s<���<���3�1���@<É}�ёg�w5=�6߻T(�:	憼"'=�Ӽ���5N�<�G�R��ן����<:�ɼ�
J�`5��F=HQ�<�gQ=*��P�<}#�_�n;���������E<l&�;a�ۼ(�Ƽ���<w�H���N=�P3=��<�jƺ��=5>����<0Q�Z-�<������)��o=l�j=׀��6��U�=�A=bE=�OL=�w<=n�=n|!��Q=Jk<��D=,`�s)c=xZ�QƳ;k��<�҇<��<q��9F�1�f�>�[�M<W�=� e+���+=|t�;����u=L	�<ݠ�<��:������;)�6<nW=��.<D)���==��E�>�o�<~�;�z~=��=�Һ<9@L�h��<<�4��<,9I���h��a(=.�;=~h�v�<�F���y=�Z�<������lu����2��I�=�C
=��0=һ:j�����ļ�B��KM���<]�^<i9��#@=�t��o����¼p.=�[�c�<	d�<g�)�4<0���q=J���c�M=+�<�<&=)v=NS-<P��Y.���ʼ'=�>���U�<
�t�5�<��<a��<6:���<�f��dt��@�<���<�VY=��#=A=K��<���=g�<�%�}���)H=ǫX=�V�=3�ʼ��4��jG=�D�O"S=�N����ǻY���0A=~)7��=DD/�)���N�M=2�?=l@�b��;@靼,�<>ƀ<x�%=f#�<��7<c�X�?𦼤b:�g�)����>�a�_=��
��d�����<��C��\^��S��`=/�A;'�p��z�;Y�3��7�<�l�<��(� �h��ռ3uc��+=��=�<$=q�:<�hJ=j�n�.�b�!B��o��t�<�:?�5=�L=�.˼�o<=��<ŷ:=��;��<�Tۺ,��<g$� �V=Ę�<�-�<��<=��
A<_/=MyŻ��=11���H�d��<4=d4=��e�m��)��Z<��K==˰b=c�ټ$]�<��|��!�A�U=�$�<�-k=�*�o���z�;�T���Ἇ��<m���i�<x�P��|�<��K=^�;��H��2=w�)� ����a��)0=D��<�Gڼ�oN�C6!<~A�<��<�\<ihV��~㼶C=U-5��"w�WD���#=�?j=����m҅���W�2ֻ�Ì��~�T=�2=A���vs<p��<A�j��\=�#�%=������=(�d�/d3��[�<�� ��mB<�]���뼎��E����3���4����<��=��.<�S�����<�<߼�y=`ʼ9ռDhJ�=;=�b�<��;8�K�2D?���<�K&=75u���<R:
�s����/���l=�C�ӝ!������i=�L)=�כ<�Q�bD�k��!��<�6��?Ǽ�Y��<C�κ%=Q�r���;d�<�
<�9= �d=�K�<|5ļ�o�<�F� o#�C�����r������	=�#=�b���W�;��?<�L����1=���<Qi!�TE�<*lF�^+�:�?=;8e=���1�����B���2�<_L�<�	=��=u��s�%�(-��b�|���{����.q�vLg=�E��8Լc��U��=�����J���<�����b��n=��S���Y��>0�HY=��=I��$@}:��]<�P�;eO���A���><��<�s�:���^y�<�E����<�n輰=.�:�: ;(��; ׻7�< ��<���<��D��)��7ؼ@�=O'�<1n=47��Zw������
<��I=�䣼�q����
<�G��<.�e����K���\�Q�ռ�к;�Yg;�x߻W!�;ll1�� T���G�A�m=�Bp=��j<UT�zf����1�T=&�����@������=>�7=�"���ü��<��Q���<}±�< �<��~=�@A��d*=j�J�;c<��Q=�S=����é;��S�F=��V�����w�<�H=��'�޶��=�"���=Ub�<��#=u �%UC�o��</C�<�����4=* �;��g=OkG<�*��E��<ňd�������=Ӹ�<�)=�</	=,��<�Q=�f��9$=[��:m4�`����$E��>�����<���9_+_�X4K<C���_A<ȝ=F;źX!�<&�}�3�H=f`;��$��R,�'0�<�<Gc���<ǿ_�-��<,���f�< ���� =P�<�0$<���=|�<��>=�"};sv=0!�<�x\=y^X=�5���<�ȻZ�\<�bv;��<��:O�`��<M0��Ɓ=U=|=!=�Zd�D:ɻ݇�}��;y�b;���;ް
=gDN=Zż�5�<�?�<D?�:���;^��<��+����d|�� ����Q=��B�C�Ӯ^;��B�h`=��<).�Xs@=ڀ�<i=�^�<�:2<�*��t]�lO�����<�.�<�1�<�<���<&/<7�d�/%_=F	=�<@��!==a�;aȌ�	%=d��<b(]=��z�w�*:�*t;M꺔z�p��\ Q��A�<�w㼞�Ҽ������,O<�V��D=��¼�.=i�Y��#=q�b=�L����=���<�c��?D=աb��ي�JnB���@��==O�1=��)�T߸<�>��9���L���T=��=9	?����R�U<�*=�:=��<�03��K;un���V<�p�;��;�h�<��<�M��o#�<��ȺE0���\<��O=;�=�7� �T<���<ϳ�<��p<0�@����<?ێ�˃H<Ψʼފs������;�t<"��U�9=#�g��>��:o�=���<��=r�<���<ʼ�<QZ�<�Y����<�C;�L:�##�;?/2���/<{����J�c<*��\�,rE=���;n@:�Q:�O_�djX=pR=�7�B�<�͚<0�h<���<���G�&=k�<���:�W��JR���;=��)=&�[=ا�<�'�d��P=5�v=���<)>�:	Z<�,�@x�<�����X��Ao��Ƴv<�a �������;^K�;d��<n�Q<�媼,���MT=D'L���.=�4�~}H�B��)�2�4K=<��r̼ṝ<᪔<z�<��G�\$�4�r�)�<+ ��	��/�H���=U\,���<G(<������iļ�<V=��ֻ;�;�3���g�@=����j�+�-=���Gΰ<��^=��<�Ί���%��F�����<�.f�����S��t�=%p=��:`&==3�<����
��U=t��!*�:����'d=�y�g `<t�'��cB<����q�k����<%�=E���w<!�Ǽ�r���M�"f�<�NY="�B��v<���4=��&���E=R�=w�=3��<t�<��U=�0D< Z�<�=o_�;ު���k=;�Ĕ��LP=h
�;)�*�{s=�+��}�m=�ݴ;"�F��_e��j�;��=���<�x>=�Տ�<D�<�=$MX=���;�62�O�Ỿ�W�9+<�U��Sh=T�/��3ϼ�0�Ͼ<��=g��<�`	<pyּ��ռîa�eOq���=1�����;�O¼��!����h&K���G?C�k�����;�������4��<><r��;����;��<x�e��A=5���`�i=KC��<�a�0�9=��R=�aW�;٪��X�в�<�J�<BLf=q�@�=�ϼ��M�����N,�bn;=Vʁ<2<�<=
6�[$<�8^<9�=+hg<-��<�	$=�B�<Ք����`�P<X�=�?��	�	=�=�r=i�\���=�<ˁ<1���3Z<��T���<r+�;N��J�Z�ǾA=�8�<D��<��<���<u�0=�=3���7X=0=��7��Q����<�(,=���=o��<�QE;<����)���0=�A�I�;�D=\��<;�ѻo�K�#Q<��h=D��;O�(<\�q�����[����i�F�RT��"�40=��ۻo<@&��}+=�D;B�/=Qڍ���F��<�&���^�<��8��A;��0K<8�<������<�/�;a�v<�c�;�C\�G����K�Y�q;�x��|<N8=�å<���;K%<y?��\���#��v���Q� ;��?=p�)<�~y=:������<u����w��Dt=��~<��H=�e��\���=�e༕��<�ڻ��.�d#=�쵼�ܵ<\ҏ:�p�;��=�b���*c=��7��=lq�;A�e<.bB=��=R2�<��K�a��p��<����4'�tPI=r=�=_�=�Ml�+,#�-[�j�=��V<���<���躱<�Ӽ�T=hnм |O=/Ȁ��	!;n�a��d<}]=��=u�
=���<i6=a~d��򥻿�.�ui'=IWi�������<=<_=�3=R�9����<~+�<Vr�=�d�[F$�� �w����W�����@�.���+��-�;(���ZW���b=��c�UpQ=U��<�g�@n:=a��<��:��<]�q�:H<v5B= ���/�<����`?� 	=Al��0=�`_�(���\<�D�X=�#F=}�f<��=�Ջ��d=�[}=K��<�J�<�'*=5I=4[��긺�����x���=�����S<�P=
+5=v��<�9�<q���M���p%�������!<)�I��!������/<��b=���;(A�<�>N=���UI�&��R��<����f���a<�l��-0C=7����߼��o<�C�<"�ݺ��<2��<|�������aH=�3���a�(�!���<�����h=�,0<h=�<=X �,f���L=��$�,:;�)m�<Js��Q���!����
�C�2�S-м>c\<���<ex�
�Q=��];��'<�6;�q0�s.��T����޼����-��<>�<
pP=
�
�^�S<�a>����qB�<OW'������J?�9��<�p6�:��<��K��3=�2ռ���F�;`p�<K��<��ռ�/&<s�<�qG�;顼)y{<�J��K;=�%&�H�<>)Z�8À<D*���9W�E��D\=S6����M�R��f�=m=���p�ڻmZӹ���=�<��8=��2�Ӎl���;X�;:�*<�L��Ob�ߐ=�[�=65��%=�_��!A�~�J�C/��cq.��4��ϫC�c�����9�B<;=X�����<^���6 �<ᚑ�ꠉ<��<����<xk7�_��<���<��^=������Q����O�}0üԶO��Wu�q��<�Gc=�_<��<�t="���̈��_x;�T&����<#=�'�<��i�SҢ<jD�<v�=x���p�ƈ8<�h���|<��"=tzW=��1��<���}��Z_0<u!y<[�\=�mk�p��:Ji����^<a�<�cP��%����<�'�<P<��/���=�c=����9=��;�e�<�����ü_ |=�7B�����(=A�]�������q���GE=}���ڿ�zI�<FAV=�XY�m�N<J���H����+���3��=:pb=����c�@� ��<�4�<�o�k(�Rib�Α&=�&,=xhQ�`��y�P��S�<��7�gI�<�ʐ���<=�U=��,���:^[`=�kU����<�k��p�:�V�>'��4V=%�c=��պ�L�� �M=Ŝ���P=�����X<�h=���'EP<Qg�;�Z�T�o����;�5���Ӽk��;�?=�y^�l�<~��3�I�=�=�4�<��B=�>�u�1�\�f�d�üb"�ʄ^=T͙���<�g��>=����`�<��غ�O���qU��ّ�9�=�*=��<��R=.}=�6�=}Tܼ$�=�Oռ�;��ռiFQ�}_<��Y=��=e�=����꼍Q���[$��d'=��0dü&�;1&��y)5����4�1���O=��&�k8~��9��t0��<��j=Eƀ�tg]���G<�e<uH��˼O��<d"�w7)��gr���.=UW���}��4��\	=���_"�{v�û��N꘼�h�&NK=�*��%���S�� A<�ͻn,;�lo�+�=�:_�ȸ�<Hzм��d�=%�<���k�J�q@^=V�ռ!A�<Z=��<�=�ݺ<bv���G<�{���g�G�<^S,=�dż�ag���=��`���<��X���<�����=B%�<<$=P K�Û�6��<;��;F.�<|�G=�y��K�<K�j�X/=�e3���
=:̼.�?�������m=+d�]Y��,6t��L�Z-;;X��=���e=���<:����y��E��<�b���<�{�;�=���;����P��<�O=����\�����<5�
=��C��N�<L�G=U3{=��*���,��C��Lh�4���A߳<�����?�?�tr��.<��<9��4�"����<��o=�	��5�_��<�w�<��<���<�81�;��n��<�o���U�n�� ^��컮�<=:yz��G#=*RE��W<��r=�gw=���2�d<�q���<%��Z�<������i�3�dˬ;�}��cP=\V6=����=D�(����=��"=l��]��;�)�����͓�=�Wf�wv�<��<�5*��D�<���z�>=��0��q�<��=9���zͼS��=����={���gừM=o��<o3���<V��<x8={R�<�l	=F�<�=�lf��;���iQ�<��,=32<�2�<^y=�`@;��k�L�=�90���<�+=��ڼ[�
���ȼ�o_<���YǏ�P�4�����hmҼ�ke�!�ؼ���Mp=�_���˼B���M=t"=�v;f`-;]��<^�<�u<ۏ,��i=�'ǼZd���GQ=��ջ����6�;�{:=HN�<��<��:�7]=i�R�7T;6f>�Da�;bf��F~9�\�ʼW�����<��=�͖�;h��;@$��N$���ԼH���w�6=����~�<�V@�7�<^}K���#=��m?*� ?=��`<0�����=UB�<��M��
���_f=��<R.
�?[k���<T'����#�c��'���;c-=J�m;6f�<5���@n^=V�<�?Ļx��<^r=p�I�E>)�����_Q�^!��=��B�d����ּV�1<�?A=w�<Y�<��q;�[�ȕ��w�y�3��Ī<�����y=�Z	�S`��)_="N
=�N=����}�k�<GCq���G=�؄<?=���9�7�1Yn�̸<e#w<PW��`��<�V=�="=�9E=���������<������^��yT���;������}:����d���=�)Ƽ�ɑ<�)='��<=-�-���k��?=�G���U���<C�<,��<�G�:����T�ټ�Bһ}x<;����V�M=Go������4���;t+#��)<�؃<VA=|f<=��;���"Ȼ��#=zb���ɔ<U=���:�9�w���U��<�Z�F�*�4?"=-\���e���;|q=��<W��=�!"�i��;���<����pR���t����at�i/�<�+�<2z��t~l�=[Ϻ��=]u� �;�gt�<�y=�<屈=u/�:�瑼��+=�&"�b��<=��B��ߘn�Hގ=N;�;y*q�$˭�B%="]<=�L��k�;|�<J�<;� �+Z��8o�<E�F�Ǹ�;a��<M�.<#!����:���N��<�'@=�ai�	��<�>=�!=���;t�L��Ǭ�%3<��=�x=`y�<�푽�z&=4=KH��"�<������;��\[;v��F�+�y� =�*=;\�xP4���'���"����<w��<��6=>�YL�</�>=�=��<)�żT9R=���E�:�$B�tܼ.�A=,^� �}<��y���u<�,�;�
g��<{p��8}����<�!=#5b<6Z=1��<�$�:���=��:J���]]=�t���/�<"�E<���<&�=e�����q3=�6�<�&'=
74�q�i�\\�9}��	��<�%=�������;G<����;�"=�iƼ��[�O#�<+��<Ce`=�!�ٻ�<��m=;��:�ɼ��=��ռ��=���<�R�:��}=�i��Ey,����<�gἔl9�z{��9�C=���<y��<�'N=X�=��`<{2����=���9>=҆4�l��=�$�:�F�<Yb��Ο���"��䉼��ǻ��C��mF�5��=��<IyG=֙��K9=��=���<��Q=T����+�]�<�)?=�B�;��<ҩ]����:2H�<�\�;']��O97���N�r�=��7�ȧ���-���-;6e��rڼ��<;�׼�{���<��*< L��:%f���C=��=�Ƅ<���<��N<�d������T�M2��S<~~V=�~4��ԼK�,=��F��ZR=�	":�=�+7=�<ɗ=�Df�5��<ૼkE�;�m�<S<�;��Ӽ�<�;7>�le0�gj�<F0���λF<�	F=9t���<��]=���Ϩ����,=^k8�k�=�)�<���Z�o���Lc�W=��/=!=�v<:�O��A~<c��:�N���=�==H[
=�k����<����^��<\<�.F��D����;ma����;+��<Fۇ��h𼤑1���=�i;:[޼���<X�"=�%!��b'=�4>�X]
�U�@�|�d=�=��<;�z4=�P6��uJ��9<�ٻ���<��H=�S�������x�=���g=B8����<�μ4g��_�Ӽ��Ҽя��Rp�;�w2=��:=�]�48˻N�@����<~W�<Dvܼ?	=�=:=r�N=ul=sN��&2=���<`5��U�:g�:#�&�.��<���-z=V!��:�63�a��;L�;�f�<Kަ����<��^<RI=��U:��<�.=��=�	=U�^�����O���\�VhO�p.�H!�}�l=��!�y>���¼�^���v�<jD�J=�a;=��O<(3H�8�<P��<g���J&��.�<2�^��A�<�o�;&bC=U�;;�K=�G`<�d=%�μ����,7X���<�5�V�<��=H�=>���x��#=ctG=Wv=!k��<8��SX�;���;_>ļ�86��쉼G�=/�V�<�w:Z�<S/=��I����ܦ���H6<�5N�c�<9]��b'��L=�ۼY�E<���9��;�Dt�]=�d=�ӆ=~m׼`E=.7,�G�J���m�j=�Z=�'�<1����'d$=��9�MoI=7�<e���29�����1=Ӌ�=��<X=�!D�a�u��=C�.�I�f�oH<�TE=9Q�<����FS�f�;�v�)I<k��<D1?=-eN=��>��#˺��<v8V;�x�<]78=�+�Wa�{]�:���='髼�1�;�����5���E�CK�<F�I�Q�3�_�Z<Gݶ=��a����<�Rb���9;����ԼI�=��	���c���=���<����ڏ�<`����g=b]g�o :=��=:R�<���<��H=4��軼@�&=�c=��R�<{0�<8ͦ�-�ͼ<v=Э�z�S47��5���W�Ɉ����<��(< k�;�ZN��{���y�����<�
�K=e�,�;M�=2�ݼ�cP�j�]<�_<��=3�(=�5O=^Լ��b��I]��^�<Lgz<!���`�=BĐ�Bf�;h���<�>�<oY^=�M8=��I���[�4�%��tY�T�<��#�p�]�C��=I��:¼���(4|<��=�q� ���9�"�5=�dH=����V�<�J����;�s�<��ֻDb:= 1_�*�^=����%#��|;=I� �|��\��<������9�h=*0�`�⼂6}�[��<	
"=�X=[��<��5=��a=��<���;�U��6�`�!��L�<�&�<�=�2I<��=� g=�|�;�k�;�¼��+���6�d�=��O�;�<R���8!�=�OѼҔ�<b�5=&��<'�<S3��μ=,<���9]!��AW<�C���q�<���
�<δ�����<����k��-��<bb����A<J8�a���Qټ>%8����:ټ�;��}}<#v�;lN;j��;�_;&l��4��mR���=[��i�=��ǽ�<A���B�<2,:<��Ƽq�s<�w��I�;���]�2�Y�7�
<0&�<�V=e&=!�?�� ��6ۀ��I��,.=p�m��R=�Z��I!�hE�<���<�]{�D�R��LB�=O�^�o���<�[�����<sjL={�=Ӝ'�(@k=�S�<������<,ť<Հl;~�t=u��;P�:�%-<�3C�i�ռR<<��|��k��b���?<K =�;���Y=|��D<e���q�<QAU<d/�<X^���z��ŏ���,=�����2�<�>V=�j=�Li=I;���<�Q���@=U�< ��{	#='�����(��p�� �[�9���/�N�-���=��=?�5=���<��8={�{=)��;T$]�$yO=?U<oo�<�Օ��6����<)�=��ռ�K"<8X=�+0��o�;��V�<��׼vg�;�kG;$�X=!����Q�~�?=d�7�0��,6=�<h.�=�<�4��ϺM4=��nd�J���i0�<�`����F����Y�<��U�����vW�i�༴��oL��.ّ<_<�<�d�<��;Ump=�=^?Y<&���E=j�c<�������;���e1�<��O����OuüG6=�><E��<�������<X1<^l=,���K��OǼp���"�<?�`<����<���U��}����<6O|<�
=U�R=cu����<���6��	 =���<5u��o!�_�<mEռ�� =�+�#�e=~�%�8m*��E���=��q=`�<UC߼�>=�<XwL=p+�<�����񍸛<k�j�c��<77�<n*]���>=��<=���u�?=\BD�	� =��<�ȉ�l��<��=��ϻ9�a��$&=��<�d��Ly�A���eaL=�Z=ޣ�<����)�<X��&�[�<`��I<u�H=�ݭ<��n����,��<錠<BG�P���H�<N��X����L�i<V�L=Ƶ2���,�2`;�W�<�{�Z�u�^x�<]�=�O)=kmi<K0�c�q�_c!=�I=���<�ZH=�	7<.�B=�$A��o2="��KZ<Qi#�=�<,=�%�Z� =�ּ�D=�?J��-I�����V�w����~�<䯜;�|ϼ�}F����*C=�d޼�Tq;%`=r�^�EN伯c���=���<�E�:�k}<��=b���#�����ĊH�*��4���M�w��C�߻P-�
��:Y�$�S䡼rƢ;.u=Čn�qvt;x��<B�<I����F-���J��7)����;ڪ��}e=���<
?1=�q=֭ջv�ۼjt(�Ό޼�s~�$����Z<A�<c<�=k�Ǽ�9=w'����<��@<�m�:iH%=��$=�oJ=�"&���!=A��;�Y�<�� ��<�D=8��
yf��C=œ'���D;��9�^+O=�"#��J#�a�$<b�5=K��<n�"�b<+���r'(<p� �J2�6j5�1G<q.���z�B��<���;�f)��+<k#�<�ɼ����R��fD=�K��;�U��<�7,�׵��e�<Sp+����� B�<���<(+��&��>�� =;��<2XL=)n<]0��c�f���w����<
�,�ʀ?���1=�>�8�N��"�;�<�G[�<��;��=r�d=��I���(=��;��n��[�w�>����DS==�W�<����<�Ā��x��=u=a,5<2u����;�7��Me��?�<c4�n\0<3=��k=a-��y���x=��ɼ��<=I~&=�[�<�~=8�ἐ�J=ie4=��#��W8=�3(=5 ���1=#|���+;f*��C =��>=�$=z<-=LrT��ԅ�:*8���Q=�
F=t�i=�Y�<jNX�ҿP=�3w<��<��$=��U=�.�<å�<��l휺�J
�]�=��/=�>'����<#�.�<��?�E�#�Ț�;�`�6�<?d��}�<�C
���K�9gZ=�Z�7Ҫ<=a�*=ͮ=Ks�7��;�h)��qռ��R�J�r=��d�=�<=0=��6���<Y�w����<�_;Z�=~m= �Լ�lD�*�ֻFA���F=�y��z=�U�<�"/���<�� �ڲ�<>(�D�'���=��K�;�*=n3I��zT�$ ˼\3,=�aS=��<�̼�)�<o{���%��?=�C<=-?u� ��&�����< �P�0d�{�@=�}=���;�;�����Hl;7=-H���2=��~=<N�<��M���vMd�;��;�-����<�����<�w_=8�6��"����:9�<���q =+��.=D:�ڼ?=�ټ4\=غ��%�+=�`>����<�����=/˃�D�N=��<7�h<��&�	��_2���)<��=Ft�o}�<p�$�����"V=�U<Ep,�Y_�;e�g���Z (��[1=ޙP��#=\=?&�<�m=\jl=SpE����<�0G=���<����(=�D=A���)=LaO��Zw= E�؛ż�1='cc���N�^;L=�'���=P:�;����D�l;(z���W���H=���}�ü�!$�$<��W�6��d�X�"=%<�Nż��*<~�!��EE��J$=�	����oc��l�o�ڴ.�YE=yܼ��=��.<c��<�22�C�T�d�=�vJ��Z�8@�;�qѼ��y�p2>���3=��k�XF�̴�� ;*��=����-<0<��8=��ӫ<�+�<�Ǽ#�ݻ��=c=��8��5���q���đ;1��<��k�V�<.����s������Jf=E�I�\��c{���g:���}<��6��t���;��h=�A&���=H��=��0=��ܼGr�<��<��G�9���z��q��;x1=�݀<=��D�nj=�1�;�/�E���˥��%��c��糼o6=�mμ�=�,
7=AZ�<�	=9��;�ߌ<0<�<�_1��%��R���	f=�Y���r�<FN4;�Mڻ�շ;:�d�L�s�W�&<�<;=+%=%�/�	��<y�ɼ��4�%���m7�&==Ar=�,�ca��0�9=��Z=����6r�d�u<4��u�'��k=��=��=�v<6���=��Ĩ<���<�t���f=�=x{��g���S��I��#m=��(=�|1�-P��P�<��M;y	�< +�<
t��l�g��\ⴼɟ<����1,��C/=d�<�g;�ݩ<��<=qh	=��X��G]='=�%��"<�<c'=sFA�ua�<8
�;@����66=�*=�(=�;���:>���B��������<m���s�;�f_=	���Q=8X�8�^H��.�z&=Rb=�E`= �\��㹼�9Ż6xƼ��:"	=ޫ���L�؁/=��� 7:�V����]�`(�����<����,��<��=:,�J�9=�x��SFI<�5�{c�fA�<�U��6><�=���;4�(="
�Q���.�ټ���<�H=�j�@K�c4�jZ7=�J��SP�st�<懖<�+�<��<'
��p�<��|��U�G��H��;�1?�l^Ǽ͖\=����v貼jb=������<%�T�B�����-�C=$S��ybջeb�;�[=\��Zy���x��Fn=Nȼ��]��{�<yB�E5�<���<> O��_�i7=<%��`�<E�H<�e����<�pr�ԃ�9o�N�['ؼ���<����M�ZӼێK;�<�ر"��v=���66��!1�?�'��_�ɟ���p=ֻ͂�͢<'���>J���=4xǻ���<8x�<A���cUm��l=����=h�c�'T��]L=�}���}���<�(���C;�|#������s<u8�������<��n�i��]%:]�V��C �K3=�VF�P�;���<��>�O�,�.=�l$��A'=����92�'�W������Q��4��m	�<�4H=��<w�.���;=�?�b�<d3W=<\N=�x=(�!=�w��"l�Ī��v��-�A��>(=|9��5����h��=�;�jK���_�V�=��>�D_=� �	!]=�H&=tJ�n�S���<�f�;��/=g�H�;=�C���@=��=y��'�<j�_=��l�{#C=ߍ{�D��� �ABƻظ<5�h=���\/����=!�ּ�z�_D�<os*=���</�j=M���W漶xe�!��;H�<aC<���<M"I=2n�^p(��'�|h�<uWg=�<�	H������a|f=O�0=UQ���U=/�<��@��9=����i�;�'���#�<,�:��Z=xӵ<]���$�=�~#�x�==�:=��<�P2�3�$=`�j=b�X<�>f<�O;�-���/�A5=]0C=_�a��j<��=�1m��o����>=�=�(�<���L���R�<
'�́�<�*���$��<!=fʼ�!��:����Ca��45=��Sߑ��t�<\�k=�(���=<ƣx<�V�Lu$=қM�Ϫ�:RZG������M�p4��"n=6FE�v��<���;�u�<���n+�<ZW���K=�*��%=��8KV=<�9}�{��o�<�y����-/�=+�<�`Y=��=>��:��F��Gj=��<)��o�8=�ɼ��R�bT=.���O\��ݻ��`�%*<�@�<Tҭ<E��<i	��S�W=a�~=z5/��CR=��=�\�<�^�?�5:�<�;Y�Y=|����F=@�g�)�S=َc=��%����мH�)�E���	*c�@l�;)��<O�<�X�<�1�A_�<HW���3=�{�=��5����;��<Lh��1<�
�!{�<�<�Tm<%t='F=�BG��u[;�=�f�K�>�=�q�71�Buټ�[���/�e���H�X=�.���*���i=	��<Z���\�����6n���;0�<�=c b<�%=I�=�/=-�ڼ��3=�6ɼ�4C���<J<X"����;��
�2�$W	���T;��a�����4I~���:��=�	5=O��l�=[�=}�#=��<=�0;=� 4=�Ob=~I<�= �I�ڹ����I��Qa����<��8�v@=�v��s=� ��~���d<�|=�=v�<W��<��;�==-�,b�8�����<`O.<Ӧ$=RW1����<G�d�qa=�]�)���,0�<���<lt=5�[=S %=��='7���wW/=�<#��2z��=�<��o=�U����j�k��;v�w�칍�k=!J�<�<��F��qE=�CA�A%O;���<���<���<;���Z=4v?=�c=`�>/=��4=�1��D>����<yn�<!����9�<-d��Z�q<�=%<��Z=�zC<栠��9=�Ze�A�E�A��;����j�	���:�z=����y�C=ɦ��"���?=�����<�X=�����<W��<��U<�=J��<�_�:�PF=���<�o)<�uG=h%
�2�<D�
����=�ݞ<��A�G"��>�=}���a<
��=�ZO#=�� ='��<Jx=�]���A=��c�\ú��=�֣��׼�e�<�D~=Q6=gZ<q��<��h�9�E����[��;� =�<�w�:�Q=�������|�����<~	W=��Z����<�<.]�<l�D�����p��tӼ�.���B����<�48=�b	<�,�d*7=�o=5:��kI���<��[=u�M�v�6; WG=(�;����,�������=\��<ޜ<�H=[%@��w��fQ���d`=N��<�0=�$ɼ��</C�F�B�=l�z�A��������im��ּhJ9;x�z<�@=n��;U���6v�;�$�N�Z;|�)=C d��t=��g<|K�<�C��^=�p�9�<���<>]��xH�<����f��l��3{9��B6�-�t�8=����z��`�== <=)C��@�9S�]�\���E=<(���r3�<�n;A�3��A =�B=n^��)�N�=̧�<�f���%=qBռ�h��]D=P�ͼX����}<]uk=s_=�:;;ϧ�H`Q=z̥;�Y�;0)�;w���Q���������'�����r�:�h0�z��O�GRμ��k�[.�����k��`=�����ּ�T=n�
�h�<��]<	E=�;����t� ���ͼE�N�S�<=�����*��=�<�,�׵b<�A��R���I�#�K<"��:$h=tZ�����=��=aN�;�*�)?�Q�<Z��[�-�Km)�	Ԋ���8< (D����� =�L;N=1zC=�����1<�J���������\+Q�M�=$Q=�Վ=�ȼ}�={$=Z$C=&=Hz{�Rۃ:-s�:'(^=ԧ=�&<��<�	�>3z�W� =��K�Ô,�W�n=3�<XD<q�;�ߚ<6��
#����,��oV=CQ�����y�<�L�:��-�F��e�<�<�<��i���<J�Q�2F�;F���
=�*2���	;/ߌ�s����誻��!:ŧ[<Vx+�J����;u	�Ht�<Q�I��kL<n�3<@��\�<kx=�aD:�&<7�8���=R�3=ȇ=0�n=���c�<,�o�8<�����\=�\�;i�= j;=�`�����%�:��=ڢR=�����h��Ӽ?1����;�:=H/�;�=�ż�R=�œ<����7ʻ;j=�=��޼��q�?*7�H��G�;Q9o���p�I^]��G�w�<M�;�16�h��<��+<F�1��?���v�|�<<�S�b�=6Ll=��
"<<�r=��-=\�ܼe)5��&޼GL�F	W=����l=u�<]�h��1L=�ጼ4PG:g���Q=*�?�f�@=����<�r���=<%��<O�!=w�0=k�<��h�P-�<i|<@�,�,"=��j=�25����<��T��5=�7��T���.l��bc<F~�?\�my�<�-��i�G�������D=�d�<4 �;�m���	��!s=�%M��m=( s�RL��-'��I�����;܀�<I<=�=�+=�N���<<��&=���;h=8���i���<�@����;�����<~�,�9&�v�7=�	"��m����v=���,�C�<T�<�����j�:Uod���=��\=d�	=R�<�Gd9H�=҆=E�<��:�H3�D�`������<��ļ�t<;Y*����*����;�+��R�<�}?=�֘;esټ�(L�?'T=�Ya�՚�<m.=�c<�� =S�<�T��4=U��<;�S=�_3���U#����~�~��-)=v!�<�cK=|���
��'y<W�P� <7=`/���'=
eM=� ����o���<E��<��８Cļ�ew<�<���!�<==B��P�_���m��<1I��b/f<+��V�6=bK�<�<��M=F�����<y;W��!TK=��<�ԏ;�U=�b�v�ٓ��񉒻v���q����Q�fW}���=Q���==��ȼ��+�ȟ�:��<��<���:/<�P�;I�<�Լ�E�<X�S=�>�ͺ���]��6�!?(����;Sny�����;�c<�	Y���<6Z=W)V�r=AɃ<��/�q��:C鲼���E���b�P����;tj���O��!��=}�]�<��<�4#�u3<��H*�d�=uZ�a災�UH���o=y=Bv=�h����w=��&=�?�X�k��K�=
F�:�����! =кi=��'=�eq=?X�<UK'= 9=A�j�Z�,�j��<O���1<x�<i�-=Lm_���G=I���n���-���=Nr�;}5�<���<"�ɼj%&���=��[�ҫ4�a5�o���~_=^�<;�#=,���(=^=P=z���Y=�o�;�C��a|C=˖=�G�<Kk=I�=B�y��~=q��<����ʜ�)���fU���E&=��w�?�E=��H2��[=,�B6ռwB7�0���˹�V2<�G�;Ϗi�� =�9���d��y�A��,Y��>�<L�<A����QH���I�TJN<s֖<?p����<l=�ny<F=*L���7�mkp�5�`=N/<H|�<��2=�D=�":=N*=�3��On�����H�;G�&�k�94q�<*�5�QA)�+B����C�O�t=f�k<��W}��l,�D22�=�-�5�o;v�G=��_���>=��+="��� ֺ��=���<4�<=>�;��༬�9=�iW��6�<\0 ���"�E�==p2���K�� �=^���id��|�<vPb�YB<* :�ބ�<�@=Z�#��[�<�W����F�=�'��e3=�&=�)�@�Y���O�U�@���=�p�<V�=+<4�;=b B��֜�+���-={T]=�o~:�@�;���<�N=�Ҽy�=�{L���S=>9�=�օ:p�3�M�\������d$.=�&��6�<�<�h�A
h�BA�<�ɱ<(�4�d=&��&Y�<�G-=v�=t�=L�!�b��;� �&�ͼ��W�f�=�<��<�6Z��������������<��;?��H��;���<��F=������X=o	�	�_=�\2=S�ں���;�{=|E�܋�;��#<���:*� (K<����&6�'=.=a���+=��n;ĸ��KC=����Fɼ-E�FN]��a=�L<��=Kqʼ5+o<U)Z=�:�<�)=�pt��`=�;)��:Fr��e�L��CC<8��<oX��ˮ<߹�; =vʰ��>���nh�;F������:n=V��<`Ҙ�no���_��գ;�N���;��f����5v�ό����J=j<-D=K��<4N4��Kh<�&z����ٜ(=	C��䲯<�{��?=��r�t��c;�&Th=�R�kME=I;���Q�)�Ѽ�OC=�jn<��J<n��=�@9=�f���E�24�=�<�7�<�P׼��V����;GO�;r?.=�7�<��e��*<� =zG���O<�G��� �<Ի�<�y���6��@q<ּ漈}2:�@=�J���<e��"T��$h�	�0=�_��H=��<�G���;��=�# =��H=���7���Őܻf�9�r�;9፼�o�Z[3=�ŀ�e>=���<"��<,M�.Fu�Ċ���8[;�!��.�<�0�<�c;=�=Q�=�*=�Z�Pا�kp�;��=ܹ9;Q�p=d#�:�vZ=��v=T^=��`=�S���<d��<�<��J=�W޼%�*=�U=���M�<=�/��B<�$	<�_q=����]n�&��&�a�gܝ<��:�E=�~ɼk�X=�e=r�	�z\�^^���I=���S=��k�֧=�_ɼ�P�n缣�<��0=H����j�����bC=S�d<���ZQ��H=��/������O�<<�%<_�h�:/;�W�<�AP=��ڻ�A�A	Ⱥ��;<=4H�.h�<�5�<T��{!�<8�e�)2�7=.��X���"n'=C��:@"�<HN7�=#�~��>wp=�&���,���=�h�)�����W=�j-=b5�% X=Sr6=.�0=���� F˼�(=�E�l�Z;���=��<�w���Fj=��K<��r$W=��<M,�<�	�<]�6�C�2=4�E�%��/<L2�,�7=�y���=$�
=�{h�g�����O�"��-��Þ<=����}3=��;�k��$Z��H��<G�<���6^$=I/w������ʼ[�j���a�+]�k=O�=��;j��	�=��|���	=��<��<?]����=95�<y�<c�$����<Zv�;�����nA�1$!<T���=I�='XI=�>e�b�C�RAI=2�E�w/Ҽ	�<kx�<�G2��X�<[��;��;3�<��<ܼ�s=�x%�lI��3m5<q��<>��p2;N�ļzh�<�Ȇ<dƐ�����l�"����=�����<���:�د9�A�4/+�1��\�I�P5;u�<�_<�)��9�<y�T=�WZ<6%<:91���>=�^��a=�=q�+=�#=�P���:+=@q�</��<�'Y�)�����@�����v�8<�w=�+�k�f����\�;g�i�ly]���a<��=,ꉼZz�T��<�U�����x��o�;FMY���ݼ�N�<C+<o���1D=M�/=K��5e�g-=k�<�]3�?��7%=X���:e��N֒��9$=�D��=�=d��<�\3=1���Ǵ�<�<�'L��0���F�'� ���O;sQ����{ ��p��񼁽��9Q<:-D��vN���=й#��j�=�{%���<�a=>E�<�8�rfB�^��<~���Z��=�DU<V=B=N߼�v5=iO1=w�E���=�� =�">�w �<����M=fIu�}<֓�<k<q=�=���<�B���5=�oZ���μ:������<�=��؜ <��<5��5��9�;=;��XK?=}�2���<���U
�U���=�;�N�w��<��漒�%���(=����K��~x�3��<�᭻��A=�Y��4\=��=�n=DZ'�V�(�J��}���g"�-`!��u޼�5�<AU�֘R�_ݻ�����|p<���:�Q ��j=�jY=��=1�a=A�ֻ�^�{����5=n�<�Ƒ<������Q�̺�<�
6�خ>�?D���q��n�;삵�$��<<J<��;6�c<�n���j<i3ۼ�.�<��Q=͒�k�x���b�!<�F��+�;��\��bE=GM=	�!�6T="FG=%�j=��h�sX_:�^�����1=�w*=6����<�ؼN)p=[�:�m�k=��ӻŌ�<$pF�e>=�޻��1��
�<1}ȼ��J=��8=�VN��%M<sZ��I;���������:I���n�=;���s��^Z<�o=�s��bc=�xe�eq�]��<f
�=Dd=��'�%��<A��hx'<s7�<��p=Q���E�</W=��=?�<z�P<�}�;thd��;$=�[���i��P�<��ż8%ԺGLb���T�"�(���<��g0=��W=]� �K���;��v=uJ����ʼݲ׼Ț�<��E=��Z��6�;Q6&=������d�M	�=��d���n�Q-g=�i;��;n;��ã�<{�������ک9�3��<c���@�C<Twe:�]�0�P<!"�=`\
=|�<*�_��4���\��ɀ����Lg��=��!GƼ�����z��lr��_=��?�QL��'=��<�*�<)v6;2���4�;��n��3�<+�< ��9��<ʼ��ˋ*;x!���)��� �3^�;):�������le����<�[0��3ȼ��(�oֽ<�LJ;yoA=��z=���<����$߼��<��������L=�P�T�l=�"��u#=~k�<Vzﻫ�-<^�O�a#6=%��<a�����żO�</J=Wd�0�j=Q��<1��`1&=��Y=;*8=�q=�=꽼j�k=��a����ú��3��<%��<K�(��*��`�<#`�;�����мהm�E�7=)�������]D�h�'���āż�V�<0��<ϻ���҃�w�<��=,ֲ��6�a�
��P߻�z�<X M=qT��Yd����2��fD=YP;2�'<�l��,�G��e���=<�l=;�$��^»$C"��%=��(�w<�ּ���<�FT���#�1p$�UFi=8�o=�Y����;Z���S���<�;S�o`J=\iu<�0s=cJ<�vk=�/�����u=�p�S���l
�"n(���A<'6ݻ3L��qc<�<p� ����������<��<3��<��漠;f��Iy����:k;���:�I<+��<��~V=Ӕ<�"=�A=$�d<ز<!�; ��`PU=h�S<G:��=8�$��#g=�=#s�Z��y�ˎ����s3<fk�;��w�A��+,O=� 0�b1�<,<)���;�;�<�XY�1@=֦G�)@=��*=Z}̼} $=��J<\c���o;&�<_x<��E=38W=�#r���C<�!o=���f8�<��	�p�;��}=�]���Yμ�i]���<�\�<��S;ґ�<$:����<x��<=
�Փ�<��8=ʹG�v��"4���)�<�=����J��u��ۧ< j�=@r���W�P~M�(�=(�=9���JaO����՟<Z%"�׽��o@滦["�	4O<�Tɼ�F�����x�{������
�=z�����<��f=iL�ۜ�f-ļ���<�z�<�t����+<��=u���R�<-d3�R�C=?��<�#���u4=��|���N�o��7=� ��S'�<F�-;��ƻ̀1=�I���<�T�QhM=��=kݑ�7�ռ`��<[�`�R�9��90<��u��؂�ƪ��/���k�-@���^=àJ�}ܻ�R<;��K=�-=P]�3�<�=:a;=�@=�^4��p>��V���:Ǯ<8�
=�Ǽ�{?�$�2=M_�l�=�Gi����;��$�4���DR����;�U��-�<D��<�ܼR�=5��K�;��<�!��3<uj�;��==�6"�Ѹ3�$���?��;#O�:��$�r`��f�G=�cX=�%���;=5���@3=�v�;2�ټ�Ț����Q��f�;���<�gr���:��*���<��I=Y�[=�#A��B�����A�|l�<��=m��<:)�<ծ�<��T=b{Y<�b_�y�	;��]<ڱ�� e�!�=�i��8#��ry'=�<�<>g��!NJ�� �:�#?=u��i:8D ����<��M=��$=���<�瀼��=I�=f��:W�u<\E?���j=���+żc�<�%=X�=����(O��q�<}�K=.�����g=Wмr�/��	�<EV��_�ü},��Hv�-o�<�o��v�<�)����;�;�Y<H�Q<!���L�<�N�E1:=Iͼ �=�����D<_%��mP��S1�?,V�ckn��;<ã��A�<a�_���(=%K�;
*N��|^=p���͝
��팼�=��U��Â=Q�<!ѼJ�;��[�%��<C��;��ͻu �_V�5ٗ<�S��@1d�>XY�/pK<�D!�?` �h�֤%�W�	m<���<�h��t;<�^?��Y������:7���������̼�ƻMUI=(�#��=;=@�̼���hj=��X=��F=�_U=13�:�N��Q���/����<��::�@_��7(���d=C.��j�y<%x%9�+����<�=�j<����<@<��<�"�:F���U��3!�<�F^��R?=ˈ=1Լx>�<M�'�������r,�:;�q����i=h����cg�BQ���F=*�=�&=E� ������<�>�<
�M�_=�T=5�>=/(�[ �<|b�M��g$<9/,��mc<<�A=y��V*6=�</ɇ�' '�'@�I�a����s=�%=���K��� =����N-�<��-C}=),3<
���yb���L�=�L��?_�-F�҉�<oQ`��)2=4���T=h�1�f<��a��$���N��1<�cs&= �;;a_a=�s=^�e��8=���]u��HV��z�<��3�GA=�d0=w��<�=M�X<@�����*��JJ�.ʼ����v�>���< F�<g��;'� �GQ����;b��p +��|<|M�i�ѻs~���=,}�<A�<���<�.w��h�<�.j�`�;�p'<�)]=dY=� <Ҽz�=��F#\�|M7=�n0=��?<�=����eq!=��O=.=(�r^X=4��<H|!=�'�1�g=<�E<�ES=y�X���B�8�b�@����i����)<�=�I*��k3<Z�-�E���ҟ,�^ "=a�T=��@�s�=J�+���k���ƼNټ��O���1���$lz��RѼ��}�!J�H
��	���/�l�M������>=�=D�lFr�:��ђ���J =Ԁ��Y��������$ne���'=�7>=�G�<�
(=x�<b�4���=}ڼqy3</E6�_\<�U<�uʼW3�~���엹I��<��"�qB����<[:��s	=�T���D<��3=}��LJZ���<�#<�w&=��<��ڼd��<@�Z=��	���=:�2���==,�2<# ��~�=3J8���ɼ-Ų;x��D�&<k����=�)=�V=��=L�<u�<@�*=(�<�i�(!����=���;�6$=KoE�A` ���=�A���	�4����$=/�p�Ό�<��Ӽ�f��=�=.nh=��ͼ̞<�4˻p𘼽@�<F0ؼ_�M��T=>�=�[�R<�_V��(=�j�-b�<�:< -=M����<������$=�N�o�=�;h�#1��*rX�9*3=Wqb�~j�<'yY<�d=�[7�C0�=C8���?=s�J=C9=�x���!��X%�Ún�x�:����<�#��I �5b�6#=�h!��<#'0�)�<�ZM�,@:���;S,g�����/���<�������U�;��`��<h<��0<�ī��M2=&YY<�i�;*����r~<6==��b<�:H����<�2����8�c��<�6�ԩ�=�#a=Xh!=�p=��l<�"��5廥n3<1&�A#==��6=<���͌��ͭ�i=x�%�u��<����<#'��=-�G�D�+<�L!=�?>���b��|T=V@9�4s=7��E��~�[=m�;[�=/>I=��6�JļŝT��
Q<�ꩼB�Z�σ���)ּ�mA=�[ֻY��<o.�<x%���ɛ����1m�<p3d=,uF�p2;��<�/R��(��Ƶ<	�C��4��o*0�C�ϼtq�<q�A=E�<�ݶ��1�<c���ɔ��Mm�<D�B��N=�m<V�)=8w���cE=*1�{�5=��ؼE�K��Ӧ����<�fb�q��;8d�+]�<� =�9��a)��V�<LW{���N;ɬ<�"�;$�s;�/ =Fp�<�󏼵 ����5�GG6�=ti<tnQ�~,�����G =B�L=K(����;�<������<GD<t#�Zi���I=�A�<�7�<��_=��=�$%;��K�̤�E�)<��&=�	'=Q��Ʃ=s�1�#"7��=a{�<�����>=�G<e�$���g�<��B<v;�<�x><�ȥ<?�<a��<ן�=\U;l��|����������xh=m���it;=���J��7��<��pi�� ��N}�;=�=]���=��X��O�B)Լ�S����*g;��J=��G�z =��b��(<A�<�'W=�:U�E���g<�u;ϭW�G＼a�	=��ʻ�$=/�\<�B=U	���g���q��õ��G6��%�;�=��2�?�< Ff��D<�1�a�M������@�v��<nzh����d���Pg����;�����p$�*T�<O�<�H�
#�RU�<)��!���5S�uD=��K��j�=}�!��$��՚�;�g�nը<��Cb�<:�<_3�;vg��q�M=�d�<��^=|��NI��aH=~�u;%=��<�v��u"�3G��{5��T=C�=IL��7�[=�����<Ҽk䤼��>=����8A=]BQ<���<�c�<��9:�����/<��M=k��}=�������c�~=����N�=��4<0^��w�%=�	l�֖W�W�λ�cm��?�=��k��}j=w��h������<��<��n=�إ���=A�һF_={�ԼI�[��1���W ���D=�|�QiH=ܾ+���-=�0<���; �=�!����<7G�
}�<��#=��S��B��+�<pnI�b�0�<;�s<�Ϭ<��4�J��j(L�6>��p[�F�V���<�0����?�yF!=���n�;��<<��;�D��=:9�:������:v�=�~<�V�<5���#�==���<�֮�!I�;�09���I=B��+9޼c��I'f=�/p��ѻڅP=�94=פ�2=f�|�G�W����;I6���	=���;�])��ו;|���H����<G�k�& �����k3�<��6<��=L�'=�v��e=��}��v�=�dR=�:>�=�6�=����;�A0��]A<W��;�B	=�Լ��ܼ*7h<�W�<
�o��8-<�eμ�.��7}=戜�8I��1���hY='�v�����V̼c>d=��;��=��=��9���1c&=B����L��^���7�m�4��e[��%���;��Ҽݹ޻�>=y`=a���}���e���<PH%=�c�=G�c<��Z���:a�'����<t��<��s=+������?�n܂�a��<�K=碗��� =+s����==3�����;~����@<�<�9V��m�:�L�Y�p
5=�!��w�ӼY�O���</�L�\�="����;�������*N6��"/=*�I�-@�<=Ы�W��e�ûnPQ;Z��;y'�_B=�X=Օ_�at��;=����r=K=ǇI�7dD=���<c8=} k=���,;��<^<R=F��<�2Z�
����ދ<��<~/�v|9.z�F���=|B��&D=���;�h=>y˼66c�����Z��{�"=���k=Ϣ���3=W<�&��?��%;�<�<u+���˯�h<��g��� �`˺��.l=qg[���H���<�{�9zI8���?=c��<�e���� ��*w<Z>����<�w<þW=w�<��5�������+Q<ZLr�dl$��C=i�H�Ĺ��0�=&�<ƧW�z7!;���<aw���=ԧ��U".=��=13��d�5=����:gy��Q�=u�7�E����<�u�<V(~=>���=��:Pn�'C>�/�L=����t����<�p���40�-��35�(d�FF<�r�=o@=B�8J�;�>=v�׼��W���=V�g=��F��F <:g='�<À��6�<�D=3D'�LV9���=+�E=�����;*����X*��[d��X�<�мl�(=�D%�up�:hE0=�B<󬼘�<��A�T%޼+�=���Q�;�}�pp���q=��4=ӹ�=����=e=Z�J;�>��2F����u�k=����I�a\(�|�ۼN��;���;���	��;%8=V��F��d@o�,�S���=�<q�<���<{�/;�#=u�G=:�_=�"�<�t�N�=�%��ķ�wđ�2ze=�YU��i�<]I�<������q=�J<)�i;I�ż�#=8x�;�K&=D}�a�<���:.=�+f��+f;��==����3#߼��v�XY��5f=�b���!���v��H_���=���;��G=S:��<�~����;����
=��^=ʳ4=-�#=��/=f�ۼ��=a�6��o�=Ě;���s��<�E=M��DGI�[.b�J輆6��Y�g:��V=�D���[;`qu=縍=+2��,�����;��;S���40��G�<iC2���<=n�Z��v���!��x�<9i=�J<��<>$:H� �.>=�>��l�����OV<ֶ�;�&=Na<�	�<f�V���<��(=����7l=|�<��Y��0=n�<��;R�9��n� a=��F��`v=R�<+E<�U�f�h=�sp=��p='=���	6���ڼC��/]�˥$<
V=�<a<���<ߺ>=Oaػx�< :�={�<a�s=�n=��;�i�g���^<�x�_|������EM����p�$��T��*�	r,�۞Q=��<T<�	D<<��U=Rt6=��;y�⼉�*=nw+�xD=���B�%<7%L�ᭅ�ś��J�`�g��l`��/����<L��И����,*��ࢼh�x>ży-=�q^<�������h6<�z~��WK=�`���b�LN�}��;� =\��<؏�=�s7�/��Ж�KJ�;�ռ_�=��=��μ�����  �;D\�!��V�H
��Ƨ��ҕ�����"���N�<.�}= ������"<��=��=q���[�u-=��X�����<J�:=춅=O.�:j[B=z�e�_| =��$�j��6/�.��:$E��mn��B<@�4=D���ί<Uy�jZ<��ɹ�\r�;��R��I�o��8¼H�I=�h<�J�L;[��<�?���,���i囼93�[��jZ<!���Vf=�w�<�����I���$:�<8��<�$��s�7R��n�����r
��^����
=
K7�j=�M�)�<{�<�E="RT��B��-=㉧�;�"��d:p+=�]���3����<F����7P�k<ȋ�<�"=�:)�qi�<�A;ߘ</�=�e=���T�ż9�T��!�Y��c9���a�<�0�<��̼1v���H;�����>F�c���~U�<��*�)$���D��� �X�w �;�Ku�|N�<ҹ�g��<����L=T�?=OY�=�8z����:Ш�<��I�Eer��OT=C�U=Q�m=�KG=!*p=b�/=��(�'RG�^�⼉�6��J�;Nʼ�b�<����<5�=��"=���;=!����tw_��$�<1�h�Fq=�eP=��S�G̼����V.ü6"��T�g�= �<�~�<35[<>|=jJ� �޼�W=eX�Ū/=񜼘�=>=�؞o<���L�<q�<X�'��1l���C=p�}=�=��~�d�O�9�o�M=���<�)�A]K<�,/=��+�o��0!,=�h���5= ׀�\�����<�NR=+~<=���;	};���<�g<U�=-��]w�3��f=@ZS�n�����Cp�<^H���`=K&=3?���b4=��s�%�C=!u;=�i4��qw�4�,=w����<�*B��K;��H���:�z��c$=��V��ڻ�V=a���(�<.��<%���L�!�g�l�=.�h=��=�⼊�l�W.M�P�.���oq=�6=g�9���[=^~=�0���,"�����Ƴ���<��=��<��=G�����<����w�`=��99�<�i=U����=�G��%�=���<�a0=�yW���%=�=XK�=ѫ��`��<�?���:�F��<Ak���	g� c<��=����	��#tv=R�P=�{=*�����;�hc<���%�/�UNz<A�t�ۏK�F�E���<��:
�t��y=H�<�\;���<�m:�[��<x�<�d}���=�R�<��"��8�<��6�+���R�E;]�j�b�`�u5�<q�]�G�c���	�ę�<7
�<��ʼ��$<,�	�K�ݻH�R=�4;�8�.��󼺧A�V;T��R=0�=�N��Α����[<V9,��2�G��;qN�O����<P�H�k�=����N��G4=2��<GZ��5MR����;�K=���;T�A�wa~�R>��ԩ��Ⱥ��jw=��=���;'�����<�S�;=�I���u;�#�ծ��˫���;=Z?-84뼰T=g�=� 4<nμ�92=aKV������K�;�@n���!=SH%��<�(z!=M8�n7)=�ٺ�����:�z<+�;}Cs��^�����I=�===h{׼ƀr�] E���T=m*�%j��?"��N=�Ч<�<7��pk���=T)
�x�K���=1����P=CH[���l����K�����<i�8��~�E��сM=<�X=7�5��
�IBZ��]b�u�g=�v��x�<l7b<�V��	�z=��W��/�<#:4:U��<��}<�e=���C�3=����P��ę<GF�r�¼�o��O�	4=��<�?��B�=G�2=<v�����<m>;�-=�dټ[;]:*�_=foE=��<���98M=��H\q���3=:�<;X�<�쓼�����o�R�^=޽��u'�_��<�Z7=��=4Ơ��cּPlc=7+#=4=�7�7%�4�@=(��Z���Ѽ̲�<�t[���Q���<�x=�f7�B=zZ^��.I��Q滐吼X�м�<틉<��;D˾�L(��᜻�=�=▖���/� hɼ
�<+o=F#=�h=���:�LI���v��k��}���DYj�5O(�vC���h<�"0=Ո�;a��;��&�&�=����h�<�%p�٢!���]=G�V�
�<QE�;SŽ�1���x7c;a{�<��>�%z��\0�	1�<�"<в��T �B��<I� <x	�˹-�dX=��[=�\�=N`]=@�<��<���<�f=5�缧�d�j�<�B)�1{;�ʼq,=ffC=_�K=� ���l>�ϗ?=O��<�B���]<=�m<ó]=�P���wD���=�0�1�#���6=^���6�,=��,��+8�T�k<��O�l��Ҋ�<_yp=ہb<4�}�dP�<��1==���/=!&�`<˼<rI&=&��Q�I=H��XF.=����M_��E"�{)?��i�ۥ=u<]�I�W{�fy7���<d�6<��=���@�?5���:��@�1�h�ټ�th=�H��#�7�U�+f�(>N;�l���w<0b\=C���������`�<�J=���:��<酉<\z����:��<J�=\��<u*b<Q�ܻ� �<m�
>�f� �*=�},��e�;c�L�T!1<0a=��o:t�J�ߏ=��K=#6���-<�tN="k�zr=�|���uӼ6�R��p<�6r�6���h��<����!(5=�J1='�5=�m�=u15�m`Ļ���<��ȼȌ4��H=���<QμW�\=&%n=��/=�e=J=�C�*=��+��b=�J��*�	�4�2�>曼�b[<�^f��Żb��<���<q_O�g�H<	R�<��<^.��}޼�*�<06=F�<-����j��&��yA�<S ֺE�{��;~x��S��<��S�v>;��f����==+�¼-�P=D(h�T4м��T="�_=w>���p�<�q=�X�ݍ�;�^B�cq�:�=�E�<&�ۏ�F�]��zu;枉�2"u<��<?�H��h�<����ؼ �*��#���>��	�<U����==o=��Y;;���:�V��<ʛ�;0��<�z�<��e<%=�Ѻ�/FּZ'(�KbJ<y��R�,=��
=H�C=�O�X#4<l&J�I4�G==hi<�ݵ�8T;&=�ч�s�:��<�����3�fʾ�o�?M.=��h�T-t�rL=g��'�<��7=V�<��v=0�*���N=]�N<p�"=E�F=$�Ҽ��o<���<�w=��J=��=E� =+k(=���;u�<�V���F��B��8=
�C���Ǽ��<)'<Ƹ�<$��;�==͚ӼhyѼL�X=���K������GF�<xfǼ�g�8�W����<1�/�"f< �Y=��c=OM��܎;C�N=<�X;��;b��<�ؽ�c D�*A�,�&=/����PQ=���@]���ͼ�Z�8i��1�;�==^��~�<�/�<��ú��Q=v���������q���;׵�<��<=�ܻ��I�.`�`�,�K�ʼ�Mp�B��.=-( �Ku$<�:b��'�}��G)żY�6=S:J��>G�)�T��M�ѷ�؝<�X=y�
=̻g������ĳ<��=��;�O
��u���&;����F4<��;��
�h�8�	�3���O�TW��䢻��J=P��qݼ�l<������&�"����<��W���(=�vR=i�����	��M��)m���=w��<��<A	=�"�<��<*��<T�ؼfC��q?7=k�K�Wߚ�q�V�MC���o7<��U<>�2=ϻ`��H3��J�<ޗ>�W��<�V�]���(֨��XD����;�}%�~"�R�
=�҈���<r*��m4��B�<"��<�7L=�o=b���,j���3<��,�sd��7=�Î��ʼ���<?��$�(�G���&=ݯĻ���<�b�<��=e��<�t�;�0W=��3���=.%Ƽz�=���<�#W�Mq�<���:
���ʼ��w(��M:����<��e=~���7�"=�f��<�*�<W�<v���뼰�B�9;t�L=P����4=Xh=[���(
�T82��81=@����T<f#=���Y�N���j�o<z������2mi�D�#�O��<]�^�s�)=��t�^�g=Ý��E<���1=U�7�2�}��ּ"�~��;��=$_����;���9�n�<-��<q�k�I�ؼ];� ��<�D��#�
=؎=H=��;�����<�)S;�uI�K/=�=K���Y�0L6=�TR�1]���=���<;�w�M=g�7L���o�G=®.<�t=+�:�}O=q�=�2<��y�<lsO�XC�Z˕��<<3.=�nh�U'
�c��[�>��N=1o/=���
v��ߦ�:��3='�<G�ļ+P�<��������*x�q��Ԏ�3g!�)~���w��0t+����<�w���=�< ,$�S�<<�<�<Uw�:Gk <���<B��w&;�u<�^[�6��!��9*��fx��J=�������<���:��\=�1���G�&�`���λ3N�����|��<i�C=\���VL=��4=�Z�<�+��Hخ�'48��U=�;=��`�	-�hd�<���6z�Rft<��>=��B�n\�<2޻�S<Y����,=�z��E<�Y=�u���ߺ��J=s[k<Wg�<�֮<M^c�b��π�<N�Z��BҼ,S�'W���.+<�6���2��}%�:	s:�b�<�ҿ�[�<�q:="(=o><
�( ����Ե�Hc�,��<i��<:E���w=o�/=9r�;P+=Y�,:UN�z(��kT�~D
����<�~t��<��<f_*�� =�U�s�;��(�~:���;<�p0<�9K��-�<�o6�O�S=�W�<N|��W!�%���DٻX�=�����=��g;��W��yJ=��y^��&@`;8@/=�!�l+�0�=;�L�������;�Cn�u�,=��6���{<�}������{<�P|;p���|����d<}Қ�>AC=�R/��b`<�K�[��;�d���c�<��q�w�:"/=;��<X��$ѼH5X����<��μѠ9�睲��Q<ӈ����Tc�i��;S�<���T=E^4=XY���f������⼟��<]=��=��(=r�H�����h
�<]�e�-� ��T��M0���(��^�U:
���|��4'=|LK��"�<�M�<;%<��,<pY�=E�<u�x=�ռ�D3�lo,=�P"=��=�01<�����e�O@�<gN===��q8T��=��=�K��VpU���I=��a=R'�<:�?�ab�;M�;:��0���=g�8�Ó�<ǒ�<��<e���*"�������/��$=�ڼ�"�� �6��sc��r������֖:��;�~�<f�����V�;
�CY=
�e=��<+-�;z<�O�i e=C�v�ǧ;X�
����<k�D�5��Yt=�D��a��U:E+�<�[I=8��I�<�������#��Y>=|�}�kg��g��m+t;��=������<ɭP��R׼m��9�k=(%H��� ������T=}|�<W�~�d�~����<�u��8�< �e�a��<(J]= �D=�)�;�
=BnU���O�����=�˲��c'�ީ�T(<=��弝?��r���3�V�B������;�;
�����V�������<Y�k���	�<�G-=Ǻ�8㵼m�?=��=�W=t�ɼ2+1�}��<�2����;�k���<��ӼI���.7_�����~�p��:��9=="�%z��`�:�Ұ���&��.e=�o�;���)�:=:��%�l����<�ĺ6
=��<Q�8=	:e���<��4�-Ĩ��˅<��<�"Ϻ�p��<K����A����9z��<v�n;���;���m,�<RX��M����t<�1���I=̓��&�~=�B�����D	=$��������ļ
���+=�9=��=?��8U)��s��:2=�=>�3=7�2<i��:?�?�E���<�x���q�<L��<������=G.��Y<[Κ��Z�=#+ݼ�N@=,Lx<j�M=O�>�b� ���H�<�k<����{ŧ��#�09=� R<����#��Z���<J����<xCռ���<��P;�
1<]	K���p=cZ�<����;,@� F��^<A��<�=b�*�#5��%�I=�D0��C=+�że]��T�?y<���<��i������_��b��]����k�*俼�%=! ��+%=�:����<�4
=�#j���ռ��<ڊ)=�e=�����.��<�+�����< ���2<A����<V�=�A6=�bR=&�S:f�0=��4���ؼ�ɵ<�ܑ��9�� V�<��K���_����<�f�<�%���¼�w =��7���F=w��<���J*W<B%�<�J�����<�',�����b�<T�;�_���6<�Ż��F���A=����3H=��C=,7Լ����3��aF�C��;;�3�/����$�]�7�2=����ն{�3=)ʎ���=b�"��Lϼ�=0%��?�*���D��ß;��Ǽv��_=���<�yG�q�=��=kvE�z�<��W=K�=.�G���񻝚/=�ڼ �=��T���:x�=U(d�q$�6k�<��<g�����q<w�9;r�@=�`�<̥=ZF	=IF�<,7����d�YR/<��=5�F<|����O==��u7U=�~=nJ0=���<TNA����A� ����8=:D�<j��<ؽ�;j\�<m�w<����Q)���.�m,3���= �H=� ���oq��L�<%��']<�~ʻc�Ӽ�>M<�<]l'�h3=�����w�����.�:�*�<:�;�j<ܠ=��<�=ԑ� �V=;fX<	 ����������	@$<���k��i��:Y�v���:=��Q=rm]�8�#�nR�\�1=
��;��k��=sA�;�H�<��H=?0=m�6���<��$��b���,=���<���<^J�<�h��!���8�a�<cʄ<@�+�`�B=��A�6I)=@�<���<}�&
�@���'f� oڻ7<��;�幻1���༜<QK�ɽ�;9G7=�V�/P�<�٢<��g=&�[�&��:$�<��\�V������<u�U=BG=y��<{��=��:�0�uN��K��ڼ�s�<O,�ǋ<�q�;9T�,� ��p9��?�f�<�7�<�u�	�z<y[����;��<h���C2=��=���� �7=�Ȉ<[��Y�G���<1�����{� ��<gI¼K�/=�"=���O{��� ���<s�h����]ɻD5⼞����H0=��=&&<�����@=�@�<v�<�@ռ�v,�*+��e�Ǽ���y
+�C�=��@=?�+=,!w�;G*<~pq��^����B��g=G%$=,�:��CO=�Cl�n��'���d=&�6=�����I�M��R^���<�"�/�
��ST<(�<��;�=>=ւ��$����<����Ԟ�;���Y�c�o�<s�>;�?�<�p@= /�<.�n�-���'�-"��s�<]�=�l�<n�Y=£��-%p�����SԼܯ	����<��)=�C&=�R=�z�&�7=B)�:�Y=l$=�
�q���C<��'����%�;��⼌ֻ8�:`�&=��;!a��%e@�m��<�ML=��=���<�H���x�9֚<�c�����%f=xz�< |�<?�Q=���<��V=��;���<��=��мz|t���V<�`$=��B�6����=� =l0 �9��<�=�d�<�Sջ��ݼ�{���ZK<)>K=Gt�<Y�m;��4=��<�u=1�.��p����ӎ��/=�ҿ�<�7"��M��6=%�o�HԼ�����Ij����=�(ϼ�#@;Tl��ZG=^��c���UE�p'9=0�]��FѼ�l=I�ɺ�`]<�(���N�823�C�<�K�<�t���'=G9�K�ѸZ=_�<1�U<I��<���xm�<>��8�<��;��W=Z��<����k�<k,�<��J=X��:N*<IJ�n�����=�|@�<4�$=�ȶ;���<��,�-�c�~5K����b=x�<[��<��&�te���;��M=��R=��<��T=�v5��2Y<��k=8�K����<�yK=������<�cN�Z ���@C<(=�Cu�+ؼ��<�-�!���V�a\J=��;��{�9�BH��P�J=D4=[IμyY��sJ=�Vb=�2��F�k=
7��L�<�pY;�,V��A7��/=ܲ|��w=��<Pr�<Ħ�<� ;�+='�R��x�<���;׌�~BZ=6)j��;ae^=�5�<���=�y<�*Y=c�<	Lͼ�~�;KV3���;| ߼���<>m<=����\C/= �=�/�:�!�<8�<��;.ס�G��p@��9C��e����=3��(��<��E�Řw�d�`=��,�FaL<&9�<�Pm����;�������O�~����<1N
���9TЋ���R��
�;�:�Y=B�7��w�#]�<���<F6��ާ���@��r�����<I(=�Q]=� M=�_3=�c\=��e:�:�<��v=�м����r�;l꺼���;-h=�c�<��a=$,v=`Z=E.���{;�t\�LüF=�,&<G�)V=�?b�M׼W�����D=x) �J�b=� Z;ݗ�<w�<�p�<�T,�:e<=�(Y��gƼS�0=̷=s�޼�͌��;r���=)�6�\�Y��A�<�� =_�/=&uA���ؼ#�ļ���<�w'���Y�	���B�0X.=JXl���.�n��<Gw<��z=W���(�<3��;��t�lM��"�<�V5=��+=�|༄9�F����e<�#�t�}<��ݺ�6��^=ێ�h��,V�Lֻgȷ<5E��B���8�<z��<�"A�PQ:�yo;� @�qF�<(�o�J��;Ѭ0��Xs<|�¼49��Ŗ�U��<��ܼ�ޓ<ܙZ��_)=zn~��Q�;�HY=��a:j)�KLR�.?=���<�5;P�L=@|,<E��ً<IG=)�<��<k^=i�.�A�o�״ ���.�Mwɼ�*�<��5;ż{	�<d���ي�;��c��ɡ<��_=E�=s7^��]�Z��<�	=�ҼF�`�.�=�]���<�^	��QR��Gx��
������=|1T�>���'[=�^v�w@�<9�:��<V�=������z�d�aZ=O=�48�-=�5�P٠�c�%��H=)l=ne=��i��cռDR�ٴ�<�,'��o`�ۓ9��cR�G!�ZY=9�%�\�<^?��(�<��<�^�<���\���:;��ݼ����V�;�� ���;��q;a�+��6�H��<.X��� V=�ܼ�^���>=�-=�p������`-=FѺ<7���ĉ��.�<��ּ��;ϲ]�B�\��Qû�żfIC�)h��wɻ��#=ZA����<��<9��(-
�'70=-�<̣�<U�=��~�.Vv=]л�s����u=���<!>]��s��;E,������<a���i�<�;,�F�<���X 4=I��<־L����9��&�O*�<���:n����<-Ȇ=i�p��s�iW�<I�
���<�t�;DX��wPռ����=Ԃp�b����u��� =�f=H��g� =�_+=�&F��v�Hj�<+�<��:��Ƽ�6)=�{f�BS<{X;�-=�Ӄ<7<��9��䭼4^ ��7=�z<ɘA=�?�� =�IR=.Z>�M̴<F�K;./=ZG=;�>=ͯ"=ц���@<������ q.�@�üK��<<����MZ�hNT<�e�Q>=J'��Y9=rq��A=gD:=�2="�V�%��5=�\7�W#�r
��q7=�S�<��a�s��<|�<)��Q8�<���Vٿ��*`�:�?�[h=of=��¼S��^n2=��/�`=äw���d=帺����<�nh==<���<Kb�<jf-:S��[�g�e��$��<�J.��tl=��0��=e=���;W�b<O��R��{R�e�|���b�*.�����0<6�h=*D"��V�<�,2�}О��7����X������;w>��df=���<������ּ~�=);q=_�	�O����;�O=ET=�v=�Z�;��(U=��m=er��e�?�Q@�-�ջ3�<�+�<|ټ"���E=��1��N=?+)<.�=�>��G��� ����ʻ�7�<�8�`gڼg����/�Iy@<����X,=�Y�3-=����4�Z�C�9ld=QG/��Mڼ���t�X�"�]�5���<�S =��(=���<��Q�ɳ�<��X�˺R��F:=��]=:F�:��)��&3=�(H=1[��a����?���0��f==5�9=�K)��<�O/<��E���k�������c��$Z����.=6:7=6�m��w3���C�((�<q(�<�།�H��c�;SD�;|:k;i�Ѽ4��<r�@=�� =��<�'�<�#;0�n�Q��<C�i<�<���������;���<�F@<��<oi�;e��<��=�E��z���첼#HQ���˼%V����<yJ�Th�;�)P�7�s=4�M;�7�V�<�@��ЉI<4�;��<Ě�Ilf�!L=hjҼ�>���=��< �=����=���<�L���=4�<�=�Is��.����<!� �H�'���)����<i�<�U����#  ��L<��P=�:y��A��&�Vlq=���^&�*|���Vi<�Z=��\i=5؋�&��dM��z1��'c� ���po�=�=��SF�I`��I�N=��*�T޿<�Q�;)�C;MH=A!��D���8�?�<@��;�.�<B��%>=u�N�0L1�g�=�Wռ�����C����<�L{<-hK��8D��Dʻlي�S��1�����9N^Q����<b�"� �O}�<�ü�
�z��xyQ��^?<)i�2�W��<���<y%=�<
'H=$�%�'l<�L��m��:;iZ�<_(�<��R=�_������<Xټ��i<�R^�v��v��X<ދ9�x=��2=Uا<{�C=	q�}��<��m��	�<�.�<��"=��w�~��<��{<b .=Y:��.��<�l�O�=��#�4e��<3���v�⋅<ف�<"mQ�{5=��_<�3=8䥼>9���ƻ�Χ���=q�<�� ���=-��A���)<�J���Y�; j'=	���>�z(�<ނ<�F<���n=!=7��:�;*#=�������g=����r�m��<X��iZ�D_#�	��޿'=��(=���:��#�$��L=��m�~y|���s�= S~=C@ٺu<�<�݅�0�
=�O><l��;��<��!=���;
(��o\��SG�ݙ�;�=�X�<��<O>� �=Q�{=��9�Ζ+��Y�<-���ɺ��Ҥ;)1��V���Ê;�=��=s�=�wn�����oV��w=̷J�.��:�/=�M=�~˼ANļ8߼�%5=���=�w����=V�����;v�s�#Ԡ<t�N�}�4�� м7���'��<���R=�)����q������s���=j�<�!��R:="MT��Z���8�T��;JO=^��;�bżC��@�$�?#м�4���@Q�=�<(Ҩ�K׶7#YJ=Y�g<�^��@=&�=̜��r�c�U=��<�9c�:��@�<7�3=��;��%�A` =m�O��<F(=��"=n�r=�R��#cC=�\�<U%���`���Ũ<-�;<z��=����彑�?!���|���#=�f=.��<��i=CL��9�=�5�w<
<�v<fQl=��≮m=��"=�1�	���~;*�j�������m�>B��[���4B=CM���<�1,��Q�Μ��`@W<��<��Ƽ��;�=Ƽ�:<r�<�?��<*�f��3=��O�$���`����{��"�4< �*�=�&;�H���z���#���M���G��h8=0�����q�jJ��c��R��H2�<�zX���.;�n�<AD��a�<�g�޴��(�"���<�n<��_=�㼘�����G=�����;�<��H�����a�޼'h�6��<FjG���[="�(�1��<BM��>u1=�1-=�<=x��;�34=X��<9vE=�
����\=�8'=��#����<�K=�K�A�c�m�e<[��;�ݢ��<0�Q����;�Yx=��E=�s��D:�\I{<�I=�?��G��:�Jo�ф�c=��=&��<�f��[�<��=��μ��=�HP=�la���:yт=D �<MJ���x�<7=R�:w�ռQ�<�L=t������<�?O���u���<��¼�@����<�a=���
���Aj1:1O�;X5뼲�!=m�o��� ���
=��U���}<���;B^u��r����x��:2E#<[��;[Q�<ӫ�<?���l���W༽�ܼK$b<6$4���Ƽ�*�lXG=Y���� =<�¼P� =��<�4���<G��c����P��b�<trS=�jN��N�;7�\w����=��(�����q�<��S�t�=�� �
u�<ښ=���#�$�)�<%���<E�=��� �=ڻD=�8r=��`�/bI=
�;�3�F�<WH�<��'=O_�;x���)r=$8=�=�X�<!��><���A�6=�:��w0�%�T��[�;aB��ǼA��s�;Y&�;�����=K�J<KM�;_�I��y�A.���=��d;���<S�Ѻ�G �)�?=�~�<�i�8=�S�6��<��M��)=�
 ��9v��Q����<[<`�j9�<��4=_KN�(��Ǵ
�@�;=�GI�jWf=��<:1=�|�<˲+�ʋ��u%<�0��;L�@=9ܛ<T|��|'����<�>����V�q��<��I=���P�:����� 5��'U='p&=�,.��(=j\O���V=Y0:�l'0=4��"kX=�E�TL2��c�<�\�<�����F=����e�|�c�*3G�u��~\2��AҼ� ,�{�9<d�ռ}6=EH�� J ;��	>����N���&=�8���Q=ɮ��NP�%]G���^��A�<�\Q=	X�:@��;��=jW;�r)�L�w<"�	<F�d���R���"=����?���];��N=�M_�*9��Gr=�ԯ�1\,�?�)=pL-=KZ��[g���=E�;��;�ۉ�@ƻ�q;�h�<��t=E����?�<��<�Ƀ=�E�OG	<zi=N��<�"Ҽx�<��4�^���Q�;��׼�A<�%=�b����D�
<%0H=��<�#<O2=�m=��<��V�Ad&�Jъ<�k5<p;�qv	=�~�<� }=16�ҍC������iM=��=��g�'=
���(`=�UZ=��d�Fu��ڄp�N�<�G;��#���(��1B�\ ]��'$<2!=)ݼ,c¼܈�;1W�:7�f<��=��-��e�<�a��0=��A��p����V�FI��ay�<��A�eQ=�$�;u�鼅��<���:�<J�<6+J=#	��Ғ�7Ń<Kw	�p�=�5<M�#=+?�<n�=~�y���E={�޺cz�r�:��;�=V��<K�<�s߼�mt�o�?=���&��;��k9=[�<(���`��<�SƼ��غ��<��h��%P��`$=5�Ҽ�<�cQ��p�<F#(=�J>�l�ů�<c`��ؤ¼J7�5�<1�v�	
=v�ϼ�ռ��z=�S�<�S�LA�:Q����YA=<߼��;�<b�=�4�<�W�&Qb�5�����<oT=^�J����*I,=�^���;뵰��]�<-�μ������<l=֕�<�8[��;�<qym=�M^������B<=�a�� �<���;C�=�������w=#ݼ;�����>=�u6�6>=���<z��<�=���Iv8l��ѫ
�$��<�x.=sJ����J��+k=/�q�H/?=]�J=�aG�%62�;~L<z���Q=�T(��V:=6nk=�;K7;��L�oP<��s�4=��r;Ԩ�;.ﷻP�F<t9�<n��2
���\=�Rj=��@=��<�/<g>�s��b�E��W����<�@���r={�g�i��:�+�=T�μ���<4N[<x�W�z\�<d=烽?j.:f{ ���=�#<�NN!=�R=����� =��P���K��<��*��!t=���v\��P�j�X�Ո��F(l:	I�=��{�Fr=<�n�<j�Z=אk=�Z�=�.^=�zK=X-����j�9=�2d����<
0=n��;$�l=���T+=�$�,Da=4�޼�M6<N��=�PѼ9�;S���=��="I�<A�=>K]�c����<�*�E�к��
=\�<a���qnI<�Y=��O��<qM]=q��<��B=_k�_�v=F��<�eM<M�K<������<�x������=��<��G�*�����0��bs=�.̼z�a=����iN����@���j��J�;B�*�+��<O��<�U%��Ճ���R=�����;�X�d=j�мZ�U��f���=&�2��,q<cY=g�<�\��+=5
I=�#ù'>B��3�<�뤼��'<���2�=�C)��H6;���k<������=��)��t���=��;#=8�_p�!�+��|9=��D=�{�;��ӼC��<��<��;n_�< �;藐<pܿ���y�l=����{ =:{M��D��pҍ���O=_�#=�I�uV��4'�<>gZ�	B�<";�|/<��,�e�1p�<
iѼ��*�<%�(<�9RrC<G �<܇%=䢉<��t:G�����������X,�h*X=��<Mm�<Ū�9��e���.<:3=�Z#='-=�=:�z;��"�J� �"g{=�k-�JUn<���<D��<�;<�G=��'<$%���1�/<�5��^O��ֆ=��&�,=Z�)�Y=�`��5�;��ԼΑe���u���8���</?���`<�������<��7=ag��Ӣ;�ܻ��F�]���E
,=@͙<k>��=�(h=�׵��Z�=�����|���R»��{:���;��g��$����@=��;�Z-��H%=pH
�-=��t�u�E=�NZ�t�Z=���;aQ������p=]q �����58��8�"=�iB=z	�4�E=��8��10<��2=��K��β��;ۼy{=�=}@л��m2м�{.<]�:��<��<ݾ�C)��SϜ:�i� ��3=�Af;U9S<)"=Z1R�����$��<b=��:���|S
<�	��<A�*;3���qY	�I!�[��H|����=�o�<Z����J�����B���%=��=��N#��0����Z�s��<Q�6��'T��F���8�0Z��nˬ<1uU=���<��=�;\�	=g =<C�<,S=�g�$1ż'�=��x�����4��<vWj��C�<����M=2�;$��9e������8�$=�-����:���<�"�qܟ<�)ҼQ�S=5��٫<n���](� `r��z'��\ֺ�u<p=���w�ux�<W��
u=����b��m�p�,�ƼE� ��ow��$��ࢼ)B0��L!����<��O=�X ;E��.$ ���K���T�7x=e4=���[��3T:�(B���2���<�޻R�ؼ� F��+�;=�$�����=�{��6=΀=á����8���,<�[��ӟ:<K�<�F�;�Z��m�<�1�<7h�T����˻����/�\��bL��v�7�
=�f<xN�<m'�uܮ;�3=��0�ћ��=�����]=t�H;`#=�p޼L=�`<Rh;A���f��6=FD=��-�� k=yW����ڼ<�?-�X T��ǋ;�<��?n<���,P=����/+:=�F=&��<�6&�'��<�=;tm=YF��������e�9C=&=��n<��̼��<���<Y��<u��Tp/= g<�k�=�7=�#���<�u������@2�����S �I�B=��<��o=6<�2��_?C<~�J=sz==�=�<��s=�=7����ļ?[R��{^=z͉:�;V<zԇ</���r?f����eѼܹ8=i����g<d�@�v�=�:=�3E�������H���v���{�0�<1�==��;�x9�P�<J]���=��==�6J=�ݟ�Q��˼&�S=z�T�KSS�i=��k�@4k<���;�Y�dм�̹<.x���(<S:���d
���-�Nڼ?�g�!�p=����=� ����^��s:<i�X���N��rZ=R���y�=<*R=�|˼:.�;=�ͼ�%9=��>��!X=�ϼ<�I=%\�rD=��d=W�9�����JA���Ƽ�!�< ��<���q�<6Y	�,3������ς*�x"=�ZE=�
==N��:e5�'�D;+� =vM���q�<W�;qt��^0=)��<l2U=o�3��wo=�����W<��=��UR���<�(=
ݻV4��[/��r����\0��
J=��<���<נ��VP;��!=&�N�z�p���C�:]�=�|:�L&@�#O�A�<���qC<���Ar�����˗����_��C��X�<;�U=�Y����X��:Tm0��ŉ��o�<?����L=�x��$�<�	=�ʂ< �$=�P<ݐ�<;(�@^��"`<����r-@<�d"=���;<O!<ʣ
��a$< Pּ}���*Γ�`j3=~�����!�@�ļN!�<R3<�\=��=�~�<��O=LI
=*}��	�
����A?���<�b=��9�x:�M�	=�:D=��<�(%=«=�w(�ɮ5�� .<S<,�<溞>Q����<�0�=�����<n� ��#8=�vR=���fe����=l�R�f�<d x��N���==�qo=�������+=�);������+=V1`���;=��[=�i����<�;_�5=���F�4aC�l1��⧀;����&�d��<{_n�� Ǽ���=�%=|���	��AJ<sl=-�V=:�N=*�T5���D��;F=2c�=�	<�3�	��<L�$�z4ջQ9�<����^ռ�%=��R�Q-=��򝋼Xc=X1�<2t;eBB=){<3��9=s�J=
d�E���2�N=%��<�s=�T�X̧<@���c�;�F2=II���Պ<�N�c�ݼrd&����;�w�;���;���;w�/=��]� ��<xum��O��;��B�<��`�L=�G�)p	=\��;��6��*��ʐ<+dP�ѽ��ȼ�t�<ޏ
� �;�b�Q<��S=�ٰ<��5���ͼ2��<.����@<��Ƽ�<�<!�C�]��;�q�:YN=&��<���;I1�<���К�<���2�=��A=q�^=>A�<}"3��\�<�m���]��>=;g��*ȼ��ia_��"A<�q$<��2=G��<^�y�&9�ۭ���?h��V<d<wW�<
:ػ��;<nx=\�>�~��(( ��Jܼ@�?=ҁ��uA<�@�9=ǝ"<k6`=���<���;���<LAƼ�#��׼��ϼ�$k�$^<��C��H*���<�-)���4��`�<�b=~O�=�4F��Ph<hGj<lMo���P��T���]=�D6='�<���=LQ�;�m�<_Bм�=�'�����WN=�6=u�(��"=�t���9<@=+�H=�o�<[e=�$	<�i�<h6�<s�-=u�9=��	�ݠ&=�g����<�M�4�ݒܼ�4�<6�@=h@=�΄�V6=����O�#��h=awϻ �r=�-���w޼V�<q�H<���˲�c�[=mf=��w�ע����=)4=��z=:`�b��]�C=@�N=�j=SR�<k��%W]=��;N�=8�l=+�����(=:�MPS�ғ�4r =Xwм�	��������<�;�ו<ї`=뭼<v4�߽�1˴<�~<	�<7�<��6���<h��:�	=�c=u@X�YT�;�����o�<]�J=��0=��Q�y�d=_j=ݿ=� ~� ���e� ��=��<t�q�a�H=b��<ٵ]=IfE=;=��4�<�C=2�{=ů=.uV��+a�=WL=q�=��V=�	m=-��<��H=�{$<j��<� �<�e��R�;��r<�~�<m0���T=+��h<�<� ��E4=h��;i�A�&s=�R==/
�x��P&'=�����B�<����>���$���<�Լ!�D��2�<t��W�������d��AW=Xt_��0ؼr۵�n��<�=Y�>;L���c�<&4=3`=x��q`�F=��=o�<��=+���M_=�D=8�j<<P�<aED=dQ��D^��1'ۼ��M��l�<Q��<ӚP��n��%X=�[f=�r=@�;H�����B=�Ά=��1��	)=���<��2��6��\=崠�}w<��7���<��U�34ռ�����W�c�	�+=�<��=4���&���H�<)|"�����a����<���n�O=�5<�C�<2�<�*�<s�^���<��<�O�J���NW�Г>=^N�<+M�ԉ�<Ѡ$��IK��s=0�=\�;�y�#=���a�V=tS�S8�×�<����������Z^�_tC<�����Q���޼�{��^uؼ�D=���-W�A�*=2r�|q<�b��Io�zH<��_�����[=��K=(���.y�E��40��U��X%=�%=���<o>��0Z�<�����F=E;�<��<;�;2�#��S�<-]'=�C���3=��;�h�<j7`;%g?= ü��l��4�<Eϼ������Nt���2B=4�ּq����H3���=���if�<mQ�]=u�<��t��c��B';L�8����=�*N=~ 伓"�<��I=R���� �<&m���ݼ�
������
2���;v;g�R^3�.i:�������i�:�<�<��%<���~1=�9%=o$=�����#{<ܹ&<�{%;cp;=*Y�:J�a=��s��>�
�ck����=�qͼ��Z��~-=��<M�E=��<��	=�}w<�b�=����|�ؼ�o=��=��y��^L=��W��Ξ�o|�<��;�9=�߼G/���(�EE���vLb=�0���O=A|���=x=$�gR�<���� �:;yI��Am��L=QsF=}�1=�6���6=�5=�1k���E���:�?"=Dz����ش���A�<ƃ�<�-� �<6y���K��ڤ;Ὁ�*���μh�ּ����Ԇ�Ays=�N=Zm��8;�Ѽ�<�;��=P�B=�o%=+^=�ο��A7��2���I����eo�Xa��?��Q1G=s�;�<�<���<��ݻ C\�7}����:�V�������=�=���)=���<��d�WE��}Lv;|K5=u7��W���<=1�<����m?=|�=~�9�Ok'��6�;��g�K6�<}���ѢE�03=pM��|Z<�"�8�����@<����h�Ȼ��;�#<%у��q���Έ�2�:����57�<F��<�ݧ�˶J����]iջ��<f�n<�9
=g�=��	=�6>�rnT�%�s��>#��š�v<C=XB��0=��<��Ｖ�:�F�J=!߻MYD�T4%�Ĺ2<S�Z=�E�=��N�^Qj=�2c�,v(�$-=�:�<�(:�O ��F(�:`��]B��������<��b=��a�����a��;�գ<�l���3���{	=x�?=7���_<��NiU=�gh=���&�;���A׼Ek�;���=ᐼ� �봻;7�7=*0=�g��Z���u��xJ���%�}�d=c@{:d�[;���<����*<q��Ar"�(7��lr�ڼ.C=d�=[���n��S����=Yya����</�����Y<d���C?�2�;��M�w����N�<jM��B?;�я<K�<
�%�u=JB�<��<6ϼj��<��ټ	0m�^\=����"�;�_��?1=��d=g�=�U�1,=��T<�3���#���%���<Q�;�	��6;H;�<��=bV̻־�}̼�YL=N������(�]vj�70d��@7��<&��]=v!�<�+��b�m=|�K=B��<0U=a�Y�(��<��	��}�@�B�%��"�Η/<�d*�������z�0�Z<@�]=�=�����Xt�{4@={����<�<�W=�8>=-	�O�>=P^o����	1e�a�g�(~�;X�!=������{���q`u=�)=:db��q��|��y=��<�R<7-<8�	����:|.�
=i�&���;`�}�F��<���<(�s=�-����D�% 
�LAϼ�=���<O.�4c�<:2a=V^<��?K� �;��{=6�&�s=�h�߯ =���<r�S�7H=�.�<%�%���$�'?�:]�<.9=�+,=v�w<������;���pf�<��<��r1=��=�$=��L=��j����m�<l $�9��r�U�L!"�ЕU��v9=G.V�2]v==}�:���;�ܼ:��]�&���)��;�<f����3<ϳ	�����t��W<g��<�6A��=�ؼѺr�֛R=$V`�u=w���<�gx�\3=�n�;�A!��=���<�B���@=����<"U5=� =�6�~#A=� �mb!�D�R;��V=u�a=�C=���=z[p��V���;<�{(=��5=��<�r|="�޼&&��ۃ=�p=�4	=���<�}#=|�"���J;��<<�*M=��;7݁=��� �<)˼{����?=c@=%;�1�.��Lx=#?=z�<�*�<Q~��뿺���/��f=�;:C=cVc������1=[�<pN=b*��Cx3<���05��O���;�!��DI�fR=J�O=�r���k;�i��I =���<>�C���Z��2��v�`�k�:�h=��<��<�&=�w���nP�ً(=>�=Z=@�J��jX={���#$���[d��_��N��Q˓�I]�����0=�gl==Ne�<��`��<�H�\fżaz�=gx�Ű@;,�6=5��<�0�#[<h�;k�j�UTۼ��]=2�H<+�n�
�V�)=_�W=�$|<��P�?�=�PԼ�E=��h�1��8�t���==�6�=��M=+���ԍ;�o������bL=>O���!5=��Z<��<��<�Y�<_c�!?��g=��<U���oE=#�� ̽<�x�<����Yw�<s�L�F?���
<(v��|�	=����kܡ���=i�f=���;�-�<hޚ�q51=0/ ;�м�!=N�_<S�7;�Ӊ=T~�(ڐ��>:*�_=� �<,C=t��<̆���r�h1=㖎��;qI��H�<�Nh�m��13�<��7<~��<Aa=~�4D���<dR��o��+Oy���=�o��x�+����;�k^=��<o׶�{&�:��3;z0��IQ=R�=g��n�U�T�F=��Ǽ��жb=�����5�����<��ɻ��d="�<=�k��3;' �<[�<���`�M�1�@�_ۼI�;�?�����y绚�(=='P+=A�[� 9=�A��|0<ѨI�5�<k�>=�`;�m���)�t�üfH����*=G�弞 =ɟ=�u��{9u��<��3<���~v���=;���;��C��<��ԧ�<�^\=��==���<��~<w����|�`61�>V���<�_
���Q=�=��=��A�����M<�{��K=ʡ��赑=:P�;8/�<��0={9��ǖ��=7�=�7)��@3�K_�ȩ:���<�ԋ�ח�<ĉ��%=7�=�-��?s��4�<�_C=X��<Cs���#���<[��@5��ہ|<�=�,=�;:�V� �<q<I�;=�8W=\W;<��x<1p�JX�<`,�Zum=c�=�?�;�]�;<#ػ��g=�=�<Wd���=䵱�&n�<3{<����c���:��>�<��ܼ[�k�~�<`����XL
�ֵ4=g+�<��.;�%=��/;{E(=�:=��#<��g)�<��s�KiżmR�<[%,�q�<�i����<�X=d=��)Lj=w��<��=L®�C-+����vZ�!C9%9�<ml�����`���u= �ռ�^>=ZJc=���=�j5���r=7 7���<��伍ǅ��&��-��V<�w� w<��R��}�;�n��#���5��<s��I�6=�%S<�Ƶ��a�<��<�Ă=���<>[D�\������/;"�:=�F���&��G0���<�<�>[�����c����#==-����)�PqD��/,���tm,<��
<���<WJ� ʎ�+��<�?ʼ���1��:]�c�Z�9<��=� ���׻޼�Z���[�<�f�p�+=���;�$6�f�8�}7�<�B2=�<_=��V+�;;��2<�\d�]LͼG=�1���<U� ={0^;���<�A=�XN��"����܏.=�]��S�48N��=�=�{�<�}�;9�D�]'����<����Q=/KS=Em.��A���8��Ao<�<�S��;>=V��<iɮ�\�=�������y�
��X(=��'�%��>�<)�<��Hx�:���+��<�d_;ڽ|��+�[�3<!�ۼt�m�K �+=忂���=gܼSUM�+=Lxm�o>��Jn4<��H�l�<R�<��	��y<o60���%�%��m5�<.�Ƽ�)!���F�0J=H��;�Wڼ��B=rC�������N=���< �<m��;�S/��bC�^j[:KL6<.of��sE�?å;�S=���;1H"�����`\0�R�]��Q�@��;�� �s�%<A�Y<��<ו_;Wr=�i���:�"�*=.�<=���=W����뻾@>=m3 ;6�%��mż�GU<%sK�o��<�r<R H��xּ�.6��%<]��<`�<�n����-= Tx;�i�<�=�h������6��q��<.�I=1�|<X�/�M���iQ[=�걼�����mo�}�G=ׁ�<&D��O�m�0_���3��s�kr=C�~�)�X�Y5�<�aʻ��y
���J�^<��b<�d3�|&�T<��%=�lf=�߶���/��'?�sg��l�<�;I=7Y�3�ƙ=��	=Β�=�c�~�<N*�:��W�F<Xa�<����a���=�?��=J	X<�;����9F�;��=��<�_����;��I�~�F���K<�A��"?=r��<t#���<��$=��+<�B�S�м�:2��
p=q�y=�w2=��Y�i��<_t�<UM=��=d�<4F3=VW�<�Z%=�JE==R�TY��c�.<��B=*��A1�<�g���'=g�J��h��`�^=o��<˷�<��B=�sݼbmD��ü�_3����3@ϼ�0��j8=3�ļ�3�%�b<��V�8�A=�^[=ʅ8=�<!]l=|(@��ެ�(y<&<��P�ҹ4��F|�����w5=�� =`ь<��?����<_�˺������<��-ㇼat��&�<��<�ח��F�]g����2=+�!=�3�;$4.�-1�?�<��'=����VG<��K=��<Qp���=����>�$��8�<���<l��<��I<|i~��|�c<<=��;�g}�XT=�O�;�
O=0��y�����;hJh=g���9�����f<��ѻ�X�<��`�^�8=�J1�wx<�Ƚ<��<�<����7���=79�T��<��W�G��T�]sw=?y<�H�<�`J�� =f�/<�盼��z�����)w<db^�d�5�*~i=�U=��h=�Yb�,ᶼ��1�N䣹F8�:�VR�8�˼��Z=K�<l��<��<H�<kH���!��U;����.=�p�:�H=}fƻH�=��;�p~T��[���<=;�&�M��� <!"�<�5���D��%<K�<�^�<���z(�;3?���_�u����<HPf�u+<wػ<�X��ԉd=����&D���Y<Z�<{���4�	�<��0;_f��u�˼����R��)�9=^��ќ�</>:=Kk7��o�<3LQ�u�`��,=3 ����w���9HK�c��<F{�:)xb=�=Zyz�V>=����<���
޽<m'�<�<c�:�6�:V�(=-5#<@QF���W=����f0����K��ѥ���9=�_-9L��9�*�;�&f=�M���Y=(A��$��<�`;�2=p�=��NX��j =i�%<L\㼘�<*E�;��$=0�V�Pe�?��<x&�<�ټ�X=<�n�;2�`=�d=�<��9���8�?�<��?;�'Z�U9�`�<�@�L��g�� ����\���<�"@��~u<����H=�_h<���=��6�[d�;�f={�#���T�?��<��<
��Q�R�߇��w�9��+�U,=�u=�s�<��91�����$��|��b
�9S9=+��;�7n�0o�<+ؑ��3D���7=<;�<l�;t�=r=��=��'<^���!W=���<�=���<W�E��Vκ�����!a@�Kp�=y��9��\��뛼`�	�^vL=b3-=!R���=�'=Pw��q�%��!��\�<ju�Xr;<2����Ҽ�B���b�G:rO�<bAk��4�d�<c�H;5���n'D�ƂD��K���b���q��0��LM�"�9�3	=I�	�_D=*��;nt=;�l�Wf�'��<�S�ü���9�;��
=�	���a=��!=����S髺�w���_�&�t;���:H�=`�;�M�;rN�%8���M�c�.=բ(=b9=�@�;�̬��^�*=�Xܼ��<����fL����[;�YἋ��<�g����:P�<���;I�+�mr�<�| ���Y=n0�<c=�1G=��9<��ϻ�m5�����z\7�}&���L=Uhv<�1=�(\<��	��_A=�-���;���<:��IN=߼�����<�vY����<B�#=��^<��0���뺊����o<�S_=��p���;�C�<
#=�B�<L���M6=k�#�^��<=�뽼��<ރ=�W�<��8�^��<T�=ή#<�=	<U��<V�;=��<#���Oy�(�N��R��Q=��O<�86���;O��9��;ı.�Rv?=�s�62="�;H���Ҽ9l6=��M�1�a#.=�|X:C0>�Wv:���=Q�W<���<T|"�}̣�}4��v����<�pq�Ǿ0���)��q��"-=:��=�Ӂ�$��<�^߼��=��c���S<��<Q�)=.���,f���C;� g	���[����<<=�=]\+��z2= �!�'��<��L��̠��F=' J��×:(W��=�<����wT=���<��<+�r=��b���4�d1�E&�<:���:�m����y�+��r]�qg�<Zt���C��I�gjH=��<��t6=(�N�O7=�~!=<J�T��=<偽�'�<�B������F=�;=>��
�ұM��?8=� �=�%i;���j=B<��X�%�	��F6�ei�;�����A=���=4P_�i3��Lʗ<,]�4��h�=2м䖵���S���=f�C=�?���xv��E�z/5=���48����=F��<)��;�q�<��R�ڎ <�(�3�Q=s+ӻ��a�I�U�X�>=>����o:�=�z�8���2�&�[��X<Om�P�%=pbV=ͼ�;"��<��L=zR<��n�?����8���|�65��y���i��;)�9����]X<�j=�A=(���y7>�QF�<�Q=L@����I��!#=!P�<�Z�<�xW<�\�3�<�j5��l� �X�1u?=�^�<�HH�D�����
<a�v�z=ZD�9�$����[=�}���<�:��<Y�0�m��<��=0<O������W=U���}t�.9�I�<��A=p{D��u �%2�<X�=Z\�tt�<X�J=��<�[���l���ׁ<'=��e��T�:_Y�<��e��W=�l������<��\=����<����<Ԏ{���=��D�Ӹ=N��;��<}h'=�j
��ZU�Jq���~0��M��s���A�^=m~&=�=�à<}�?��y=�&Y��
=}���I�t������[�e᰼�*�-3�|�<��� �E�2���[���5��Ż�� ���x�A�I�n9���<v.#<����"�B	�[Z= ��1���+�]��<
�-=U��<d���*F<��� �r�;X��]�=_D=训�� ���k���L�<�û\�7�ԋ"=�Q=��u�S��J41=��;ȁ�<m���N����*m��uV=��w���6�Ƅ�P0<��J=gm5=�gռ]�i�rW�:4�T:B^�;ew��s=ʶ�<8�<!3=$M=$���\����(���<�5=��V�kL����;��;}bߺ"�\UF:�=<<$?�ڮ��+*=KVZ�Ȱ��Ӆ5�/�<�)��;�=Og�=�� ��;33$<F+7=�v�<dND=��\<��輗x'=����'���=�����;���P`��5=��"�yC�:?B=)5"=f\:M,6=0O�<a�L=-<�����<p�<ʛ�<Wp���+�\�N���o=P����1=�;�<���: xy<!lw��t��Ȼ��3=u�=���,�z<�)=�(��-(�� <	<Uw��:F�ah�<!6���"4
�1|=�g=�z=��3<M9=�6:=�UY;��_�G}�<<؅=�FY=1F=��=�o���pQ=.�=���w�7��<V��ڂ�;|ϒ<[R�hc�;q�Y����<O�[��<18����������,�9����'=ɔ]�3�P=Ǖ�ّ==�����D���c=�==�Y,:�����,�����:<<>;�eg=L��
⼕ϭ<|C_=~� <�������޼��s�������6N\=���bdp<�>����ϼ
�a<�Ց��!���Q=���Ӷ�|��;�#P=�θ��-�<��K= �c�%Ҽh�-=�i�4�=�9��߫Z=�< a�:×��<�mY=�N��Ӡ<��;:�U��8=��`��E'���=-�$=Jc��y�U6�P���<;���1��ME�� �O��-1\=#=2?T=9�����Ka=H�=:�¼:o,=�%�<��:�JN=f-�r廚����xڼ��B	=$��<��ຮ;5=�P]���k<_�|����<��3<� ��N7��&F�	Zo��uQ��ʅ�=�*=�ll=q��<D�2=o���$=,�&���F=��Ҽ��ɼ��/��� ���м�O&=ڱ{=��t�9��=�A���m���ļ������si�/�ۼ��X����;��9�x)=� /�(�;�!=���B�:�dE��z<�c�����N�ͼ���mh���I���,��Ӈ;s�M=*7��z�U=uF=�;Ǽ�D
:�;���<C�g<��L=ƅ�>+<ۨd=+#H=��:w���c�\f=�D�<�.�=o�=��#=�=�f:�x<Oq1=����;�߷<��D<R�3���M=��F�V����=#=�?N�r�J<�="����g��+8H�
c�.ʼ�&�<{�N��z�;�;ټB�s�<%\ټ�J�<����E7	���<C �<Ic!=�QO=��;�LeQ�x�<k*=Y��,Sv<$�5���i-ܼȳ�=�'=�:Ӽ-6=$u;<�i��$��7��J�����T����diȼ�J�;���<&�B�����	=�e;��T�h�=>m�T�,=s_���%=�K=�2=(�=���B�$���P��z��
U�7G�<2�;���<:���L>���'=�p�<=
R�o�=h[�<��&=��+�_9{²<�d=�{�����/=�k<���<�ϼ����
=^~�t4!��<�;U��<��?<�;e��,w�}<9YW�,�_=��`=��]<�N�<��K=�]��w�<��z<��5��>���9�ѹҼդϼɕ=ʹ�=9�ɫn=W��=��b������z<��=A����%�;h� �����i��2;=���<sk^�6�8�y����;�#�Vd��b��1�Q�4-���2��T�<=�;$vB�+�"�fb��Q�<Y��r��<����B�!�� ��"~	�eJ�*�4�����"����B=�ީ�s�<�l���#k���ּ���<�+=U�=CӺ���;NA�;��J:�r��w�;�4D=g�{=/G�M�2�Cۭ��5��<E����<�v�Lx�;E�T�{�:=��ܺ���?��4�v^��9I��R6=*�L=��_<S_��w�=� �;��\�<ˠ;��p=�bƼ�)=�u<���< 
=�uK��'@=X�&���c���b=v�U=�rK���=l��<�u<��!=�l���R@=�����r<O�G�̬=:j��2?=�2�������"��Y8����+�=S��;�1�<�Q�f�0��*==إ��8!�E=Sc=�H=H�#<�q�<��2�t*��&!<a簼A��<��<ADv<mם��"n=Ê�<�F�<r0A=�v0<�u)=��oJ�:г!<YE=��K���S=�����
;�fG�b:��(ۼ���f`3��=��4q�<ߓ��Ƞ<0�<��2=�S<��o����<����@/��X19ޱ���';����1�h�E����p=3�2<s�<���<�����﷼$�#=Z=�����<&�-���꼵�*��񤼻�I<_K����Y<���Y=R�=���n\�>F=��=�`����輒�*��W]��٠<��<�+��%�<��<�=����v԰<�����@=�H����A�*���8<ia����*��0ݼ�gV��JL��:=�:Q�����N�;�|7��)��O�v<
@)=�y<vT;��B=������	��I�<��z=-�,<�b<�q3<��μ��鼯��<�Q�;'| =��_<�WX=`)==��^�H���#?I���Q=���;^t����=>1=r�>;�����=b\y;�u4=��=�1��64�<֝�<��b�Jƥ����FX���;��P��󼡬��J<��%�s�ź�z<��ܻh-��麼�=�Ҵ<�|&=v��<�;V=�Ge��j
�:�+<�T���=�%����=\x���H< �{��Q��c.J������ o<�y�<�8�<�^���O<<�A�#�m�}!j�k�=D�_�;�KY�bg_��E�<�U<2���<��-=!�u=@X�j�"���`<��f�R6��ic,=W��@/=튼M��;9�?<x�O�txP=M�>�g;=�n=��:;.OP��+������T�c=-	��{��5�\<PL�=�	=�u���,<z�i�o̼n�'�rT<Wo*�X�h�&fQ�j�����-��=��=��[Ǽ�ً������I�]ZA��u�<����E�SOҼ1�?=�;����c=��`���!�O�<�bؼ������<oZ��xͻҎJ�y��6�(�'���e�H�s=�M6��v�;�ߦ<��j���U�t<�AY=fŉ�f~ =\��<T�<�H�n��=׌< I&���<��<���]Ѽw"��E�+=��Ƽ�7�<dv��[�Լ�;W����<MA:2
!<c۶�_Z<�1=��|<T�Ļ�����=�w\�F��<�<z)�De=�5
�2�=ǽ=�y����y��;^�p=�8��}*�������4��OV0���<#�H<�h<�R=�,9�^S������;j]����7����u=!�H�΍��.��i}=�7(=; �j;�<a�����R����<:�:�G:��漝�����.�; �/�<4h��=�̼�@�e�� ��"ww��LK�t�I<l �Cx����4;p@<�'=�N<�Cͼ�����<S����^_=�8�c-���p=(g=S�(� q<N�C;�+�<�p����G<��Լp5;��/��<��<c�;�w�<%1K=M��<-qn=ߩ4���ۼ������;<�<7�j��	��R�+���뼼b����\�r*��w�3߼���<�]��*ջ����s�P ���|��pӼ!=��<U�g�߻�Լ�� �<�Ʃ;���"�=�*T�0�����v�#����	�,Bż �^�/<{Ǽ��<a=�;ʿ7<.d3�U��0_�<�1e���L=b�<�~^;�g�<~� =�a���<�<��<e����>=�M�0����hq��u�<\�Ҽ�8'=��=�Ȫ<�6V=�B�;�c<��<�|l�oJ�;�B�=o���\���|4��|K�p���A���<�U��D�=��7=��~=~==�=8b�,��<�f��:1�|�#�8�<�H"�H�<L�I=;�<��9���C<�#��<W�5�9�Xp�;&���ܜ���C�=G=�`a�aҼH'E=jA#�q��;��<����� ���<F��;u:�<~�ϼ2Wһ��=^/=M�=	)3��%�׽=�i#����<|&�*���ٖ����*��9N�p;h�H=ʏ���9=�<e=QM;$X=N��}Ze�^ 0��'[�E4<�/�<�O,�LJ=�,���V5<�G�<OB7�nʖ�!2=��1�6g����/=`���?"2��W�'A��<;�<�"���c=7�<��A���!=JbּŁd=L[V=س���7.�IWe�z>����=�)�eU<]���u�G���s�� ˼�w^��Y<��Yꂼ�;�<�-)=�;=ޭ�y=5Xn����<==�K���W<{jg�}���Dɼ�F����<��,<�ӑ<q�+��a��%]�0{8=�4>�)K =�٪�;�f���<Yg	=-
��e��Ș&<��3�Eu�<�����߼��ǻ�d=��;��C�p�ۼw@p��<�;�����(Ļߖ�;��Y=��0��DP=S�}���\=fa={TX=����S<�.I=��<xsl;K��&p<�M=�:��'=�����=���<���ϼ(�=!�u��c:����<������,<d�"�Kt�;�h�;�^R=�����y=9�6�Ĉj<u��<�{����<p��i-=��<��6<݇�Xe�pp�ON�<��Y��2n<��n=q�D=�Һ�B�а�=��D��K;gn�<0eL='�T��b�T�V=��<���/d��2=���<��^�-��;	�<�a����{l� ��<�A��L=�<�29<�n&���o=�+=�L���ͼ>�+���R=�������b�E_Լ�2�<7��<��T=G�:��}b�<xZ����<F�;EA|���=�
��T���b�H=>�V��<H�j<��D�7��s�<�zM=B=)��:Sx=*XW<-v�o��;}nH=`H5��3=7�2�=Q�P�W�G�|���D�8=ҽt=kS5<�;o�=Yݗ<��F�q�0����z:=��=�g<9=	W�_�h�)�}=� �XD�<X��<�R�;_a<��L�lڰ<�:|=r	���|9�2Ժ������<���;=�[M=u�=]��"�̀y�h7=$7=��x=g��<��}���+�=uWƼ��L�,0��"�j�N=l�S�І=m�<�k.�.漐e�;���#�|���F=��(�;�)=s��<=�L?=M ��s�_d	�-11��=`AG��z���<��|H��μ��;��<k�w���=8c�<g�����L��h<<	�m䥺*d��K弨}e����<�d<�G;=C=��&=J�<�Y;�͑�:U�=�&�b�M�q��<N�<�fܼ�_<k#�p� ��PT=V�=.�Z�MM�eW=�J =
�o=�6#���=����
Լ]�P�j�<1�;��Ff=<N��F�l=ȝx=����r-��P=Y�H=b!<C��=��P��;�=�F�r11=>7�i'�>4*�t/Z<��<�bH:\�=6x>=|Up<T�+=��<$\<�o���1�����"|:�S���p]-='��S�<���<(���6�<����Zd�X�</�P= �/���/�&�<u�1�M|�)}�hx/�M��<&����;�O�=���<u�<�8�.��<����j��b3���o��@�M :�B�6���3=NJ@=	E�<Є���=���� ��=m�H�@�ù�}u=<]<_`��Q���e��L8��M��b�<'ľ;"�W=���;��r;eo�<����L��d���*�,�M=�.�<�d�wȽ<���������<L�<<��=�J�gݲ;#�<# ����l��[�!�.��<^&�<��>=n�W�hc�;{;H=�U༎�Ƽ9XżL���=&Ed=$�V�W�G����Gڼ�a==tȀ<�=Iz���9<9w�;Y�;y��<�H�<�7��@�6=�Na=n	��Ȋu<������nyk=�¦���n���	���ܼN�=C=��8��䊽]�<�;�$=�񡼄W�<���<ne��2׼��U�2<�c�1|=�=QB}�ti¼�==AO�<�{�<��<��!�`�/�z���=e�<�Sɼr96��=�U==/=�@=nČ<,��<;�<>�z�5���1��޼,:g��X�?� ���<(|~=M�<U=�T=�q];b�=��8:� P��e�<l�mޭ<&�9<�
 =2����*<��
=���<d�t�eI��D���;�X-�7��Q�t=WM��"K�bZ�LN�<��=W���W=��.�|��;[�ûV}?;�<��ug<Uj=�V�0I���b^�_�P�n��hW��b<�y'<��ݼ�X�k���*����c����� L�<a�K���:��<��T�2d���<�(��،���~��C=Wt�<���������=�Y�hsv<9 J=
C�;�+����< F=�{���<�_Q=��<i�ѼO	Z��W�<j:N���:=�7�=4#>=��a�;:�� dͼ�����D���D��b<	ܝ<�"~�3=�;�i0��J=&���|=��<�z:n�;���N��l\=#-��xw=	�W<�,h�N�R�jaJ;�@߼�ϋ���;Rnx�m 
=qۼ�5^���#=Y?#=��6=�	�<�O��#=d������X�^W\=g5_��:/kD���N���<X�T�M����ۻ�1s�����o +���9;i��Y�	����=�L�;��>���?=a��}.=�9f��|<�=G�=U6R=e;= �F�!G�<�~��e;y�;�b+V= �W���-��6=D��f�=}ʏ;���<J�?����- c��8=K���Ƃ
=.s}=��2��ir���<�����<�¼�:)�!���d�<�OW<aG⼤�P=�Ѽ4)�<�/=L�Ѻ�=~�<]�<H���L��.��%Z=�y�	�<���'|K��N�<�����"�)��<'�/�G�<2%2=@eY��߸<�.=����j�ɲ{<K�Y�]��<��\��H=h3=%��ᢼ���=��K=R�˱�Ȥ&�L�$=C��<8�=��0=e�[=h��<�˼�
�-� �(�d=ɮ�<���HE<�s= ۻ�i!��P1�F=z#K�p��;8&G���<aݼB�]���x�W�,�Wi=�;
=Y�6=ǿ�;C��<'3,=��\�]�=_�u:�I���i��i��'�����@��qm��^�Q��ݼFMC=i�;="� =��A�%2�<({
�=J9���x�=#�?���D�$��<`.<J�E<!Rǻ}_�����g�<�Ӈ<�&�<���; Q�<^؂=�v<)��5Ru���Q�7<��>������@<
����5;4沼v�N�ri@=��9�뼉�"<��;��5�y;�<OA=�r��F��>�e
=�d=�dy��	=o�s=��>�������3��h?��T�F�{<sϸ;��<�ư����m|�=Ne�Z�<V:9=���<{�(=^R=�	�AB����<ͱ����<��<<7=o��; �?>��/�C�TQ��Ӧ:o��;qc���<�0=d�=�r_<O�ջ�6h=o۠;�,��E!�:�_�<�?��Ͻ��Av��њ<��[��L��7�a�<�/���h�<M���Yj=��]�����{��֑�:#���A��J���n?���='K<����3=7&�������{���H;�f�*ں��=v�/=K�S��uC=��#=�y=��<A��	��D���=�&=����]��w�0��O$��r�;��&��"M=&gN=z�k�� M��ۛ<bX�<u[$<y|;=��N�<��=yo��X=!�:� �<������ 9缽$���<��Y=����<կ�뙼�ֺ���7��*�;���:k�<��4����m�7Q
�D�:=�X�< ��;/B�<�麙����U;�o;:?�<b����\żV�k�W�;y�a=WR���o�;k����6��$����)=u�;i���(<kF�<� <�c=B��;d$�<�C��!�=�6=· =�h뺽a��=�<y�?=�d�;j��dD�8�W�cd=�f�����'�;��;�&;�꡼�OY=jT�Z;=���<͓t<������ƻ~˳;	U=��"��\ʼV��<��S�=^x��G�yRs��y�X1��f�<((�t��CP�w���-�<��7�3������<|�7����<V.=4�Q�v�d�-����Ѽ�X�=�����ߺ<�no��7�<(����f�q��ڎ>��U<��6��\�<�8�9������<���<�:d<K�P=7��,p�<?=oOV��$��\��~�<��㼧i4<��S��N=6��:�b\�	�<bI%=:'=۠G�,��	�R��Ǽ�T��PM��ŉ�<<9=]`�#��<:mF�W�Q���=�(;
J�uH���$𼓔L=+�U=C=�H�����W6=8��;�6=B�!��t�<�����~<uHs<}n=:=����iU�Vo;fb�x&<B=�B=O�5;�=�������`�)=v��#���f\�7����(��M=� <��K�0�f�(Kt=-o,<u��ي.�$�b�譁��gn=�12�(��=f��]I�<�d�<��ӻ�u=�II��i����W=�U��8�<�L$=ۨ�;�ve<��;;EWϼ��L�=u�u���T�<���'�M=C�L=���<�̼d��<劌�w�=�,�<zBN=kkG=�%=��<�����;� �Q=u}=j�Z:�o2��$!�[$�=<=��=<Ee=v���R?ɼo�B���=�H=�	����;� <F���*X�g�a=غ�;�:�<EuX=(9=�]7=�D'=�';
qT=/)=���<i阻\���
t=ǟ.=5��:�� �s��U��<��9�|�f������]����<��=��W����>Lo�#.��dna��c��$ӻ�s<�|��򖽲<���õ�����<2�,=,;�<�$�<�S�;�k?���� ��<�B�<�ܼ��;�R<�B)= �w=ե:���<!d=	^��ុ�A�=n%0<�dw���;��Q<��=�@�[��<ǧ�0D�5G=�-��҇�<�f=�[i<��,�<u�����F�n�#�	=�;A�-��.�'�a:��<��tm߼��B=,��<��S�<�=���;.,_=T!�:�BI=��`=J=�G�;�=���+1<��,��c��c���@[%��b�{,
=���<��=t-:���=�2l=��S=���<��	=�6�<e��<������#�����Hc�;@��<���^�R=�S���7�<��'EN=u(=�_�;�5ɼ�1�t�<q����V
���]��)�;=�T=�ᅼ��l=�:'=��7����6�<ԝƼwm8�����Y��M��@G�V��<�Qf<��=f��~�<	�<��a�������+:�+=j�=/�9<۾"��Ԫ;���<S_��ų<4
I����<�L��t���]�����Qc"�h�c=�(< ����C=T]�<�|�<obl=��Y�K��z����x��_=(�1<��M=B�`����� �:he�;��l<�y�����;V7=���a�	=��Z�D:WR����#�-�g=����<%;�C����i<�=A��Є=�b�<�M��� ,�ln<��s<��)=�^ټ�Y�T�+��<h�C�4�=��k��2�Z�m<��<蟑�x*���������<�,%=#�@�d��<ud�#Qa<,�;AeX=��<�⼄�P=_=�xC=/���๼�r��
��*[=}��<�=g6$=.<=�~�@v#��=wҼ6�G=>~
=�d���T�����<��g=Ow�����ɫa<GR���K�,}źC����i�GPi���2=���'�V��.����<���<j]� �(;�m����3#=3�_<v����[����<��=�q���<�*�;�R�U����V#=j�<@{/=C*4�����j=�b}�)�<cܼ�87���a=�����.�9z=��+�����&�=��<]����}u=*4=>z���Z;0�G<=��=�W��ؼ��"��_]�;p:Y��=w�'���Ir�<�<w���4��جh�sm�<+O�;�Ao=ɱ(==sr=�b<rY���.��B=�r!=K�<(���D=D�L���{�_�<FSY=�����ż��_���U<L`&=7�;��=Jr�;g�\<>�[���=�ʠ<���</`?�+������f�=�|���7�~����=kڼ&�輋�a=��ż��O��[���	�<�,��╼�F�3�=d�d=���;~�b=۵$���^��:����~Ƽ��u)=����08����<�Q�o*<DzX<^N�)������ε-<��D=��=;c;���lP����<���;U=��C<I���]x;t�Z�9k�=�C�}J���A���&(���＆E�~?�;��^=+cW;�,�<*�%����<kh��Y(=9��<��=ۨ<�=�$M;Tm���=6�<�I=�4��3X=�(=I���(=0���wP=��;��=��T�`0Ӽ�QN�˿���+:3g���CH=�h���oŻh��@�?���t�"���)�{=�K<�VL���{=h�=ۊe<��l��↼�z?�s��r,���=I_*=N"���<�,l=�E���=h���<h�=�RN	���f���=O��;��r��,�< �<-.}=0 ,=f2��[\�@��DC�<d�y��_��wI��7�<�)��3<y�^<4<f�#�U�<��^=�ּ�����*��U�<�
��<G{@�jU-�4k��ܯ�i�-�5��<����D�<�
异��?A�<�]=Ɓ�:k�6�=��\��0<�.J��A�;X,��k뼁�<���<��=3(�<o0����E{����<f'�eh��-��;dXU;*&I=]8��<=��7�T��;�7������sʼ��y<��$;��K���ۼ�ۄ��|A=�d�ٓ.=T_<��<
=��E��N�����<���A���e��<wK=�� =%l���;"���t=���<_h�����l�4���]��Ӟ<-�׻i�;��2��o��<s��q�;bs=�
�;:�J0=�Rq<�:��=l�O���=�VU������/�J=�yʼ^��(1m=b@�<��<Cj�;���<�<��J�`�k��n���6=ǅ��-�Ӷ�:���;��<f^�<�ǋ�M�<;k=q�
=��$��M�<Z��<?b=3���s=>;p;E�=�
�<wZ	�rZ|��G:=�i(��F&=Tq����<�=f�伔�D�� �q4U�e�<>D��5M�����U%���=���}C�;r~�<0�;���2`�G�Q���<���Zu�<�K���0=��B�q�?�񉰼��8���\��U���l�<�c�a����:j����<d�l���)�mQ>=�Ü�+-�L�<�j���u��%���X��I2F=�U��,D;?��=�Z�;v���3!�<��_<�	�<�j�<ƕ�<Q���(�:��l����E#=��7=06����V��o�<���!�&��H?�+���$�B�}w��7G=��FV����;����7'=g��<0l�;�m��#F���=F)!=�I�|v��ܼU�<i1�<�!�(	=a,޻DxR=6>����=Ǯ=�{���:=��M<�MC=�襼$H^��wD��ͱ����<�i��^��#G��:<�l6��� =�_�<�=�ܼ%'�əx�z@���W����zob=�]��������<W`=t�4��'<1ȓ�[=�;�<U�7;�=�M7�儩����<��S<��0��W�<���<��u;;T�<�`ݺ1*/��N�n����Z�;�k�CvP��sf=<;R=�k$�B��<>/h< �$=�II<��-��*�3�+� ߟ��Y���<�E}<,��;�zH���=
��<9TQ�y�[=憺�V��g8��a�=3Ps=[�C�n.	�Hf<�м0'
�0ln�Y�<]J�<FO�=޼��j���<yB8=i�=��=K��8.<d����#���=�J��6�a���J<7�X���:��.�l��<�乼C��<|�X�kd9=nÄ<[�������*����'VO�kî�8��m�>�L��rU��9��
����<>V=��P�?�P�;#=1j�<y�=\(=��=��<��]��n@�Aļ�A���.<(�ۼ=�=�p=�5=��<��=k�Q=�䝺L{�=�5<�kH<���KH�0˝����[��;wk��no�zn軐���Y<b=��2����s`=R��#}�_�b���M�M�<'���S�<P�<��H=���<��żC�=��=s�-=j��[='#�M�	:,
l��I�;z��<|�:A�4����������	=�(��'�<܆><oỆF�;�NH<��3;.GA��z>;�ۥ�����/��ZP�T ���\m=��S�9�v���a=f�=@�-��.��BZC�`=v�%��:eѺ8J#�X�Ҽ,�=Y���m%�n�"�����ۍ׼y��;ۮ����<��$=��D=�S,�>��V/_�v�*=5�S�p���?=Pp���D�<zQ*�_-�Fg<��.=+�<�,�;��<���=Ѷ�<��y=7�;�E�<��]���=m�$=�dW�O�=d���P��C)��WT=��j�
��<hj�<9�s����r�H��@Y<�<#%/=T���a$==���<Ω>;
`�<��@��$=c�<�+��T=���<"��<����H$e<#�,=fo�<�]��9ü��;�\l�<{�F��(�<o���6�=gt=
iE��
�<������<�����-�NL<��<NS�iV	=`��1��S�j=�<��`8��I�$x�<N��<�l��������e���v�U�C�8Б<8�<��@=�q =U�i=���<�':jSc=���x��<O�<�T����UJ=�9=�Mw����0΃=��W="�A=��0<9�,�̳���z =�K�9YwȻ����ۚ�P��<(-^;o�g:�*�����:�
'=T�<��� �#=%[�)�eEN�ё=ڮ;w�	��3���n�=U>R=� �
���G"=$��;�1޼E��<:X�cX�!!=�h�;�����4[=@`�RB�9SF=�/5<h�ϻD�Ӽ˵�<��9� �<4����v=ap�<��<'[��=���ߦD�2���Fd=�x��X<[;g�02`=d=�b|=�Ns�x4��2���&�$��	��9��	��f��N^=f^U� f�;-\$��5T=: 5=mY�;��%=-�w=�iA��u=A����v=q���n�;��c�G�W=]�=�ī��7=v�<rF��O��;�J�<�:��o=��h�P��;Jl\�ϱ<"N�<�?=1�N�#�=,&=�@����f=pB=�&���*��!���2��h[:<�ӥ<ݙN�,�G=�W�;��C��R�<P������<Ԛo��
�>V=g0��"<�RQ<��+� he�U2/�N�A=��S=f4P��c��໻���1��	<��<���V�hMa<qC��;Լ��OO3��n��s�]+�<i��|u=�W-�6��<J=�`O<�=��B�ƻ-��<��=��=+k�}ؼ�K=$����(o!���e�*ڼy:h�5��zY���h���9���Ʒ<G����&=4�ڻ��H"= �b�eʁ85P���<�#=�qἭ<�.�Δ�;����ʪ6=N�м"[�iIZ���=�� �������<N	��%��;D=[A�W�<�ʼ�Ȑ<m��vլ<��1�;�Y=�� =O)=�zv��ʈ:p~�<^�\�!ܼ�i�<ϱ==ȝ=����H�m=QK'���=F���R��; �s=�����<�<��=QE�<#�=������ܠX�1�s=�ꔼ��=O�<�y�M�N=�_ϻX�2=)���<��<�|�<��B=��~��<��e=��Ļ��=��E=��=u`����:�:��;�Gi=��<��9���*�6-<7�=T,�֢j<\= ei�a=�<�K=Y���+M;���<��a�w�;=�Ӛ;�ּq�������D���� �����=���=��+=S:C<������5�����=�g�<an�;�<�t���萻����Ϸ;:����V=�`I=�<��=ۆ�����<)�=�=x.�;x4�.��<�_�:v\!=H�C�X!�;m�T=g�=�����2�.��<��*= x��L)��=�<'�?==�=5�<K���#��w���4=��<=c�:��q=e�;�)E�6���,ۼJ�Y<����,�<�=:�/=��G=��?���Yo`����<%��;ܿ��м<hR=�O��
v=f.=���06=)� �F���t=N<+C0�7Q5��h=ɛ�;N|=���l{U�����**=����dY��<o��b�d<p8T�(�<؂>�.�*�ʵ�<�k<=5=b��.l)=m���!%��|�*��<%��;��<��S=I�3=a=��s�_��<��,�/=�vͻ+����=��=���;�����B<ը�;{��9QЋ�.�.=��:SDۻ*�8��r�(\k���|FS<�SM;��������O;��d⤹�������Cɼ�̃�BL�=��<��J��;�6;�(���M�ڡ��]z<��:���<�ȼ-'�wԅ<{�4��0�<�e�<g�S�po?�/A=�y�N=3��}H<D_*=��;sth�>!<j<5��ټ�Gc�+Ǽ��@�j�:��<��{�=��<�Y��&�;yz�<�T�3tϼ8J�X\
������m=\��<|!��׼\{�m w;!�=?�/=<��<����V����<di;�9��<@Gd=���5n����x<4ɿ��b<������<M�Z=�����һ�6=��<6uY����<qQԼ)Q��t=�D���	����<,=��=�ed=�8���e����<=�(=�C���|<@=ob�?=�ey���'�V*7��o<��`= G�9�����i���-<
�=��p�<wgB�&�	�g=�m �;�;�	�;o��"N��L)�b�����k��k��u��#H� gQ����o�<�n�<�(=�څ<���<� �<�P%<��<�e;[Gz<��������C0Լ�O�<��:y�^��Qļ؀(�d2�<���������/;��=�=A��<כ2��Em<Q���q=k�=�hq<T/:=�=?=��<<�]�AMC�947=��=�cC�^�1���U8=��\<����@�<��<��=<H.��"���g�V�y��g�s�<�%M=��=�s�<�B�<:l8�#wf����:��<�����N=xm�U=���[�<ܚi�~k���D��+R<��X<�)V=|�;�S=:�q=�t=u�|��K�p��ss�v�<�2���=��ǻ�}�9�B��:��w�1��)�<r̄<;�ۻ��Ǽ��H��Ł�;￼��*�嬵�h�Ѽ���:��ͻ�{L����<�N��zF=��j��M�օZ=m#����:ԇ1�}����я;q����=���<�׼?���=�c�&=���<��W<*è�s�"��D�<�g��\ϼ�β��1;H�6=0�J:��<�.;<z&I<��<#�/���=�h�<H�N���P=�� �*F=���<	�]=�n�<�ޅ�?��<ڀB=���<c H=ր?=>�缵�_�T�I�Q�L;��<6��ygE<�`�_�Ǟ�=����/�ۼ��A������+��&=w��<E�c=ߋ<��;�5���� "=}R�;b����~���<�L�?�e��|����<�=�E�3���1b���%=Ѿ����E���=<F�F�������F<��(�P���<�oq==}�<~^&����lл<L=�c8<D�<4����/A=y�<�p=�m%�9Ә=Ǉ[���;h���N(���=t�t��.��d52=:� :X�[=�ü�a=}��<S}G�v��<��Fm�=�>A���
�{�S��	e������ܻ��G<<f=j*�����^\<{�d��e�
\�<��<##�F���H1=@p:}1=3�=�ox<0��:��<F6<=D-�<����P��b=X.�<,�=)z�;�C8�������[������f\�:������;9�g�\���2=m@<+<�!3=/<��D=.��<������=�
����[���P�d�<&��<fd����=�)I=*�_R�;���<�Ż�N��ro=�F=ܥ<L�4;V�g=���Z��<���;-�h���c<K	@=��-9��<��z��}��[�R�?��TǼ�����t<B�;�qǻ�:=�M�<N�;�ӪC=�;�ɶ�?֒�1�1=�Q�<܎�<�w��� 	=f6F�P��<�x��t#�\�=��:^M�?�&=�;0K?��
:�c�<��;�&��o(<�/��� ���Ƃ���_�hɼ%�Ļj1̼�+���<"��\=� =�w+�0~�j%@<t�>��0Z<ܮ=��H���s<!BL����<��;7E=�L�̄��\����q =�0׼�nl<�%�<Go?��4P= ��=		#�5'��0R=k{Ѽy7<���� ���Y=@A=7�B�E�<��B��<����<o\U=�/��	;�a:�;vo,��w�=��8�H=yq��%�;J�I�fN=<Qs-=��=��F=R#=�D5�8�C=�#t��
X=\n]�+��!)�<��p�$=X�1=av%���)<��2��Ԝ��t���,�r�<o߾<����,�f����B=��<%��
��<��S=���<�s���d�R�o��L��i
=��<����\���R��Is;���<	l��.7<���<�;���@<�4�<�8=���������<at<="@O=���<��i�E=�?Q==k�u-J���w�e)D��CʼQ8���=N�:�a=�ソH}j;9>=Z�==�yk�#���'w�� <=+���u=���?�/=fIm;�U6�Q�!=����=���<�>����n/l�f����B��8{m;�"�$�;����.�;�jK������@2Ӽۋ&���{=�xG�s1=)�5��2|=&z�:*=���<�� =M)���N.��(<��<��������7��<���<ƈ���R���<�
=��<2��<]^��y��n-=��7	�<o�t<k�<��<oq[��;�Fr�<�U���:�<��<�/�<��_�vX=ʛ���,=�ց�$����<�����r��Sn7<4
=>:�<��<'�ϼ�<{�+�V�S��w=��"=�=.�+� ׼���;�%?={��;E�@<����]�U=�ꄼ�Z�A�h=�K=�B�1M����0=�A�;�?��ЗR=��w�8�+�3�j��=Ӎ�<+�
=�b��v�*Yp�gs��1�F�c�={�5<��<�3�:�bȼ��=X��<�C<1d<�3�� �ܻxZ!=�@�6&z�D<䃩<��ؼ(�����v�7��F�������D��%���h=��<N9 ������9uF�U��<�+(��;
<Q>��͎�<V[=w%\�>X���m=�¼(^�<g�z�[.�<��;=�I�D:$�l�09|=��r;i�1R�<�r5�7j��(�;���<tNa=B}�;�'=�*9���= <��<�� �4��<1|Z<�\	�����(=�ه�ݜ�<>k<�9W=[=A�x�Z��1ݣ��v�<�Q�< !=�Ux<C����B�֭^�X0���\C;�mE�P4��;��� =��x��W=��(=��i=�A=�x>�>L��=o=gb�<�!�7CN=��,�h�k��bV�]8=$�9=Z6r������L#�<�nG=�2h� �<�üK2�zZ�<�]�>_�s�==��==R!��b1��p.��O����/<��k�~+B<=E<%%=�D2=D*Ἔj�!��<���<��J=��O<k�8=�iW=�@�k�r�PlX��&�;�B��=E27=�<��_�ȼ �<��߻<ȑ9Mf �%r<�V�3�`��C=�9D����S�6A�<���;'M2=�7=�d=��=�:=%�I��9Q<����|��<�W=����;$�UJ=��+<�-���
=���!����;��A =�%
=[�߼� ��ۀ�;ۉ�<��'�w9<5e�?�\=��;�[�<>Y�:��=�zü�.���3���=�n}<�e3�.��1h�<�1=��<�
"�Ij���^=Ċ)��3��{
<O��J��;ϥQ��"������񼩩
=����P}X�U3��\�;�(���&=.����.�F�U�w��=:p�D&=<�=a��@%�����F���:�{T�����Q=���8�=� ���D�]�<����v1���qn��=�(8�
YQ�C��<�������=�#h=čR=�o&��#E��]�<)�`;a'g�F��ѿp=7g����~D=I��l�X)N=Y�Z=����_=������Fn=��3=8D<��(���e�<�껚ջ�w�I�]<�\=�.=j|=+��<)JZ=P��@��U��9�<m�<���<��G=���;+=4����/=oI�<� ��77��3'=7uW��q�<�>y��8g����<�n
f��33=ĥ=��a<!%�<l�(�N�<�H=V�8=��v=ġ�0V�<� <=�T��rU<�F�<�H=m�<4�4<��ѼT���a�T<q�<��Ȼ/f<�3�!�;-��;��@���!z=X��;�N�� �<qD<�Zb�(����a<�7�<��=���*���@@���$�25=�>����kcf�e��<<��E�1���}�O$M=��L=}b�f�ؼ;xk=;�4�94=(�=G��<�*	=�\��gc[=�T,��=>w�Xg����=�-�Ei�|�]���<����<�	*=�w=!!�<!F~�QV�����D�<3'��Qg=	k��O<��l�+�<�ڦ<��r�G�Z�c�'��~�<�ʸ;�)��0��e����=}��;��<�6;�@ɼ�\�<|F{�w@_�Q=�����7���s��R=�g���	�o�<�HS<�'L=��V�&կ�B�9�,=��e�<B�E<�'=�T�<E�2=���M1=��_<I�<|\�� f�<�T�<��M��8�<��2=�@-����<� <��ݺ�h��kH��}��s$=��<�gU=�3��u7����<�9��ü�\�%�k�^�Q��tE>��A+=q��<�+� >!=��t;q,=aw(<0� <�cd=}c=pc#=�Z��к˴ټ��=a=��<2 F���<&�e�'=�T�<L��<*�������م�<c���VF��h��z�CY=:�<��ϼ-�E�Ɂb�gC=yPL��T����:�3*��Ն��*���>=~	�;�O��h=Y=k#=z6H�딼*����F[<�nF�� <M���tx\��@&�pJ:=��]<eZ��G�	4��v�<)�s=)���2=��=_=!K��I��<&=G��<|�6׉<�=�f���1�;f�]<����2���<�$=JYr=�Ԣ<.�#<JE<=�X����;�L��g�Y�Ԟa<'9���;��=s��;{=߷X�8~���N=,M =�?�����i<+B���*��!\�<W@h==u�'n�<2�ż�j==�=��q<Vu;@�v��y��_�<[��<B�=OlY���.:$= w�=^>=�]O�t�F���R<~��<�İ9�HO=	=O9=�=� <�T(=Z����+�/�)�<��.<���<+ED<�"��VD=�~<`��<$]��=�P��iI���:5[�l(@�y�'�񎊻wsH=L�ü����A�:��<|#�<	�#�!q��０�K=�;E=�xu:��3�r�����x�w=r�Ȼ$=���<$�+=3~������Z|#���2�3̟<���<�c<��W�F�]=m�8�[a�:�?"=c�8�cGm<�7e=�G��kT�u�1���=��<&B�J"ۼ#5t<�����<��<�;a���<��<;�@:�2�I�=Y�O�~C	=���������A=;A4=I���(�<�i�
N�J;�;���<��;���<�*�;a#ּKiS=�9(�K|I�E�2=���gPڼL�_����<ȹ�hy�<��=!a=��ؼ���:R�6�5;R��'<�Z���z�:�3=?:=�^ɼ+<;�?<S[<<Ag</�z��	�<�����?}�A��96�<���<�D�:��=�-�<�z�<J21����<'�]�z�]=d�3��m<�B=��B<�r�<u�;
���J� =z%}�#R��\ �(cb�gȁ�����V"�k4V=i�ݼ��<!�+=�5��f�<��=�!<V�_�q�/=�-G��qf��:Se:��C��=uH`�K�;��/=#��;
u���¼�D��<�kH=1@(��v=��d�t��<�&����Ha�[,={�;�a=�;�#�A<����P�<b����<[��<PN?=>�$=��!��9�40=v�Լ��S=�B	�V;^�9<��J�~<�#�<��M=���<���<�|$��� �a�j���;N�4��<WN��(X��@H�h����<&�6���=*�0=w�<cNE���U�F�Y�A�t|=xJ��*M�<����)1=�@\=c�{<�����<d�S<��G=�H[= c&<2D���<�&�<�<�����q���j�����m�d�T=/�<�ĸ�3Z�<�Ҿ���B�Y<�\=+Je<w��<}�L�`+<���<l����&C< ��<��L=� ��i�#�
�x}ܼ�b��󃽗�=�=��Z��t�������<%��	������D�;��%��L��k�/�`}W�=�R� �ɼ�(O=@¡�?a�<�{�<_�q�z7j=]1V�P����#[;=�[�;��<�K�B��<�z��6��yO=���z�7q��7V5=i�T;= ��<ā�H"F= �{=鏽<�P�<��;<#���4H=������L_���<��}=�o�)�K/=�Q=�ļ�l�<�!���<@\���;�9��ͺ!���u%=�Oۼ��f<9}=���$H�<���<��;v�e��Y,=��=�=�x,�9�U=��`<@a=ð#�)>����<�@M<������=��P;�T�<E���ݸ�09�<&U�����nm������w�k�G�H=�|�i�Z=}�V�ثj:�a�;+�5=�Q=W5E�݅r<����	G=� ;��4�yB���\<ѻ;���=�
��ef<N	=���<h�F��Q����h���%�2N<�Z�]��H���_軼��<)�J�@�3=[=�<�=���/��L;�#$=d,��=�꡼��<xJ}<���<[Ĝ�h�<"�"�d�=nw�<�x�9�<��h*�<�o=��&�2�]��IJQ=�렼���;�]����<(�B=A�=�#=��Z=Z����1�+�5��"�:��=7lO=��4��?=�d�����=<�zO��,�<�i����J=M�*�~E����:D��<���:��=כ';\��� =jb�;��!���;jvU��n컝��Z�*�NBU=��H�C��=$�<<�����=x#��$]���<�p0�<����\=ȉ��,��#=q9.��Ǽ
�9=��̼l@�P������<�"P�+/�K*�<βR=�	D<̈́�<�J��q��F�=��I��+�D���V�=K�k=�{�<b(G��;^'m�D*�<��6��\
�)������;hU�<��ؼoa�<���<�f$�,�<ӨY��[=��=��������μ%�<{�-=G2^<�����W�� 7=����\�<�6��@�KN=s�<�����d+�,�A=���<��=�w��5��<K�˻�%=ҝ=�dļ��=G�P=��L=�)�����`=7�~�V�<J�[=۰
=�v=��]=Ye;���
<Bx�<<�<�~��9J�1q;$T�p�^���Y=����R(<�v��,}h��a�;���<"|6=m ͼo�ɻ.��<��=�$�V[�0��<~[+=B37<�:y��o�<���=Ua�V�%�A����V����;�<��7�/�Ѽ<�[��g�a5�<�G<s�>=j%<<ք<L���%��}�мCW$=o��<G��<^d8=�,;����8�8�]�O7�=Z�<2v�<	�<=qu���S�28!=� V���V=��)��_�<�p�<g;M=��������d_/=]�<P��<�,��]���༼^S<��^;��o��M]���<�_�<��m�1=�f຃Ts�t揹D�"H4�4&==t<ӂE��E�<��1�n�<¾�<���45�<sRu=K̼����=Vy>=�	�<&��<���>�=��=��?��=�-`�T���;};~�y���U�d�<��}<�JN=}�o����<|=��J=x!k�t�9=��&�Ӆ���>��PF�I�<��׼���<pK�����<!EQ�$)�<�=�kM�A��<�䑻�0^;��=�[=+�_��^<m*��wZ��g6:������Z=Τ0=��< g��h�yP-�w
�?�i�M�p�k+�=��/=�[=d�5����<%�;�E+��ն<�/5����<�_�:���<8=���q X=�<�=|���ϰ<��A=�~�=�<��C��Ǽ�ζ<!��<�D=���;_)�:w]����(�E�K��绵�-=d�8;��%��B�����V����=����>=F�1=���ڿ-=4J\=��f<�d��=]= =��P������ ��Gۼ�Y���s-=�%�<��n=?�"�E���+�<=�ÿ�x����<�/������Y:�m���� cǼ/� �Vo=�T���9r<zC-�{uX����<� 	=�4;�E��<$�=�*q���3<���de����;{纼2bG��)�<�ﰼ�\���4= ��W:=�R	<�Oe�*�<� EF��?=,A��u��[Z��5HN;w�%�%+�K4R;73i�	=s�O=��"<�nQ�T?⼤�<�m�:|	�<��5<���<��Ӽ=@��EϼpJ=g�=���<nbf<O�=7�O=�RR���p���fs�<�Z�<l�;��<A��<�ռ��<K68�����ej<m;_=$=���x��1�<��0=1X=�0n<7�p����;c޼�۱<��I=�8=9?&�W~�;k��L=��+��!=S3��hy�=���<�==��P<r9|3�<K]���=��5�O��<��7=0���L�<4=�'�B��<Jq<�S�<V.��>l,���9=�s�<	I= 8���+<*� �
�����;����/�>@*��Y= Q �_�U;3�^�=ѕX=BI2<��M=��r��Is=���<�b';�#��.V��-�<�@=�T+�@��:(O=�y�<�&;��e���<$.���k�x/O=�1^�(?�<8��T�s��<��d���<]�<�A=���;�����4<Љx=$�4��3�8�-����wJɻ�<=�3<L�.���g<�V�;�Nb���
<��K�޻�U_м
�E��3@��O=d3u�#?�P~�<�8��j�=}�==�T ���P�J(=��<�e�<o���\�¼�
�<�1='�U:�ȼ�1@=���i�C��+=���;�Ę�7ڝ;�6/=��=�H=���<��l��=��O��p�<WFd=�}F���3�݆~�7�R=�g\���$=VVB=��:�=�u�:s�o=3�=��<��t��F�:�y]���/<_ǘ<���<�֟�Λ=��8��9,=��<8�'�!���мT��;V�\=��<�<���&4=mxr=������<�}N�(2=��c�_5_��'�<}�ʥ*=1�h=��6<�o��5+n=^ؿ<��<��:��T=�Og=���⍼UZ���/�7��<k#C�'�=�[���Q=�� �s)B=�62���W<�BA�(*鼄K�2h����'�m��!�<�>ڼK��<�t�ۤ��=hh��gҼ��t;��Ȼu͗<�����W=Pۉ=o�<ϝ~=�2$=�6_�P6=~�<q�G=��=��:��D8<$YM��e=۴/��O��R��<٣�5�������<ʎ�<n<\�pX��}N�0��<���8�iS1��|=�_I={%=�|V���`�Q�;>�I=��2�U�]�<��j�R��vU�<�m�;�=��+�-e���U<՛�tS;��Va��R�<{���g�,�I�wG��y��(��iOλ�T�|$�1`e�W��<s=i1����*f�]h<�mt�(��<��H��l�� =3Q=���<��I��`(�hs�<���<���<@T��>�=�3<�y��:��<nq<ֲ���<�$O=p�
���o�3�~<�5�={GR�j�2��G�]��!W=Q�:=��=��û8r�K��:���;��K=p
={��L�=�J.=,0�<.�=���ا7:���x0�<A('=�a��5x=�{M�e�k�CR���v�Dڹ�A4���=��<�3�<��k��.;C>_��E�P=[3�<��=I�<�E2���<|�<�e��2�&������<wB�ʸ<6�����<�F=w��;�L����g���R�h�<`H�<��ۼ#Lv�%$w;\�1�.�i��l+��8q=�7=��V��	ѻ3^�+X�L*_<݃�b>�=!�<-r��V�<��\=��.�TJr�G�3�{�ּu=�e�< ���a<ˀn���A�Pp�<:e2=&��97h�l�=BBͼ#�(=��.=2���au="d=�%i�Vif�����="�=��=�	�<S<���<�i
���4�k��<���<"A<x�L=X^����9�x�:��vj��r�D��O���=Lo��^l��
TZ�EeU�g~��3�;m񈻟�ȼ���<Y�<e,=�*㼛L=mֻ|ˮ�LdT=L�&��07�C�|<x�<�xO=��/=�\3��D��Q���&:k=Ԇ�<%�j=� ��݂�������F�j�o<W� ��A�<+�)=p۟<X>�<T�=�0<`�[��&+�� �S!�ћ��`L=4l=SX���*���<R�)<%Ә<�ڞ<y<=ݡ̻���� �:��;	��=�g<�5��s��vZ5��y�<ȁ�;�=[��Ǆ%=���<|ꂼ��X!$�@h����=�M��7&/�#F=s'��^=�<=��\�s<�(�;��<��ŻC�=�<�<�CF=�H)=p�I��%�;i��f:�D����&�)�t��< g�<�o'�����n<��;W#��,:�d�,��:�<�H�<O���v�ü��j<!�߼��]<.�ϼ�q�<�hm��6	=<��U��_=��`���t<�&C�!~9�	뼼
���hü$��Ϣ��.�2=�\��h�<Y;p��Q=��O=�ب<��D=u�<��� !�=���=q=n=P�<J#=<{Ň<���<�=C�=��$"=6�C��Ȝ<mV���������:̙K=�h���<Sma�~�3=T%=\y����;cǜ���>=�L=ѱ�<�*y8���A�v=5�켌R%���
-5=!�<�aϼH��o	=Br"=%��L��<�p�;L<��ۻ��%���	��.= �J�����$n�̉0=/����k�i�Q������$;=�M��8@��!M�?x=S�f=̣��*��qdM=4b5=��<=��{��9�;̕�<O	
=�Ğ�m[�<k�����Th�������-<�'	<7IZ<=�:L���^A�_5M=ʵ�;.���vxc���켜��u��N�h��9�9
����;�6��[��<H��;Z	i�؆*��n��eU0���=�Q�<��ͼ��<C>ڼ܀�;�C�:�~���)��bJ=!�=�m<�EԼ�U�:�=h�.��W�
&=�q�;��[;1Sf��=y���s1=�'�<��9=�0��;mW��@=�q�4)�;S�˻n��;c���53=��Ǽ��g�o�X��<����+��� = �= ���A�A���M�*����<���H=��<�j��e��߾i=��b��<���Uo���<��9;�¼�x:]���w�[�p�w��jX���;���(:4�����<R<�<�YӼ�zm=�cR<�h<��@���U=:H�����'�U= ,�V<�rJ<3�Ǽ[��<�h=p!�<��@�>�=&�?<%ɚ=�_K��r��FP=���͹e<X�I�"��<��c=�G=��==��="��;@KW�v����*<?��<�8J� �;wsm�x =�?+�����Im�����ɼ�HW=��!�<�_��;І�9�<�0=?����ϻmF<ڮ\�)�2=o=x+=��J��f�8��0;�2�5��=!��<Ch=���揼ր��F�̼r8��?9�<��H��=rhj��0'��II����<ݛҼBj���K=��)<%�'=�F8;�/M=鴊<-]�<b#\=a�n<�MK����^N=��/�Q�+�;2$5=���<��D��6<t�S��!)=�����H=����1��w��W�:=�"M=d��<T񻼖l��D��<$�_=m���|=���� \���9=�`z�|:��lD>�Py�=�����(�s;=�̜<��8=����4���e��JM�]��<P�¼��<�}��=�v0<��p�%�<�k�:�<=�Z=MV��lw=��:��<��
Y<b��;������S=� ?=ɏI��/J�4t�Fe&<}�<=�r�;�U;?�
�,AF=£S;m:;ʞ1=��F�<�a=R��<�pe�c8�;p�ܼ��]���=D}���C�>;��%<5~Y���#=B71=(�켆���eN�;�j=$<�
���P=tQ�<ݳ=��1=M%�;i��S-q=�����!=�[�<�^A=��Z={v�<>l�;��p<�p=sn�� t����o���,=W��<�P<�L=������1���+�el��S�i��gD��n�;}N�I�0��߰;��P=����,=�_׼D�A=H��N.D���ۼ��,�}[=�p������<�*l<��Y=ԃB�%#�<u	=_Ɔ�=�	<�{������]<�k<c+=�~�=4�����<��>��u�<�45=�5� ���۰�<�L�c3K<6f,=��<
$�BD�!|��#<=sX�;E.{���⼤�=ٴ�U�<̱���D3��b=
M�����D���O�����;2o�9m?]=)E����%�~:�󘣼0�D���=΂:n���,��h ɼkL~�B=kq�u�/<��A=�i@���<I:+���=��:}$0<CxM���|�X�T��<I/e<f�ܼB�����<��;��� �^=@�h��DQ=-5<�w/=�R=6�)�3��<��L=�b="�/=f$����(�,=��z<�x�o^m=Qk��M.=:7��O�w�Ƽ�M<A>G<ݭ=��������[�;��������t���x��[=��%=�7<y�=$м+a�C�v<���<_"= ��Z����gI=��<hG=wt�L���x�c���F2G=�ŀ��?��r��K�,�\?"�(羻��b=��E��w��b�y�G<�z;��b=F��<W�=T�:��.i����p���=i1�!���4�<��Ѽ���oPP=��;UZ<� 4<��?���ʼ�pj=��<az^�؏<?��<�dL�:��<��8=�O�(x��F?�J��<��=�=k�;�Z=�='�o���=���-�<7�5<�����<9�ںR1\��\;��m����<�����Zf=�>>=��y���,= $_���=3k=)��<q�=���:��=�[��R(=��I<u3t�`G8=o�;��/��2<�d=D����v1=^U=A����^�Ÿ�<+==�p��n	�E��<�Gc==�<z�¼@�ֻw�^=�=g�7�=���˼�SK�v� ;�<>1= ��<�5U=2!�<  ���u�f��<�Ǽ�zp�[O�<Z�z<�<�p��+N�v�+=��\�����T��V=Ź�Q�A=Bb<ĵI���
=����H�Ƽڟ�����VBq��(��`K�mK8���~�<� �<t�.=��E<іn��b��Id�A� =�r< ��Q�M=�>���d�<��]�dd����.=��<�O=Gᮼ����R�.�AF"=5��}�N<O�;�0J�:^�<�s|�gv{�O"����`�c�<�=�3m�U[J=� =E���=I��_=���<-|�<�C=.���B=�㑻Da/�K�B=���<���j"�����lK;RQ=�� =�B=D鿻7���g�e=	wJ<=;�>�<�t-��NY=P���n4=�c�:֝꼿mq=�����<�� <��Ѽ��6����<
��;4l��i8�v�X�<u�<f�i=�#f�ȿ:�I�s�dK��7=��;=NM=Cl�;ɸ=+�	�j�5�+�;C~h�_Uٻ�4���=* =��⼶`0=@�J<�ȑ��D�<�E�=ܳ�ܳ,�3�\�Ǝ�<�b߼p5L�)L���|<d�:�ŏ=��-=����cb�<� �=�<)�=�D��<â =�\� |*=[2\��1l<�4�<n
�<r�̼Ɇ�<\��)g�;/a<CS�<�<\��53=V
�/)Q��������t=2�];��q�b8��p�]=���<�����=m�<j�R=��;��5���H�U�;^ϥ�H�f�]\;U���<��f��=�G�<�5���x&=�ꇼ����=�O����<�]Ż���:I���E��ر'=̲=��=�l(=~��6|�d&O�r2ż��=�ť<T�\��#Ѽp��9>�5���8��+�<�Mټ��=�'ϼ�ad���'�%�<��G��rS�3L*������E!�<v_*�[�&���8P�;Wf@=�+#�,��;s
�<ʞ���ǼL,=2f0=_��T{+�
k=����B5<p�L<�W�����!⺖~�;��<���<r�Ѽ�4<���,iy�n�L�W��<ٳͼ/G	��-=����6��<�=4F�:	�c<$�V=7[=���;c='y�;�r����X�ƌǼA���v(�a��D=��"�D��<�W���F�~v��tn=us	<���<W�;)Q��G��d�<=`�w=�C���-�7O���g�;�rV��_��)Z��#ϼ�1�<|/
=�a<�4.�%���SU�<�컻Ģ��@��HD������t��<�?��\�Ӽ9l�<�	�<�XB�Ҥd=v|8�����K��#�;<-<�H�a��_�2<L0	�z�b<��<� ;~�����1=�zd��<w�p�}`<B�=�/=�:��Cw�=�Ŕ��у�~=[.����<�~7<F�;�� ]�7_߻���:�0�	=ے�;��<���8�[<>NJ<�:»�{ ;�א����;��.<�`	=��<�X�<����<�/���^�;�Ӯ��q�[�7=]BR�Z|1=��=��]=i��f�n�gH =��)=�����������<Ƭ=�,<H!4=�g3=flF=���<��9H��q�o�t�?�q�րw��<�T�_�JE>=j��</�\��i=�����T=);����;�jZ���J�V���gaB=
O���E�3x��K
�[��T��<e �=B����T�:N<[=����H��k=]������T�=�\U=Q�}<��N; �<��=���7����g&=��a��F	�I�=s�=�r<oz�"�M�R�n:���:��M�V��<]��A�V<g63=��s���<�P= ��<v=�&=�)���,�u K��� <�k=�֠��K���0z�>�m=�
3���>�q~���򼃴j=�s���T=kbI=��<�'����.�ͻp�
���;�<5��<o�=�=�值�빼$�Z�)=]������<&�J��.f=�_=��=� D<-=N��<+c<=!G=ۭ�;�8���\=,=�\�rD��37�<}c<���;D�r"<\X�����n�<8'�R��<��:�%=�� �O�	�	�h�m���Eq�	4��U�<�Lf�)���a==l}=OTq�"�m=?L1=aM�<y0�<�/�8�,���<-��<>L>���{=������żj&�a���`�<O�!���<�{9��sH=�Ew<��ּ�7:s�k��jҼS¼���e=�;�<5�<�&������VR��9@<u��<��,�@�R<Jb=`]1��4=����W�=�
:=U.F�ZJ=��"�/�R��<�o�<��=1�e=�=����p={���>�dy�R=l�-=� B�z{�A�b��@<��B<��U�+g���iQ=�e����<�)b�
��!��	�	��b���K=�~U���= ��_�3<G�<8<��q#�<.~=�C(=��&=��<)"�f�<�V*=�e�<����O�8B�$�<����'���}<��E��lc���8��s�:��c�L�����<ٯ��`���3<:���zk���\R�}S��-�ڻ��M_;=V5������87=3[=��3����<�s�J�<1/s�|M��P�t���Ӡ�ի�<�N�=�7!�d��;J��]�9��C���V=�<����y%��C4;J=��=�n��]g�;Bs�<��=��$�>E�� dQ��*�<J�;?ee��D��;;�>���Ӆ�kxI�Ċh<���s�����zc<��<���;���<?R�<�h�;�R�<��<Uvu=8WN;����=/�=n/�</
�tv*��P;�Z=����c�y�];�h==bs��R�\��s�;{�S�����Q=�i?=� �<��#���i��o@�"@$�ge���I`��8�=��=�rѼ<�?���c�1��<��ͼ���<��)�)�=�j;�^����i��"�;C��;#| �?�<�=DvY�L=H�U�cN���7P��w�<� c��R%��\�;�U;��X;�X��ʳ��`*=xK�2���� �)$+=��;z=��<���<�R�<W�S=%T=��¼9 �;�^F�><[�f=��+�IY(�us���W��.=(�o=K��+~%=����&W�)�$�(EH�c�6=8��O=gA<;/K=+��<mN/=h�-��]D�^P==��<j&�<"��b�<���<�}=�fB=^L<�`�(��������^=��5�wC\�6�=��,<�]96��<fm=l��<��b��<Ԓ]���.�n89=n�
:m���6�<5�$�4�;H61<ⓛ���8o��)?�<�I(=�I�CA���N=o64�X{Q��-�=�RN�8����}^���N�6���߾�� L-<]�<9��M=�Q<�僽g�U<��m)ܼ՜w<jj	=�$�KYw< �żF7�<U�<Sz6���e<���<f�==�f=kqU�1+2<�a�;���<\:{<�If; ���:H��Y�<��'<�<��[�
^���1:=��5�"��MI=T~�<�
/=i��<�&g=d��L¼��f�zY���<%h�@a[��5�=���<UC=�YA�c2f���O���<��<��ô<uq=Ai��[=*-Ի?ٶ�J�7=3�a=���uJɼ�^	=�<.=>n�<����Y¼��=6(�<�oF=�]�:�/����;�|q=���W}*:g'�<|移'����;=�}w<l$;�ض;:�=�b =�ἐ�.=�S¼e���xƼ��"=5:��eڼ5}��yAg�� �)f�094<+
b=�zl< �
=�i<u�=�~�<��E���=�g����<��7�k�B=�ܛ<����0���G=��;�R��
��F�<3�1��W=���:HiZ�k=�N�<�p�<~T<A���!=�`��̨��[`=AZ�/ښ<��7=�K}=��_=�x����i��-���է��"G=��L<mxۼ���<�wm���
��l=���k�(C="m�;�Z6=*�=���;�|<��}M�W��1 <��^=�4�#8=4�;��������k=c�5=�<�'�`����<��=�qR�	|ʼ`	 =�O/=�x=���E��J�8�^�A�s���<J�n��6�<�=<�< �1=���<���<�7<��F<�C����<���<�q=R6<#��<N��<�r���n,�Ux�<�m�_�ؼ��z=l����Fn���)��=�־<t���|=?������)��;
�=2�U=p�"Yټ�<V�%=ɏ���^w&�!�\�*+���&��<�����<)�=�f=X�$����;9
�<w��J.=&�:��<<�I�<2{< ��<�*=`[�:��:RN=ڢ��4�<��!=�|�.�V��N%=7|);��Z�)Y$=�aU=�<d�<��n��<���<i:#:�H���5=��;_�H=|�,=��4=z��O�,���<6�<ڿP�x�=hAU�/C�"z�;.�<i�s*=�H!<8T*�',�<A��.�=��6=d�<� ���d��щ<�>�<}ce��.�<��u�;=܉�<�`5�m�T<��<�^=E\��u-���
�:A-6=#��;F[��Ds������IS�4Lo������+��Y�<<Z�<�=��;���;G�$sD�F��<���<&�; ����<�ȑ<��<�)=6�&�	;Y=q�$���<��;pb�ʫ�<fl7=Qu��CU�<���Z�ڼm�+<�S�G�=v�ʼ�u���$��+=fq�dK>=2ٸ��s=�SL=R�@=��m=n�C=N�=ֱC<�K&�}�/�Z��<�%�Y����!=�[ϼW�Z<�������58�X�W<����"�n�H=�y�<��B=�6���]
<{�k�[�W=X�i�&�;�:��:=|Z���<i �;�"�'��<y6={�=��=a7�<Zr0�ml���K=��=T��z��<|���*=���=�==��Q���S�9$����=���I�<N9�;�롻}]_� �L=��p=@�=;Ϟ�<f��: ĉ;������=�<;��5�O��<���^Ϩ��I���;�ԏ���Q��y=n��ʴj=���<x�h;Jt�<6	�<L.F�J�q�IuE=va�=K_��aaܻ�i�<0�t=���:9�=�(=(8b�R��^�M�T���7t������tx=��<�xa<uA�<_��I����������g�Y"<p��<��=�Wû*�2�J�⺶u���BX=�������; �<����.��uYK�s����<�����������C�6B��{���j�`;��_=Y���E<~��Q"{=J=1=L�u����<3��;�;|�l����9�Ϊ3��o�<H/��}1��.
�Y	�<���<L魼7�a=�ʗ��G��M���@<8�����;�)N�0T=@��<֥��$@���T���r+���,<��<�=��E��<=h<��[=!��Dx]<��,;y��`$,=42k=Ax)=�έ<�A$��&O�3���%=D�B��ͻR,i=т �+��<e/����;=���Z����=�j\�b�&���M���X���c<&ؾ��<���X̻q<�uD�¿�;�	=J'�Cm�<�����T=2�?�3D2��A+���<�ך������F=F�<E�N�;��<	g��4͊�I��0��@�e==Qڼs(=�Q��;��I�� ��4=y`�<r�3���;<��<"������<�}<tQR��BQ�j��<j0�޿�<�}�<?u8<@k(��W=1�Y��24��7�<��J=�⼌(=��6;��
=7�%=���0�=3�<-���|�!=]|8����<2�<���=c_=�̵;�h<ޒ�2F�N�]=BX� \��� ;q;�g��:P<=L<{L�<B^='#�pL����(�����N�!<�X#��P�<΀=��=�J���&=@1�ػ�� �=rd�M� �,k]=4�M�2ؙ<��E�<��-=!�=�S=N����ý;���;��Ն=�����W�\�6=��H=>x:;����*�M��j"=�TY<_�<=_�ܼ�]Ѽ!< b�<���;yxq<�s�h�$=����;��"�'�<�tX��]x<�cX<�4r�Wc��/�<��=�ݙ<i��c¼�R=�<I�U��� k��T<:�=<8���.;�TE=���<�=Y��1=�.e�<H�!��f=�ܬ<�L7��n��EF<M=D0 ��0��Z�<�Q:���n;JH��7��4��`=��X�{S%���;C@�<��<�ܑ�<��{��{�?K=���<h�e��N�y=G�#�g>0=&��(^%=x�.<�X�:��!=չ=�LF=K�_�TRټ�<���<�_2=BF=�2���]=A�X=	(l<\� =� �<Q̼����m�'=���<S!�ߵ���;=v5=`6F<c��<�Xg��!@;n��
�4=Qs��`�<�A;=�bT=B݇�ɱ���M-<�Qb=R�u<6����r�LQ���K���<O��;@0���!���Z<�i1<�Y&=-�����b����G�b���"j�G���x�;7�~���ͺ#r$=��-=�u꼚pN�7�v�γ�<]_2��v�`߫�� ��hl�m'�<�ü��+V^=����d༭}�hF=F������;���μ�:]�J=�W��*W���n=!쮺<�	�4�1=}pH= �<Xr\;�6=��=O�6;1�a���y�,�Un����+��,޼�o7��T<c��<�9K�Cd����O=�� =$K=�}J�PZ����L��q�=S��J	"=�q�bf:�ܼ�e6�}O�;�D���;�R�<�Df�Bk�[ׂ�]�=]x�<��A[=] ���k�0H����O<�^���c�J۹�͉<���ԯ��ǅ���K=1�i=�tX;����/t��&d=-�#��(Я�z�K�e��<XO<=XP�<�/׻��-���ȼ��6;\U����m���'=�c�:i�<4�`�s�<����︼,���<%g�<r�i=�,s=��'���6���x� R��z��=�<|��<��E���:=nF5=s�c;ߵ=�E���ͼM4�=?���H=�`�7�<�㠻��<}90�xj�oU�;�����L��@����<:����l�׻�=2~+:җ;Dv�:��&=(r*<r��YtѼgüe=�<�<��@;6�T���m=�fi;��м�+�<�R�<	`��k/���Լ��>=;J��C�C���<Q���
s.��G&�f�[����<S=��n��=7�-2p=�S�;��;ږ ��g�f3Z=�p:{�C�C=P�+ �\�<΅��?=�=�G����s��=d�;�Ps�����<�=�
�<i�6<h@�;���< +�<��n<<1��d����*c>��)���ϼ�����\=��&� �@��l�<��==��#��W�;�'=�ރ�Nv��-�<��/=:H)=/YI��`$=#B#<�iY�9�=T�<��O�T��=�V	����<*w������%�!��j=֚.=|q*=8/=�A,�?`�<��h=�:��(�@Z�<�.<������<���c�|;�X��<Ȕ���{v<��<|D�E{��?g!�NF	=�Po�V�V��ƪ��:ϼ�l1=�p6��_���1;�^<��p��[R<�^���[k��C><���������O�S,��hb=�Vܼ��<T��<�H=�]���Lx������1��<�r=�?R�D=�;��~<q� =�;,�r=��D=�.���w��"b��^���f9�9qH�<�8�<2I9���⼰u���ʟ<�^�<5`.��],��ϼ:�W<�=�D��1T�.=d��<D��㿼3�1=C��<�)0=(su<\l}=��<�x���R��G
=�(U=�)=7o!�fno�@P�<N~i=�0�<�H�� Ѽ���0�<�q=~Ǽr��i�M=�8=X�;;�;&��虻�o�<ʅ��.R��2b=ţǺ�g=X����g�<�6=��=�����1�p�<#[�����=� =�w������0<=�uI=+J����#
<=S>=�z�RW�3�=<XH���E��<�A<դ�<�Y=��<O�N=��`�e�9� Q�$����T=��^=���?�6=��+���=|+=G@d=����=�;�<PM�>i����
<�ε;�<=3o"=����`�O�'�>d�x��Q_J<$�<��(�
`6�>:#��T����;4p���=�<���2H=�� �Y�o<F��;�'�gkF=�
=�~E=]�d�W��<*�@=ƕ�<���<��W�
�Q��/��~E������5���<��9;�9׼���;�}� P)�L���$<���XM=a��<*#��h/=��ż�(=� =�)<�.=�����$���y=��1��Q*=Z7i��M�<<�ټ�i�3=ަ4<ii=�>�;^�&=+:�t�Q�^|
=�oS=K�<���<��W�44ϼ1�<N����<�_�<�[g�͆ѻҤ+<��}��^���5�rIZ�e����6��`�_����r@�:3����o�;ٟS�@5�[A����I��'|a���=C~����L;|�<\:����	�Xw���+�<	�3=���u?=Jɓ<;�&�R=�Z�i�Z=��H<5L�ه��k=?`=�˱�Wb@<A��h�<٠g�A�k=���<!.(��\?�<sL���ռ#���M*=y=G���nI='p�����<|LļD12�>˲�.=��n<j�k=��]�3A*=	�=AP0���0����<�3�®߸�˻�,����<��=բ�F�8=��
��/��;P���6��}^c=m=�&���������y���,F�	�y=i�t��(�<%`<��B=��C=c	:��,x=�Ig��<���@<�����@֞��n���g~<��A=�Ck=R���<Ѓa=*��;�1$�[���mN��o=߯3�o?��5��<�<An;�r*�;�=�<�͎�Cyϼ_�?=���;��8<�z��zI,���:��w�Q�V��
�/@v�)&�<���<�G��e;V�\<���L<һҥt�n@L��Ҳ;bռE)߼
F=�j-=�!�8��><=�a=W�H;�TѼ�����C=(ZB����;Nqc��9��A=�9>��%�<xJg�025=Ğ��`5=O/�<���<_A��Q��XI=t=�ͼ߸�=�k�<��@�0x�<�=�ZT�k��<����iM�vht<���<6�<xa	=~K����
=h����zZ=��4��y�+DH=z��9�g��������T<�mQ�tlм�=;=gZ=���K�<N�N�
5*�9�;���=A�Q�%g��t�2<��;v��<~���;�9��?&�z�);��d<�_-<�{�L��<g��u-=�~=K7�]~;��P�[�7�,UL����:��Ӽ�8P��;ժ߻�#�a��Q���Q��;&5 �*�˼���~.&:�P=�<��=]|K������rĻ����<��0�1�ɼ��8�̵<_�<g�<�-
��y=�<���<�U,�о<N��<�d���<fs�o�<=���#�Z�N=�C=���<Y��5=�;�<�ȼ�`)����5;5�ٗ3=�������<'u�<��(=�4(��`I����pv�+wZ= �;�ŉ�K ��Z�<�en�&�I=��<��$�.'{=��V���<���k�Ǽ���<�]<��$;c�2��I��dM=��5�ލM�$���1����d��S=��$�Wr�<�����G3��XC=��J���(=������^�оD=��d<����(b=��I��H5=�V�Ξ;3��<#�0�<.F<5�=<1c�<��~��M����<M���K,�<�M=��9���<��{=�M\=7NS<A�D=�@]=%�<sL����<{oO�d-�<x�̼�wC�i:�<5H�<G�����<���<��=(�u<�Kx�ǣ+��b�<?x�<�/ܼ�Q<��ڻN�9=�8�<�l!�\T{�4���K���#��#��=�Z�E�c��tw;=}o=�㭼t�;�jL<��E=Z�;AGa�;=�	�I��;�uM�#�+�S���<������<����^�����`=7��eI�ID/����5q�;1=�e?=���<ɜ�=���)9	=��b=[&
=��m=�0Լ�4-=�dX��"���Y�<AP^<�ɝ�@<|��S=��=�a�;S�=�uw</0����<iEG�v�켸�������z<w��<�A2�!�<j�l�7Zh=�8����9���p<5YB��=^�&=��<�~}��Ȼ��<+�ȼ�v=�=��
^�<Q�պ�+%=b}��=�-PA��NC��:=�Hr�8�d�� �2m�<&��9/V�;;'��07���@�6rK=)e��7=��&�}�@<z�<k %�v�=_��p=Y�<"�"=�x�ku�G�j��,�x�?���8��"=N��<����);"���zF��廟�׼���*�ڼ��p��i�I=�W�.y<��e=
��;Ň7�b7>9�\�<�s=��=����J����<J�[=2 =L�="��<�$�;�D��f��8U��쩨;$���E!=�=��=Sg�%$?<%��<�Y��H�k�k�_��?
��<��+=Pd=�^�=�_S�w�A�u���ck�@��:j�M��+E<��<}lA��K����R�QU'=���;O4��� ü��";8R��[R��C�~�u8�<lh`=$�Q��,=\�<!g���)'�[�r<yۼÓM�	V�<{�X=�Rv��p)����AL2=�P =�&��\e<�xN=iw��Ɖ��u��k(�#�T<�2���V����B�6���������~���=���;��g��4�*WO< �>�T�<�`
�N������:�<��ļ-�׼(?��rF��T��;</�Wdp���'��s�<ӵ�]Y��8��<9��<Jv/='� �j�ɻ���j�<7S;��k<9=��2�q���b9��`=z(�T�t��!<�{�<�W�<���;Қ�<��:�,�="=m�9�ksu�X�0<p^N�\���H�=:�d�; @.=%�U=�gV��:I��7ؼ�X=ѕ���8�<�=�q�����#u@<�*�,&M��S=����z�J<�#=¹�����܋�g��c0�<g9;����;�'�tX;q(ݼ?�Ҽ�,�=��T��ʎ�J��
I�<��[<b>�<x��<"��g<=��M��üJ�D������<N�N=){g=C�<��)�W�=�;Yo��|�8=p�a�W��=� �<�
��o=,��F=��)��)?���(���ʼ�^<U�R�u&=�<5;?L�X�T=GY�<=�d�m*=[p��X����C�X�Ի BN=;��I�@S<�=���:Q����w<��<3���RQt<22P=��i=�[����=��c=�S*����8u��պ#�0^߼.)�Hz5=EP������,=�˼)�s���V�Y<�,A=�F>=�6�;�3=��<kN=WB�� ʼ�㼙d��7)=J\�=�;�<8Z��N�=���L<��M=t=�n=�|=W 0�U�N=��R<�7�;�\A�*�-S���ޗ�y-��ݶ�n!�N9���~=I�\��>� ���+�/=Ƨ<��F��;�-�<o��< b�<٤=|��;"ٻh�t<2���j�����;��t�k��;�����=����%꼵��<�8J�v�=4��< �2=s�<���6��<��=�@&�9lY�Tor=d�<N<���B�<ѓ#�`h�<�G@<���;Q��<z�;�=�"�D��<Y�D��6�.��S)�<�u<O-=�T=TZ=9�Z�Ib����k���(���R�i/�=�@�<�G=K_�V�=���[庼���}�[�9e�����v�W��q=�����\=ve<��-�Z1 ��=o��Z(<SS|����<9J��lH���m=='��=.�L=�n<�O��(��ꄻ��;;
V=�ga=X����<}�e�D"��vA=h�E= ���{<��P<�-�<.�}c��05����<}M�<τ:ż���<�D���7<=^�<v9=�k�;E���s^=�x�����d����N�<��<n��<�ry=|=C�=s�<Bg�;�~��� Z�(6.���,:�t�/I�<<7	��9�Te �{.�;X�M�,	i=Q(<�1J�<9J=��\����Ղ=>X��'�TEJ�]t)�A�4<�#����=]����`=.My=v�9=4�3=���jz<:~��=�<�����<	�<�s�<_p=�:c��w=��<*5R��}=�q�<U�<�;�컱C�<�軺%��FE�:8-�6Z8�Y�F�G����i��I=��<���$==�8�<S�!=��'=�>�:� $�πn=mI�<ӒO�e���xZ���`Z=���_Y1��ʼI';�;)���?=�QP��Vo<��Y=�+�I�����<�"��~�=��&=\�~�K�|<Y �<��|<�<��|=����=�<cD�<��<�A<�^=���=���;ޜ�<��8�8��<d��< �J���
�<=�HU9�B�m�!�8!����<�[a;

�=�0O=2�=?R,=z<�<�p�:�l���V<�SV�=2��<���<�C7=?��:��ͼ��;YҬ=�=x"]<V��Ϯ<̧�<l=�l��;��=�"[=t�i=ʂ;�kD��5YA=�AM=+�<�*�p��<\#/<H[�=��=��=^\W�ӝ:�J:w<W;M�=%B><uT.=��W=P;������3�{M;���F�oKc<��	�\ j=� 3�(+�;B�=$I�<��3=��=eM0��Uü�jT=�h-:��M=�<��O����<C�4���P=60�<K=�p�<��j��a�=��<i^�������9�`��x9=�D�;��`�&=�X'=ڂt�F��:J [�OVz�HZ�j	����<�	$�5��/ o�>���Ht�;�Ӽ�a6��z�<]�V��'<���<�� <bU=�K������O������7=rȅ<>�!=>�:���;�y�7��<��]�]֣��V��v-=3�l=�	�������p��	(��t=?���	%��` ��׍<�L��'=��'���!�Ѐu=�.$��P�<��<+����ü�31�,Oͻ0���eF�	�<�}<<=j8=F$��>x}=]�-=�=�g�#Bּ�V=[eH=v�==���j�C�\(&;�r��D)���)�2�G�?M��߄��<�b-����;�q'���<��A� ���\<m�0�)$e=�j��]"�?߄��w���<I�=HS=���}���=1�J;�;�<��D<c$&<�yC�O�=��;Ag=�z?�]�*��[!���j=�9�ؑ �^��<��'p�<���<���<�U<�h\�N�%$��j5=�T�;�G,=� ���`�<X =��';Y�H�#�, W�d8V<uR�<����(�:Q;�<C�U<&%�̈́���溾`�<�z3��IѼ�W�<����g��<�[9=�n =9k=;
H��𩼏Q=(�P����;ϔ?=i2=e�+=7:,<)�}�s2;��#�N�:�U=ݙ+=����h��Ѧ;��r<�s#���c��&�0��<�i�<�M�R]0<��=�$I<��=[���}J��Fr=^���ΰ_=()O�Ȫ�=��=� �����ʎ<#A~�-���b��l=�%$�G?�n(�g듼VY,=���<vL<O�)�tf�<0�� �d�����AE���=���\�<����.=�Iq=���;��=`� =~�<�b*=m͂<�$F�1�w=��*=�~�B�,��� =߲9=�P<��js`=�↽<���v�.����;g�r=�& ����J�,���:��j���I=�D �Z� =��4�X��{%o�N���|�<1;��h��1�üں)�.m��}�1/-��&V�V8=�HW��K(�Zd��]���<J�D�=��Z=��;k�4�u��<3TH�[�;5�;�W`��J4=���L�I=c=���1�N�+����<���<���:�,��X�12�P�=p�9<�Դ<�����o�<	��}0�;ޣO�q{�����<a��<�a��)<�~���1��=��<a�g�*�F�5D�:C�]����/�T;������j��Э<�(��I�k�=�����r�0&�;�;��<�յ:]Zb�6�=o�<!=�<�d��<l=��<*8ۼ��C=	=�<k_=3�)�l��+�<���<j/^���?�'� �a����� gM=��=d�[��G?���=��=�uļ>P���(�<U���'�<S���eT�2���bB�<���f����<�] ���=�}����;���<	�A=3�\=z�H=�x<��t=��<��<����>^<�=c[n=�
6=ᦲ<`l���]=���:�"v�&�;f�Ҽ)@<=SE�<$I��cv-=He�<�U�;^��w�:�?=���<��%=��=��<���V���\
��S��zL����5е<S�
��>B��\��kɢ=(��<�a���2�Qu�SE�=E펺7#9=��м�<E��q�4=��<�Q�
XT<��3=��LL9#L�<�����)=@���K�;�ټH=ڻ�7�ԇ�<�ἇ�R=4f@<nҧ<�U5�����Y[�;x�b=���<�]=���F���;�j�a=]�<�����K�kUD=�]�;lNμ|΃���������a�;m}�?��<[m�%�<A�<pa�<�+�<,�˼���w̼�<�`��c�<]+�x@=�Rl��4O<(׃��.Z= Ma�jH=��8�_�G=!�5(=NRh=&Ԉ=Ү�<|�0��O�<KX=�=��;��� i�;�#s<��k=�9`<���;�h����(�V���;/ ;���o��)�<#?=L��<5JA=�4���B�<���:2�Q<��A�Y�2:|�*<#=��;�����l =X�g���E���M<��:�{N;2��<��¼�/��� =c��;����R��<���M��c�<�=�������<KH6=�]P=�@�<gjo�L-A�ɺ4=�i=k�;�<��r�<q���p��k~���<̨=�.�q=�m��6���0>ʼ_�G�N8��R�<��:l]��N�Y/ ��c,=�Q�<ﶡ<�g�6�B=�|��ߊ���<-�5�r�J<�%=qG���_W=@�<Z=$�~�d��d=�k�\��;Z�h<<�����:g=�V�;�@<ɚ�<��=�XO���)��6=��v51=�x�<�y=�c&��8���)�5A��;�ؼ��Q��[{�@м���Ok�<��8��
S�E��9-� =��μ?"=�4=��zoؼu�=���i�񼨬%�xS0���4��]c�lE�<e[<�[\=ty�d���?=�ڶ<��@=�F�U�����<��m<�lB=�b<=ˆT=�]ܻV�=2i�
`���h�<E[#��Y�<u��<"�]=@=�<8S=����<�$ɻ�����1�;�xP={-V=���<��{�����j��％el=6{�<��N=�J̻�]<v�'�Z:�<��K��!Ƽ�M�3��X��<}�=I5=Ѳ_<�~/�P�0��N���=�:8�LU��}$�t1�;���Z���Z�2�6<F2�6��E�X��q�<�����B��'�<�`�b�ŻG�=:k9����b�S�,Z��i<�IK=%�J��x�;+�Wx(=y��;�C=����>/_�^+=y��<��N�S�]=���<Z�8�=�;�Œ�'�==n�;�6����7����{jS����3A=V�x<��0��N�7(\�܎�S:�<>�-�����Tۂ����<ټN?�w�d=�0�<�.=���;8���U�=�6�:��UG�t>����ռ#���G��<^�u=�Ea��6U<����@��s�Ζ!�]9����:���%����#=������R��&�<ٞ�<�<3��4=f]�<��K��/�<ۑ����̼�<��	G=���<��F�=~꯺���;E�^<_'=/��;n��<O�i=��6=��D=�O<`-�&D0��J�<��
���]=ҝ�<�a滻�컊H<_�H��	[�l�:� ��������f���n:<�zּ�>=J"�<�x.=o�5�oP=~����D=��;����� h����_<UH���F�Z=xm���PO��uY��tf<ɜ�<�v�<i\a=�#=B`=~�;짼��L�Pf��I�%<�p�G�@vN��}#=3�]=�q�WU������$ʖ9�?��3=��I�yf���<a�U��q�<�r(��~)�5mN=��<l�<4�%&P=�]��gN=D'ּ�FW=!�Y=�d=�~<>rA:�^����$=�.�<��4=o�=]Ib=z����A�{���1��d�<|\�<���<��=vb'�� ��=��k���<go����<���<*9�=���;��<��� �Ή<�����d=x~<5��<}V%=��Ϲq�=&��;�n��	='k=�F�GA���,~� 1꼁<=x:�`�𻁓J=ڈs;m��z��;jɔ���w"�<�S���uC���<�&���y�AO8��w�<VF�ؚa���=OvP��n[�!
N�A�=�Y�;q<m����T���K=�b=�_�<K2?�6�!��^<��4<y�ļ�\�=�<�JQ���ü\�);Z�����d= ��SW��_B=jӁ��
��=�R=%���S�;�`�<Q�<�A=۹
=.� =j[=}���ߓ�t�!=Z�üU���
���K�ԛL�g�#<`r>=�B�X�_=e��<Q�2=k� ;;�=Zݪ<� �7�=YT1=�c=�>�XP8�dFi=�-,=�X�DO0���<�j��z�;n۽:�5I<v�j����?�<ְp�%�=��=�$<t��<i#2����6W=�we=(�T<��Ż�:��� ��?��hx=�r�<E�4<�C'<e���'�^e`=)�<p�&<$ϼn� �\:����V="��<�2�e�3=�%N���$`0;s�V��U=D0={,S�$=�(�HX<��<6�jrR=7@`</Eĺ�$�<ő=l酼V:D�I�ȼMu<�"�<;�>=Z�v�[W�
�4<a>=�2�t�=��u�*`}�P;��=p=��B���T=��<?P<�(w=jR=��%=&�=q���z�;��e=9(:<@\`�M?b=�"�<��_=?e�<e��ݼ~�R���<Å�<����q3�s�͘�s�>8�<�i��s޻l�l�YL�<"u�<��b=��|��(/=E���P@=G8�<��Һ�e=�%�<Dm��U༘�g�Kx��������<���͸�<c�E��zC���D��RT<��V=q%=���<�"V���<t}���_�<;�<AP���<�7w=����9�<ܮ�B�<�=S�<�I�r��;n�h<;0=���?���=I%=3м_B�g�<X����~=t�<
x#��/G�,�p�{�^q�<Sc=������<)H�<J��G8��y�}�==[�X<��c�Q2/�?I<O����6�FQ���-=�����#��`���v���ؼq��:?����疼����ۑ�>�����I�E�d��⻰�3�뷖: 8��L�<@��<9��([�<V��<"��;6p�{v�<�qC<e.<�9y�-��<ʒ=��<��^==�;<�¼Tm<s�R�V�;�<��1<x��;Y �O7H��큽:/�� ���(��pI�"q=<(�:�_D�1|�J�[=~^]����<Tx;P�D;5�����	����KD���w�;V=�����9p;b�;=�/<��1D���W=��y�QJ�L�2�(6�<���:���py�;<�7=�4�ȥ�<tu�=!��<�ɼN�k;~ZA<�+�<gHv<��=��=�X����<G�<������?�y���f����Z�=4�:=ߊ�=x����y=��i=,���=���:���<5L="�
=S���=,�ռ9D�;��^=��<^���$6�;�"=g�v<��<��};�<�Ab�-/9��F=6O3<g������Hk=��<C�5�i����H��?���	V=�ڼI3����\���3��p= v����"=�B�eǵ<R��Vڰ<w�.�_a0�Xs#=X9��'�<1F�6�ּH魼��=���<Ъ�{�<��R=M����=1-�]e;O�<(�U�&[�=��L��|�<�G��:�	f�7�4=We=R�e�����hrb��H<��K=��*�I��3���f�7����]��;c�һ`�>=[�2������%=�wq��5L=�v)=Id<�=^zS���)=�ּ�?<�?=>h ���<�&;͌H=�������<��7=eB�;'�<�$=y}�<���;�'V=R��<�ͼp�%<��ֻG��<��f���	<����r1=ћa�*��<8ؼ�%-��	��SG�c#.�,q%��^���C���f�+:���U�;V�]=�3=�n����<�&�;(�<�M'�]9�i���Ti=^p�<z,X=��E=�ϗ;��̼�j�<��<;"�;����9��<^:� �<Z�A<�<�0�9���ּɋ�:M���n�<�-�<ܲ^�mS)�+��.���;���;�M�<W�A�7\��,U����<�k4<q�M��� ��>^��.\=:@�6I9=�Ѽ�(=W�J��`�7.�7��<�V=��4��N���9=37�<wL�v�C�9<��?��["���;{��<���� <5���͘�/M<��<���;֙)���v}	����8P)_����	E����ļ��J=yHP�;}L������o�O6漃n&��S�<��g�"�=���<G���rO7<�"����A=�����X��:��|�<aS��B� �?��=�zO�������;c�s=�r�<�.D=�ռ�֎< �뼛�!�7Ww�����#(<h����;.}=������ǌ༓Mh;j�T�G�B,<�:j��,;�h�g=�;��<r�V=�O��j��#��]+�J��<��<��?;�c<1�<�Lc��
o:�TY=���;)�=��;�%D=ÉT=��=�~�����?*����<D�|=��-=��G�gNۼ*�{�1\r=א[=�w8<yD��{�<#��<#�-<�?7=SO=��=��?�E�=�A#�����Q���&@=;�MȄ�蚜�.�gI=�p�q���(�Z�H���7��x�<oL�o}=�k$�]?#=�V*����c���[A=�a8��Lf�I��<���<~{"<zM=��g=�Z�<�rm�JY;���\���`=�=��`��-S=��&=�N���I�<8��(�����D<W�<Ѻ�lk-���<|[�=F�X���a�j�,����ݕͼ�����>����T=Y����7����+�]=
���VR�ދ��*�<	L��@<R<e�����v�=]g=��+=4�����9JH�9��e=��1=�/μsN=tq��$���V���Z;ݐ��&+��h�\=VM<vDF��.��˼-0鼕�!;��=�h8=���6fʼD'q���7�8�.=���;j�;@Gd�%��<뜁����w�� l�<H0Ӽ֬�<�Y=���<�N*=4$=G�� .+=�YD=q =����rG"<̀8��LJ=�~��u�˼#��;�B��=�A&���	<I- �դ���$=)S=R(;r�r<@2��]0=��<J���-=sD�nF��W(d=΍�;����Fd0�q����D;8T�<hl=��T�}���w��'�:���s���W�Ƿ5=1�;�m;:��b����A=���;Y}Q=Lv$=��	���!���4������M=��8=��6� ��K���=��:G�y=��`����>��Ԯ'=��;��Z����<z�<�y
;��<�U�6=���<N1,����A�b<�0�J8?= �=�S���=:B9�+�=�[(;?7!;��9�4p1�\�c��\���h=.���:E�;>�����G��D(��Xo=�IG=Θ����'� 5!�R�=��=�c��0�⒑��g>�Sb<S��<�`=�,�<ZSh�>@[���<��к^o=:��<Eꑻ3�o�}�<mk��)�.=��J=A����=z�-=���(U=W"C;�F<�:v�e{k=��<F=0�=�J=il�<���/=�FG����<\Y��'�<=��<��<�����.���9)=�<�;x=�9�c=o��;�:a=�=�r�����W�=��;=P�7��8������%<����L�m�<(uz;s@<8�"�dI��>8=,H'�2d��5�g<��¼ɵ%<2F5=���<���n7�Z�<�' =_qH��2���-�g�<_8H=?����x8��d�.Y���Av:\���釽1h$< !=�=0��:N�7<�^���|~=/��<(N����<f�M<)�<[�{=$6̻���<�uL=L��g<W/6���C�cۼ��t=R,��=��'�Hb�~���:���O�~��ŗ�뾛<������=��\=Ml�< kU��K�<��)=I������C��r˻Fk=��(�m�<A��5&S=�2<�D켪�/��c�<��ʼ� ʼ� =>3-��%�<�����M$��Y��� =��'=Tw�<��D=�y<}<C�<J躻�[�<z��;|�4������;���AD��q=ڛl=������<#��<�D�m/?=nZ༘�ʻA8�/�*� �B��0��DI�[+=�n������b=�g��u(�������=�A= �#�:o޲���I�<�K�4 =vq���:���n<*�	</�����M��������2�`Gf�`�D=o��7I0�vʴ<T,����<ˠ=I໓��<U�<�i=!.d:o�x�b�ʼl�8�9>B=��w=��E=Nuu<I�<�Ib	=&�)=��	��LY;w=ِ'=���l)T=�O�<~�1<^����<EѠ<д�<u��V�;p_��8<��D=�� �&�}>]=�%�<q��[
=�^��ڼs��<1"`�>�D=�uW�:~m�S��<���i7�ŅC�P"�i <\c9=���f\=Я�<�[����S���<e��<�ϭ<7�/<��^����J*=��
�%�Ѻ@׼���a�A쇼�:��kxO=�����<uC�:�_J;E=�9<q"�<�o�<[�A�a=�8=��)=�xx�C�3=Q��<���<���������T���3�Ϩ`��Lܼ/� �Fg��"�%���j�<~������<�5K�}�<��l� �=/J��t�Y=�TN=��<	�n=�-�ՈI�
y�<�F�Z�<H�I�ImZ���<�X0�Hx���H6�;�\Ｘ�#�e�~=Z;��1I<��;f^s;~�.<I���.<WE�$��<��3<(�t��/z=���<�:;�_%= }�21f=�_�=�l��ƻ�S�<�~g�4pL���s�l��<�Py�d�<M\,=���;K��=�z<N�r=x}^���2��G����;d`V=�K3<J���B<�b�m�~��	����,�S=��'�d�=
�]�I'��,)���=2�u=�镼�?=<��W�=�+��<��h<�ԅ��&?�W{�aF�<����A?<+�/��<���^Ƽ*.=V5�X��;1^�'���߻ԾT�̲�<��)�0=|C/<��=z�2<�W
��mE=�Fo;Y�v<�w6=/$���y�U=lTj��<5?�<ʸ����N�!b�~"=���<�4�<K�5=q�Q=='M=4�=S=xX\�j!f�������;3�{��I��7F=��u�<[�N��>P=��I=�vI�*�$=�~.= b>�Ąs�,'�;��<�����Z<��;d=A=I)�<x��r@��Yq��:�<0e�J�<z��<l�^�N�ȼK�\��c�<�+)�I���
��N�<!��1=�Ĥ<A%��Pۼ6��wx=[I���-�<�=��5���Y��u��D�/~��E=��^���g=�R6<|�J=ȣ=ǫ�=��*����F��<������%��-Z�5%<��d�̵Y<�r��$�=7�={{=�9)�!�H=���6<T�L=m<���;�54=B�2=�}��}m���k=�ټ��<fU�<*����<Q��3|G��a@=N�B=�a�;�A=d(���=&�9�ջ�z=H��<_��<2/=�Kټ����ˈ<O��r;��2=�X;�={�<d�	=袮<K�=������+<ieY=���;B =��%<�:;�{���Q��W=:�P=wGE=�`C<�̎;����9ݻŦ��*�<H�����M��:=Ȃ��vi=��<�@����b~:�7R�^�<��!=Ϧ�<�?=�N�b/ۻ�~B���Y=�6 ����<SZD�b[H��� �I��<fꢼ�<��W=���qꪼ�F�=%,��V���<e`=�U%<��^�5�<�ׂ<c-U<٩�T�=ߊu���X��B=��=`�<�vА��u����DT�������0=��3<8�d<"r�zo������=3��h׼�O=Ƴ9<j��ҋW=�n`���)��/=�ܼS�\��k>�K#�`?^���==�ߎ�m�ͼ�~�<��<)�<n3��ajX�N�4<t#-�_]!�#F\=�'L=��=��|=@/=��.=~.�B�=UB�=����/�1����Y
ż�nL��z�<�-]=�����K���H�=+8;�Э;�?�<	��#<. @=�)=j�3��s�<cG=�)s=e�e=R�<&�C��t=8�������<[�=�l����=$E�'n�;<&<d\a<�M�� �Ӑ\=
�p<��v=t^���=�X$���f7U��<�u=x߱<��q<L��<v,=��<0�K;{�+�nUf�g�!<�p=1ü�_�9�p�=/ �<x��;Sp=��q=`��_O���2��>�<de�Xm=;�4=��5����&hA<z\!=�Kq=��<ߟj�pq������h=dt���ļ�����i�<&Ļ�<=�6$=pp�<UF8�#���.�����~�ۼ�<������ZO=���<dp_=��%=�LV�Ԏ<�6���$=x�d�Q�;��	=:vz<Iy�;��}�U�#=lS���W�:�8�<�/����<��g<�����.�=T7<�k�=�9d��vH� �ּ4tüޅ�;�ź��=A}�<�C=��=�g���h��	���<�_׼���<�b���y=��I=�T&�sSM<�78���>�~�=�B�r7��x@�V�q��U=�BѼ�2�<΂�F$L=�8�<	���=vW�^bQ=�H���;�Kg��Ih���G�<�đ��]�;2��dql���<W�q=r�<Uh8�����N��X��<��\�jo<��=Ob�<��<#7;!��u�5<R�v=����F�;#*=d�X�`t��MX�
i��9�ڻr�^��^=&�+�o�<�d��2���d=��_�K3R��@�:�C=���<��Ε^� F,=��?='�� -��4=��=�4!=� =��0�s�<���W<�
��`+�n��l�o;��i=��G��
i=dV5��J���G�I犼DQS=/l���S���������
�4������
=P�U=��z;c��<��*=C�=k&=qk�<=�<��(�F\q<.]i=X�/=	L�q���:<��<E:�R#�{�E�y6=n�=<Q�����<M�><yCջ�iż�#�<��	����<vb.��2�<^*d�Pl�"=��-˪���;�!���1;hZ�*�Q=�L�;-�$�9�|�!��<�)��.C
=:��|(��D+=��=ܹ�;�Q{<���;l��'�<W�p<�4=���<���<*>=y޼�zҼ�rj��V<�j��	�]�;�[���<��=�	C�;�9=�s)<x�<���jn	;�P�=L�C���@=���<�]��G�5���<���D�=� =�V�<Cs�����r�D�F'q����;������l��/=#+�h�$=u�;��g�R�;�P��TU�(��<�I6���<��i��A==;�<M�ӻ	h��l��򜻜��=_&�;�n����<}#�<�T`=�
�<a�t���=q}�<��߼�7G=��<=}<��Q�<�1s<.<:�<@�=a�H�xBC=�q��JK;�B(<�e�9�.�*8����<�F�D�����PC=d��9�D�M��/��6ȼ�
=��=�}-�>�$=
��� ��{�_���<Ϸ>��=�֮:�1��F��ԝ;k�l<�ޥ��C]�,g��|!�$��<Tg�<:5]=�l�=f5���r.�(m�<e{�<l��7͆<�<�{��?=�$'�9'=�Gu��D=��h�J9�<�ɢ�\	�<�;"�N��a�����PhO=v��<�3�;s�	=�I=_K�s~�=�?�<��ļ���<��<������;��Ȼ����;!D�O�I=��ͼ׈;�X�<j�3=m/8�'h
���E�XQ�kb�nD����<�=�缥y_<ܸ�<7�<7�<���<�K`=.푻�N�<�7���¼�@��[=P�����<,�e�&���|���������*��ᑻ"�����R��м��+>=����:�-�����Q=��<P3]�ߑ輻r;
{�:� �:�lҼ���`'���=^��;ݛ@=4̰:RY����p=,�G=,t�MQ=��m<c� �X�=Q�-Q�<r��c��[s�������Ҽ.�<cmR��iK��P���A=2��<�ƾ<�v���<J�J�e������.��%�?B�QV==�<X+��4�<�j8=�'�<w��<�(�d�^<�~�F=7l<7���'s��A���/�3<5Dȼ5�/=�U�ԓL<��< � ��廉`�ݽ=���<��<����; �:���T�	��/���	��T$�*ᒼ�����Ӽ��b�z
<�5Ҽ�����B=�2-���y�DV%�GT�<) <��|<6�)��	��Ϲ6��Kq~�v�;����<K���;	����!^��I�;����o�d�U{�'�}����z<=�xc�Y����/O��N�:��<n�Ӻ�	����<�Ip=�Y�CJ=�ռ<��xN�U�����X=3&��XG�{r]�ή�<n�9=��<) �ʬX<7ᙺ��D=���)T)<��Z��^h��󔼉x�xi��v�F�=~Q�<DZ=�<S�;�/��祼���<���<��!�*ᗽ������4���<��&��R<��9�D�Ҽ���<#�=��</%=�rD�E׎���;���<^\�����k#�<w_ <D�<�]*=��<jax���f=��#�#�<��d�;�n<=Q84�9�`�{4=�s5��!�;B�(���#�� �䌼��D�'����*=��t������<v���I��3�<Ds�<�ȼ�������֊;l#��c�=�<?މ�Ş!=LuK������d=�3=u�/��-7�s� =�{��V�*=V��oˁ���f<��<��`<'%���(���;��<=���<�j���9I<9��xhQ=��\�2Y=�C;����W%��E�	R=��p����^�<�G�;��������v<�y�<�¼��p�;��=B<4=	2`=\�ͼ�=ӡR=78�)�<�j*��ܕ�����=�β<��)�L�������9��N%5�����4=��<��/��M�<-r�=�e=i/A����w��<1^��)���;��{=1ݯ��
H����<�=1S�U��;	�<X��mQ��97v=�+��B�wd�:Y�=G�=t,V=Tv��ʼK�Z���E�׼�B޼-��o��:�;=���ڻ޵�<�ZH���D<`d=�j�<-^�<�
F=G�8=`Z���D���7��v|<T�`�tM<.�L;	�����}�j�n�
 =9W��i����;�||;�z�=d���d��ߓ�x�<4¼9�a�������\�<b�2=E�h�>d�=����UҼL��<<��o8>�\Xͼ��s�m��<�V=ž/=Wb3=�\�֌<`�\���X=J{'<�)�?|=��=�_=,ֻg`=c�(=E��=�?��d��<|�9�A��</2.�ڔ*<9�+<��=Js�Έ=j�ȼ�g=hZ�;D�s��ɂ<!G�خW=L�C=���<b�<e���]=��׼>c�<N���:��fa!���Q�u	��0^A=� {=�ɾ��<Գ<knb=�7<z	�<6���@�X�~�[��=JZ_=S�P����+`��jǼr��<j>�<|��NB8�=)~�2fp;)��<��;��	�i9��_Z=�FԼ�'=Ŗ�<FK�:+�,�s=�%��A�v�ܦ0=��$�3��<LϮ<�c�<��ƹ�H����w���=�pMN�B���,-�f�S��j=ӏ뼾�b��l�<G�����S�X�_��;����6=���e�U����<��=�g0;�N[�ՠ�=@t<��r
;Ȁ�=6h�����vü9�μe={�5=�s���������	=6Ln�_��;���S3�a���Ζ=!�+=B�<FA�;�폽:���4�y=0�;��6KK=u1=;��;o�==�n;����u�����Y�Z�6����ܢ<v�t=1�=6WE=��=�8n=s�!����< T�<h��<e�<�:,=��Q=e��<!C�����6(�<aQ�<�w
;UEl=��ϼ��_�9P�;�!��ȻB�7���O=𵋼h�><��i��޻�
�e\F�Xr;���7琖��cA��d�Q�p����<�6;NO�<Z����1�<�"�<d��g��m"=�f����=�,�1۬�TY=^��	=��=C� <:΁�2H=��<�o���%L��6�=��|�Ӏ�Q�<d:����ռ�!8=�tL=Z2'=���;���<��0=��9�+�<�eʺ�c/�&�,=�!=Ƈ4�ok;I9<��l���c=g?W=�R;��<="�<�4Q�x��n;ʼ�b�@�W��^�껈�,��X��l<c���,����;��ڼ�*}��ø��07��j%=u_�<�<�|	�5�=��2�	�,��%���� <~��<cS_�P�w�N=�)�|u�����~g�]�׻���_�#=��R�>�Sf�<��<#H��0��L<��Q%=zr;��s��<-�<�p��q�?=���b�o��]�i�Jh\=��b;9ه=�%u��o����<d�P��(��}�����;�RO=�8(��<���z��=��<�;���1=�se�w�M=�`ʼ�9�|�8���=��={ ;�x.5<C�.<�<<�_=��;���<�]=�#<�C�;<R�G��s�<���(׼�X4����<)iT�⚻3K>=1`S=������y�6Ղ<�:g<��K=����m;�z�<��x2��ƭ�]�w��%���h=��=�4)<4��<��W򅽮�<H�j������޺Kd=Ya
=6��<�=�\�=�(s=��w<�o5��ڻ�w<@�<���c�=���=D_S�n�����1`=2���������<�F�;7�L:��=5.�I�;�2�<0��ۥ/=������	�;`=C��<o��骎<��x�#�2=��<@���̋��U�=̲<��I$^=�� �?=���<��̼m�n�(S-����<�X��i�<�J�<EY<��=�R�;�0=��W=�Ma��<�я�M#}<�̰�@�"�?�<BÇ��t�;��G�Q)=�yu�C��<��}�J�<�'+=õD�d=F̩���7=:D�<� ���=��r9�|�<.^���EҼ5i4�'�5=KI�:q��;Y�<��%��l�<?n\<��5<�;\U==*��<:M�I	�<�m˼,@�<���jCe;�$�i˫�P��<k�μ�
=�@ٻ��\���:�#;�HN={ Y��L=K�=\�|���Q=V�-<�֤;쌅�_v�< \���ql=T����z�,-'=	fc=�\���Ed�C�=�s��XBL<�{�^�X=�c�Go,<�պg� =��;<�)<�S��|;!�\���K=i_<�h�;��6<��/��ż^f༢���������W�;ݯǼU��mu輄�U=��M�~a'��3�;��<�vl:=�����<��N<d�ǣ�<�i=8����<Э�<�Y<(��<Ss��$����n<!�YJܼw�G<�a��
p=�/ܼ��=�Cg<�����<������z�/=lŒ�2�R�=�ǼG�<=:�����S��;�:�7=x�-=�G=�<�	�<�-�;C:���D=id޼(3p=ƑY�����#;���U<��=��c�T�<��<b�9S�?="Tc=�1!�K��<%?�W�:;�L=s�k�
�,="�=�����_b;f�����.<�8��`�*6<ZPD=y�+���/�f[7��d=�����`����X=�m�<��=ׄ|���0;3-�<��;��2�<�4;�mQ=�;|���n<ru�<�H�`���<��Ƌ;zw��̒X��_���)=��n�����ˍ=m�[;@��Q<�F ��1=�`�< L;��<�5�<�����μ�gK;r�{�t���r���ؼ"`�%���8~�INh���=1��<�:
��~��]B�h��<�_*=��U�4?S��K �����b��I=SC���oH�6��;��<������I=�=̼Tg=��F�e��<�8�<�+<=�O��4��Ij�i�=�=��=�<�����ׅ=�仁�e=�^==���Ľ�>^=�\����?<:r��8��:ͱ�1���LlC;Gj�<�;i=�h=n��<� ��w%�c?�;�<V��<�X7� 6�<V�=IZ��.Q��#9��=9�=��἗N{�]�#<�}0��=�><go]�8�*���;k��<~xk<,G�Uh=])=)��;Y{�<���~�d���u<M;�<���h�����x<�L=S[�����v�9;)~+�.�a=�;��J��oJ=n���UaI��x<��)<��=!Y��Q�<t��<CZ�<��R��&%=�T�<ed�<$7=����1Us<��U=�P�<��j=�dI�yz��1�a=|l�[׋�X�c�������X����4_=}��<K�H��LлR3&��=+N��	ڼ�5�<�(q�y�K��/ �����`����Ƽ�1�u}V�Ѡ��X�;;®��R�@<��<���<'Um�#9ټ�O3<ϼ`��/=�/�<�摼��c���<�-=#ݐ��{=+E0<��=�?
���=x����G^=ޗ>=��7=���=��=)1��懼T{׼�3����<T�n=D��<P���u�K�+�-=�==R�<,j=���<�{n�'�L=`�l�{f軛w�<�G]�²$��l�<�;����MP�<h)���1��\�R��ho=~�R=�vd=�,�����t=}>6��|�<P�N�A*�<��G<>�غ
3�<ɨ��x��<X�=�ɼ�G=*=��|=��<�#�;����ü/�!<z��aFH=a;c=>촻�n��o��<n�M��IM=�L�<�ܝ�i녽�o=�ۙ<����5�<N�<R�9���=�=<��<Ne��!�$�a<E�$<�y��<|(��g�缂��;�ᓼ�=�v<��<�';>�=x9�����s�<���,�<�z���=�1�<*D=�y=:#����O�_5��AP,�v�&=ە�<��]���<;t�=��b<��4=.!�<�x<I���S��x=:�<�+=��<��;�$���7<�/	����<�S";�3����TZR�l�<0l@���'�។�b�<v@8=YZ<k�ݼ�QS=���b�>��b�<�n�<%Y1�ɁB7�G;|�㼟Z��b��w|���d+=���<h��<�#��#j=>H:=\I�=C.�)(����
f=�	=(�=?�G��\h=Z��<;V�.����Լ{�����<������<�	�<�n6;O�ͼ{��}�<h�;u�=[�0=-rR�x�;;�k�x��<�p+��,@��h=�»��M�ZUq;"q=x�<W+<VF=P==�gF��=м�7b���<v�:G��<;�<>�p=�
%��L�<��ߵ�����D��<��:����O:=`t�<!�<�F�%輙�0���'=�^=Ҽ=�X���3��*=��;�3[3���c<l?<��3���=�>;fgG�Û�<�e=�VO=��K�5�����e=�5�<�e��E==1vZ��x=���>4#=jV�<߮�h���i/�R!p=6�I�]�I�������
C0�e"��+==�yP;���$6��̳</lM=��K=醼��<��w<�v�< �꼾ϼ��<
�)<*�=dBe��Mt�M?��M�<�N���l<��';�!�;"A!�;�V=��'��(�9y�Ѽ�ސ���n�˹�:T�\r໅`s<uv_���e<޺F=�b��*�2/{;���;�'=��P���4���l<��:ã���
�hЙ<��=ݼؼ6@��jB���<�� �LD=B.=��]�໴�X=�ic=7�{<�~���h=	�<};�<�/��z4=��=I;C=��D�J��D��<����&�G=ʵ���S��U
=fi�0ӌ;s\I��L=��s=����&=�Y<�17=�%w<H�J��_�<�X<�h=V��Z�<��(��'=���<�M��@Z��a�G�2�>�9n==	��|mܼ���.�P<֖Ѽ<�L=�Ǚ=w�ռa�����49�tP��s�<l;�M�ۼ�����'=}G=�m�=I*<��;,(A�	ҽ<FL���y<�)�:�P=<V\!�h���X���Un��ߍ�.��<�>\��P��;0�J,%=�#=��Q�-Y����</�����<�Y]=]�< GW=�n~=9�=��<U�=ԛj<��$�I�_��M=+�<�� �	OL�č�< �<^��;��2=��I=d�<x�)��i�$}�<֔=��<�*O�� \;��<
�=�����V<�8��(��U�ӼV�<L��Df=�h4���-�d�J�Y=����-~J�8�N<��/�J�ʼ��^�hᗼi�[<�����<���s+=Y��<'De<C��;��<��9��0W=5B���<��o��5O��z�<v�<GL��R��<y���ҵ;��O�w����N����Db�</H<���<��f��<20�K�:�O��϶<�Q5=�RN�Z92�'�8=��D�vGc����='���������2��k=��ݼ���ɼ����V4=4�<<�k����ɓY;Q��J�J;$
ٺL�<7�;�c<F���9���$5�;�1=�Ş��t�c�C�k�:��<kwq=�[�;�ź�湼Dʻ��-�;���<w�=��0=��%� �<����Oo���p���걼�^=�R����*�o��;�J=()�<��<��=�(���o=��5=[e��$�7[=�T���6=�Q�g9=������<~=�	��w�G ����<f=i2׺)�S=Qۺ�O���<c$<'�(��pJ�k���t�g��*j=_0�����<�F�EՄ�R����.j�m�O=V\ȼQ�S=�Ѐ�L��<��*=��D=�vJ=��l=b�Z������X���@����¡�ŗP;�����\��0�<<�]��2=R<�����P�"�W���ټ�Y#��=GT<�~G<�1��T��<Yg
�.��u.�l����;R�<�d����d���ͼA�^<h|5��=����z�<��\=3;1��:j���D�(,�H�b=d�;�q̼�[�-"'=�-=U?��	�+�A��<���<!c<��gl�# �|��l�<�N�<)��=�Ҽ�c�:��<�����=2؞�MbL�|�E<�s]X�(�=�S��L��~,<�(=kٸ�+a�>I#=~�:&�޺�n���9�sLM�_5=��,=P#U��X=W��<s�=V�.����<��<�*P��b�ն,<����=f� �p��=2��o�A��^=���<`�MbһM�6=F��c��Myd=�v&�Τ���t���珼�P4<)�T<�*���G=�X`�ȼ<�ʒ��o��^5��]A�m����!=��K��l-�R;.#C<0We;���<Xdy;��<O&��m�E�g����ʼ�'=6�;\�=W�u=ˌ�<^m��r�OD=3�<_Y�A�9�=?�c����(=K�	=���<�-ȼ��<�����=w�<��;�( �d[��n<�; (�ߌF=W	X�����<�E�e땼�aH=ۭ �f�a<j1=x~���B��0=*T��E��<е���\j==@<ad=�-=@ڨ<S�<F�ܻS�J=�]��;��zz�.�����E�8�w=�F�<��D<u���=���bD�r<<$��<sJ�n�0�=��<E]'=�#[�Ԣ>��z�vU�:Cl��,S�ߟ����<�?<=E��}���I�l=�Ϻrr=GX�<�v��1�m=���<�8��8�<eP=�cV=�R<���;=���7=��=x�1=���J��[/:�>=P�����:��p=�pR�|ۿ��瓽NZ6=ju�<&�<U���/�<�u<P���m����4=͋I�%�1�������}<���<K@=�s=�+＄�]���漌�J��\ɼ6�C�U�_=�����&�Y����<���<��=��5<��5=ɹ	��|�QO�<���to�<����=�v=f=�n2==*�H_Y=��!=��t�GL=¿��!�:P�=�RN<�M����=�H�<�!=�aq=�,@�����6��X6�`*5=R�E�VLἺk=t�<i�%=ZZ�;�z�ةj���ܻE����%=?D�<׬��t�����9��q;N��AL-=�w+���D=B�z�`;7=����<+�1�}I���D�<�k����<�n<�LB=�f�<T޲�-:�#�X��<�Dz�V�!<2~�(^��Zg=:C=��=��"�e7+�2c��d=�<�:c;@ڽ<��28�<O/=�IT=�id��Z<M�=��4=��=���<XZ'������Q=π|���<��7��[��(��<��<a"�<�%=#��9X�:��0=��{<+=+:w=�����R];��<�w����?�Asi=D|ܼq�j=��9=��Z��-b����4<~�+��x
<������ =��G��<��2���ͼT�_=��]��-2=}*j=��8��ۿ��Њ�/ź�	����=�%�<	���Z߼�R����d=5s���c<!�Yn=�MW���^�́=�7 =�l�5�.=��J�3�Ǽ���Y(=�����������E=,Mz�p���b"�o��<h���='ǐ<�!=D7t����<{��<�SL=[�<��<�O=<|��U�d=B���:�=5��<���<�������<U�<��f<�;t�<���<�e�@`D:ʮ��4I�WXl�CV"�$%���..���m��	)�< ���PJ9�PZ+;&۲���u�M��.=A*:=�F_���
=��<j.��~`=~�7=��=;!+=��G=�z���6:�h�=T��9���#�s��<��X�`?��Z=c�ټ��˼�$�;e�&=aW��F��?=�����4=�V)����<,HB�:�N;j30�\Td��m7=X�&����<��<x�<FJ+;�<�=��A�W����<���<�w��<�����Y{<8��<�/<��U;<�;�bm�-3t=L�\���� ��f�9	��=���>�)=EG^�	[T��ῼ�t=�ͤ�0
�q����e������R����-=�P�<�H���}<A��<t�V=�:WM�F�=cNp�`;j�Z7�e
��~Qx���ѺH�6��ͺ�ɻ�%��}E���:��պՕ�������:�>p��T�B<U��<]��<�s�;0�|��<P<�hD�O�<V���2 R=g=l=��9<�$H�!G=�/}��tB���?�n�Zg���y���7=f�>��Y�<xy��ļkϭ;$��"P�Ȩ6=��]�h�ӱ=���H=ѳ��S��	|�<j�?遻��==1�*=�O=����#�:!i�Q=���WO=�yҼJ��<������!=��<^�Ҽ��;5�B����<5 g=�E
=�9=��=��W��O�a�K��*>�� z=;�t������.=2�7��.V;�t@��2��jv�1��<e�~�,X���\��^֡�O<!=�j=dj=�;��e ���N���	��hr�r��;��>=2�P��X&=��[=�a�;D�0<�\�-�"�4�C�*#=��<�X:���<��5=R9>;�96�C *��y=�U��;�3=��g<TF޼~��"I��Ԁ<����goO=�۝���J=��ɼ�B_=q��i:���_=?�2=T�=���� V=�\�<q*Y�@�e�y�=�o�K=*�D��}1�:��P��|������BT^=�(e=PS�;YNP=��ٻ�&=�@�<ϳ=��<)�&<�(�����<��*<y��=�p;dY���
��#=7�	=��=�D=S�)<��=�Sx=�%�;��J��=�
�<��0<R�$�g��<^�8�o}=}KH����<��܃�<2ۼ��Q=�B�<I9.�u�`��F������5=2\�8ɼ���<��<�a�ʼ��r7=���<T��<%���Ks��|\�I�F=��"�;JB��]�<`�4�j����<��;�A2=��p����_��<94Q=t��l]6�E.���}�<�7<o!=�aw��8�����j��S*%�E�"=�_���<���N�l<X�9=R�4=X% =���<G�<�����~����B���<R�Һ� ��c����?=��4=��==]_�<۝ͼK�r����r���1���A?=Č <{��<A3�;<ϔ<	�H�%WG��WH������<�L���:�j��勸<�TQ=΀P���<$��:�ST<A�ؼѱz����<���<CQh<9Ӽ~��</Q�<�5j\;Z�ͻ��;�R=�U`=p^=t�,<]�-�Ѩӻ#�<��3�Y��ȡ��9��<���_Ѽ�a%���<(�V��Y=�'=���<%'�;�V����<��;���<.nE<y�X����O�=��p��:�<��4��bc�F{g�(10���~;V@�<�輧��<�Y�Z���l�<+�r�q�Y���<,#<��»��8��SR�G�Z���h(��Jb=��H�#]c���c=��.=Ao%=:k.=Ѭf=/�1=N7S=��ʆ=,#z=Y
k<�F=i5�<�Iȼ��.�?zw����;��0=;?���]��}�������`=4W=i�����?�..�<�Q	=�J=��f<���u�:��J�U�{<\���_ʼ~)ͼ�C���Ϻ�bM=#	�ղ�<�}�<�ȼ7B<C�<����}<Ą<��g�/��<$0=���:[C<8ܨ���8=�cW=M�9��@w����=���;���=
˼�[=L�x=��=���1��;Z��:_��<6w,=,1Z=�`�����L�?��:���*=OR=��\=�l����;��<�r�;.��<F/=n�u<�ʼ�<���<+�P��W7=��<�#��l���
e��A�<+pm��B5�Y�'��T=���N�<��ռv��4����.=�x�=,��Y�<U�"����<�X�<��<��!�C�;���<EĘ<�2f<̹Z=�
1;�==V?�<���;�μ/��<O�A=z\A<ʟq=D�=!�G��Bh����; �6=��;=#�Ƽ��0�_�����<ۇ��M�;�	�'���b=�Py�����d�F=!��;=b^�����������v���=[5��
�%��<��4=N�<"L�����鵁=,�5��8)=� ˼I�=��=��4=�0�uSC����H�D�(g;����<p�r<u$=mm���s!�w���;�.=�	<2�t�z���2�=Wqe=�=e�x<c�U<*b=��L�m|T=,�`=���0!�<G���FH�?�ʼ��=1<�<jP7��{�����7;��׼�1�&C[���;z5=	2�<�8 �c�Լ�������;�ͼK�S���=�s<74�<�/=�v<m����ň<�� �s=�i�0{Ѽ��R<��<�B<��y�m�;ޑ�<%��MI=6䑼6N�<lL⼃���-h��F|�<o�<�N	; ��I�I���Ƽ�d[�~�e=�=�}%�w%��[�;֑O=ԜM�2(e=�O�<�Ij���<�z=��6�Z=��A=�YؼK\R=��(�{���W����q<����r=+K����<�I���'���P�I@�<m�0��	7��A=?Yk��{��@���ט��n���=�r�t��{s=\�<��ûO�⼸����^=5Ҽ�]μKgV�բ7�ޫ�<ȓ=��&<���:�<��!�?=�}���)�4/�GH�<5H6��Y=f$����t�� E�י��Cʎ�$�Y���ټ���w�,=�z<m?_=<�a��RɼΎ�<$�}��}�<�X=B��:�6<3,I=R`�;ZO
=��V=����<o�d:c��5	=�$=V3t=�9=l �F�j��P<�Z�Lh<�D�<.	&�]����%���0�SY;��=��U����T�����/Cm=O8H<.Ҽ/[R����:���<,n,=0��<�}=���< �<)#�<9R�<0E =M5=eu<lļ���=�,�t��(f<��<=�8�����3=�J5<q�[�Y�<5��t3O�Ґa=<�<���iM0�9k0��k�<�>���]�!��ˇ=4�f<����x=�5��_M<k��<��b=�L���Q�+a5�����L|= %�;hO�~ց<G��;�o<uIn�(UT��6��,�=[Y�<'��<�=�K��b=���_"ڼ��l=n�<�[;W�Hs[���<xe�(�"<=ysټ�'X�T�A=����g�+=\f<��{<�4
���=��g=W9����<j*����<=u�<�!=ȊD�Hf%<}�@=Oet�/D;��G=��$�CT;h@���<�|��Q��g=X�U��2���0=�wX�?��<���<*=���;yA��>�u��Ǽ�z"�ŵY<F�U=z���L�N�=���<U}����˼O�<Z�=��<_�?���=B�I�`��`<�x;=��=ɪ<S2=>5S<;��c��,(T=��:��c�<������F <�	�ϼ�:	�f��=��v�,�/=}K=��j��\!=�٠<���<�]0=;�[=�O!=μ<ZQ�,�ۻ�f���:�H;A��<0�<m��q�$=�c�a�=�1'=k�k�w�W=]q ���B��� =KȺj'�<���<�7y��?6��- ����;O�;=F׼��;�V!��Q�Uu	��q-�R�$<>��<Oy�:��=G�O���w<Ύ�<�<,�,�-=l��<W��y=��X��M<m�<o9<���<&�8�	�����<0��WQh�Qɉ:�&=go�<�X<����W�.#s���p���7�Kxh<&A(�p�;8t�;��>=�ؙ=�� �ph0=�Z<Ǵ��V�<ZH=�'���):G�5�'V2��}�<�0��c�{;ˁ��)-<��M=��A���?���h</S���(�������m�$�=����[q��7����K}a�T��;���TM��)�K<�-�8ؼP2P��#;����$z?��0�<���<Z45�X������<����e��lJ�F&���ف�~�=�g=lŅ�$�ͼ�=��ݼ;�%<6Z=kF���?��k������<��;�� �c�t=u'��q�=�F����<:n<�i=_h�SKz�m���;*��fu<O���3q�(�i�hZ�.L<��g=�;�<rS�U����;6=��'<fم<s.�<�<��b�z =4�,=�/=3(m��V�C�>�pC���2<�A�<<�]�@Z;��=jbJ=�$=�)�&�S���������D<�w=UC�w�=��]=�Tb��� ���;5<5���B=.�J���ϼ?�=%!���?B�~��<��C=
k��%Y�Eyn=�`G<�~�<���Q���!��S�i��:�~T��ո�$�h7r@:�]�q�Z�.=���<�k���=��G�E-�?;ʨ#<6[z=�vX<�:���O��'?�(��;%o^�2��<�g�;<[=ViҼE�M=�_�Y�0=�;�I��M�6�R6�<N�I�8� ��<zzZ<}A�:ߢ2��2=��+����¼X�X��;�r�<�P=
\<}h`=�-k�ǽ=ϝ���K���=/��<kV��d�v=��PUO<�}�d����7��"�uMi=5�96�{��Q0<�4ɼ� $�@W�<�9�����<�ތ<�+�6l=("k�H�<��4�Y+���p��d��<=�F����<l�}���:M�1=�hQ����<y�<�/�q����-=�+��Jɡ;m~�<�	n;d�<�x=��H���p=�U=�Rʼ��uQ���g<r[��I�:?{]=��v=t�<S��<;�Ǽ&{6=�O<��u���̍<�.=hV�<?T=��=%��<�D:��j��jc���{���<��<�ɯ;C]�<yr��OL��<�<�m=.�6��<l�<s����=��ú"�L��kE=���;�<��߻�0=��=�$�m=��L]=��B=w	2;�7��9Y���^�q����+��$����M<~P;�N:��!��=pÖ��*6=u�:N��n�<=���;�b�<��E=u��=c)�<��t��7<�Gr�x��g�=��L=�o)�ci�<d3i=��H;N����4�^��@�<�n��v���F:<������&���Sx�=ἄ�C�?� i�<����b?=��g=BC����<���@�&��sF��f�"G��==;�;��#<�C=�!=�	���:���e<]�ɼN�<\�L���#<!%��_qk���:�~hJ=�A[<����	�JY�=��<�мG��<v����=_�y�L�8��E@�6�=(�5���1�Z��<_S8�A��zaݼ��<��<�V5��J�=�,����Ҽ�{�;F?=�)^���<�5b=�t�<��E=�(���<�D��s��<�\=p\�m�����Z=V�8�uo�;
kW=�u�:��<��=��<ߟ�;����l4<����i��<O#�����Tn��g =�j�*���,vG=*B⼌=���~��/��!��;Le:=b6�<m1�<d+!<�h:=	z���p=e�<�-�:p	ָ$�L���b<��E��<��;=�R=E�ۻg�1��u�<��<[�B��<�O�<�;=�ki=�������؏��4���<\ͪ<�&�Bq���<�r�2�h=����;Ƴ�똽���=^��:z�3=v�ɼ�r�;R��<8Iֻ0�A�	��<-����������=YӾ:�җ;�M=�,-��Jؼ@�< ~��C�=n�v�(<�<�e���仜+Q<$�Լ�d=z�4<dE$��.=t�F=��1;�k_ =&H=����8�Q���a7�����<hY�<��	��=�>=,�;���x=���~���+<�.<:u���<YN0=��<�>(�QP���<y�$�=�xR� �=��o��a�x�;_b(=V4;=/K]<w�<�Z�02�<��ἇ/E����;#���oλ-87��t�	H=��j=�Y�<�<���;��5=��7=�Ag:GǏ<��<�Z=]�=�c;O�:��wi����:fO_���=�O=�.��K�<��=+Jʼ����=�Y<=�)=�}]��ㆻ�W��<S=��=�_��O�һ�3%= ּM����l�������<�~�q)=o�<1���rk�P�7��[�<��Q�a;׼�)��hՎ�(�;mT"�Ȳ�=e-=,&�<��a��U ���l�\qܼ��%��qr=)1�	0=��ɻ�(��Qi�g�μ.�5=n0]=U��☄�0Շ=�2P�fp	<I��OS��ť;VN��5�Gkf=�p=]�U=�
;�Aw=��/�o��<�2��F�켉56�lV�Dʝ�қJ�V��<O�<I��:Q� =K�ֻ7�C������o�ѽ�<^$��bR=��/�v�=�N=�4U=��G�Xk�<�J%��1+���<G�=����ӵ=[��<�#���<��<m!= A>=`
!=4�Q�nJ�;L�8<�x �K��<��j�@\�<�}ټl&ͼ���<Q�F��`%=��A0L�8@��N��fH����M=���<S�~={�n=�w<�Q���1��7�;�g=놽"���۠�5N��NN�M�;��ͼn�a=�ل;�ˊ�$1��bh���<~?�<���/���C=�4?���m<`�F<�=e���t=u�J=��nU<����;z�;=!�k�
��9�M=����"W���Q=�	<'�<i�?<��<jHM=��J<ء��(=��h�����̟��==L�R=|�;x��,�*���"�5z&��yB=��{=���<�����0��1����=��<��<qm��\n���E=e�O=sJ�5���+;���<�v���~�k�<�i%=
vº��=t����[L<^�8=�]��=Z��<�Y<�و=3�x=��S�w� !=Q���=z��<j�c����;5�d;J\=�w<��W=,�G�kh�<L=�3��=�d<��*�!��<	5�<%j<��5=����;�>���N;���;�*==��<o�J��¤�s.S��bݻS�]<bH;�5缷��;� C<��L��m=����D=A]�<9�~���=R�L<G㦼;�	���E��<l 7;�����=�s=��82=�����<�H�<6�E=��V���������4�:�)dܼD&+=�Dt�f
���K�Î=��'=�>=�B���<ff�:̇#=��h<yY�ig<�:�����׼��T=�=���+��<�ɻy+=^;��߰�+�[���6�G���-���L��ӼĦ5=�QJ;X_P=3�<>D����2�<�{�	�]=aS�Py=�d⼟�x=yMƺ��8�R}�P�2=6��(UJ�Ϟ�<��8�������w����<J�=g6=�e
��9=��ڹ嗀<��[��g����=!W\=J(�<��]�F�J=n�K�^Zh���O���B=X85�bm��U:�}�����	=^G�<�A=@�v�8vo�ID�<5j=�%������t����Ǔ9=�F��t�>�{�<_�=�5d<�7)<t'I=^N=yy7=׬_=�kv=3�ݼ	X�<I~���Q=���<RЁ<�+�VX�<�:�<�`<�]=v��<1Mx�i\Z����<��1���<��<�M��Y?=��)=Z��;���n�L��EI=t����<�1�d�@��P�=�{�Y�Ļ��;��-��=�{���1l=�!=��u�;'�se'=��[=��'<��9���ȼ�z�<��q< ��<-d�<v�&���6�	�O�k	=Q�<>rr�9�=Y��<��!=�o���R��
&=�G�<J�=*=���=YM=fqܼ%�P���\��1G���-=�����	��(=��<�O�<�	=��=���i� ;^����<e0���x;<e�$=��)=fU=(qw�/�%<3��<{=���;�a=f��<�^�;21;=0o1=�V#=�]&�d�Ӽ1oE=R��J�D�M=&�Y�IC?���<��=x�r=����,j�/W�#R�P;�#K����<���BO=�}(���e����<���<�p��-P�qŊ<G{_��r�K={�<M�A=�=41�%��<;�ɼ�2;��<�m6Ǽ������]��]=�� <s˧;U�+�C+0�<�G<��<�㸼Gm�<L�G�4@�#[���=&�;Y��<�b�=S�=��I��g���8<�/M:*h��H�6�������L=1L=>=�?��6�;c�f�~wY=���<�N9�fJ=�	�d<)T�O�<���<�uX=\�+=��$=�ﻤ��<���~P��h�t<G/�=Jޓ�5�<]�;=��j���;r�'��ZM;Yj�<K�V<�=�F8=��=A*�<
<�;���򺓡�<�]=ab!��-<�w<��x=�+ּ�;�<��;=��:hz<��=�Ӡ;/j�<8[=y�><rI=��Fͳ;��t�,�4��~t<&���:�9�,2� "%�S�8=���wK�<<��Z��ip��<+�=�ś<��<ҶF�dt���-=��E=I^�������=��2;[{�؅�|Y���C�<�ϙ<�?<r��<�k���x�*�U�I�%�JFϼe%=��:��2R��m�I�<=�|��RqGV=�(�c2��o����<�H����X<k�g<�e�5>�w`�#��=�A��E���X=D���B�����<�$�;�,<�=]CҼ�Q�<�6��ڼ�?���,=\|=�2!�>Z[=�b�8
�S*$=+���z=��=�:t=#�+<*$='�=Ɛ7��1��D6�L�S��5�=q/���6��]h<���<=��<ԁ���v���K<b+Y��r�<\d0=�R[=�d�<5 M���=�M�	����P<�B��C���=��;��+������=ԪE=��=A|��9�{=*�M=.��<^�=y	B�6��U����p��
�#��:%-�I���1=�@�<��N���9����b=���=�����F<�iI=H4�J��&��:�N=ދ��s��.�D<����u�9��<�#��=6Q=_�&=k����P�<���$)i�� +;L%�lH=�<]�-���ټ= �<62��� �K����/���n�:�)={�<��;ܵ��\=J&�;�<L�=q�;������=��;0�?=~w'�iwN�]GE=�坼�5(=
&< n
�����1��<����l9�\5#=!�D�6��d=�*�{�u�v�6;��'=��B;�
a<	AH�xh=�R=��=�ZB=�����:̐�����]�-=X
Q=�s��Y�m<0�=+��:�<M@�;�ż����Ǿ�6tB<��<BǼk�<� �>�<CW��@R�D$)=Ñ1������28��R=�]T�<���<j�=��)=�˼S`���NB��xJ=;,�?���;�%����{\%=g�K��9���J��r6;ù9=����PG�"���z��<鳥<�����Ǽt��ID�:�o�R==|���3=w>�<��d���5��*g=�&����n�YY�;��*����e݋��E<8@쾼��7����:]�$=�E;�<E̼��#=`��S��M�<g.E�9rT<F�<���<������<P����Gw��\B�d�$��ُ<�vJ���<���$w���L�J�T<���<j�4�Ҥ�<�4���?=v{(=W踪�����9<oka��Vl�|El��g�9%{�=?�E�;�8���h=w2��6�;�?�<:j=�zX��ԻRv���1=FAJ=l \�WY=�ռ�^�<_�;F���������t;��Qns���<��V=C-�:�=���=�c���d=�lR=�z=�V̻�I;H��<��:��q=r)L="H8�&�� �O�"@����<��b=-{:���=S��]I�ӯb<���{2O=�o=��j�Jwh=��9��&=�v����<� �<V˼�0Ӽ&��;4}���>=��5���9��=<o6�9^H�|s��=$}=(�0=�z�<w����{7�ւ�<d<�<�7���=�hw=	>�;��^=��C��}U�ݻּ4a���7=�1$��M�=�'��]=י���L=@�Y�ҴQ���o�ط<kf�<Y z�p�.��4�<^
"�W���}�����y[�m�<Q��Ƽ���"+=#]>��������]μ*z�<T���"��Ƽȁ*�5��\=�*N=�V:=��=D����<��<�.=����=`�=���x4��?=�aμ�#��a=+w=!$�<f�<M\=�k=�;K<�W=8̘��!����#���<�� =B,X=�<)`0���<��M�.%=��0=�������:jl�b��!�K=���<Kj&��T:��̂�Hj�<�W=>�=XdA=ꅫ��zS���]= �D��\X=��c;
|Y<(���<�B\<A��;�!W=��6=(r����<�Lo����n�p=��<��:���<pҭ�׃�<S]\=q�^=��=���<��u���E=)��<a�G�<�@�<WQ���������+\�<��N=m'���j��`=����zz
:�4-����<�5<�w<u;=V`?=m��<=�=���|!D=!#�7�.=kF�[�T�KT[���=W䠻"��<�a�^�<�=o2¼��%=R|:],";5E�<�<���<��=(=D��|n<./[;�!�=N�d+�=�.g�b=zD+<a�8=�h��b�<��"=�!=��v�YX=���G�=�0=>[�DB�<$ú�oB�<\���4t<>Z<�{�6;3����a��� ��=��y�R���n<_�;HP=�6X=��?=x���,�1��;f�<M6�<q�<�)&=#���YE=�=:��<��[�Z���R<�>�<�����&�m<?�<O�@=������<��V�
+^=`�M<ep=WF\=&�t=���F����j<[c"�p=���v�+���Ü<hS��t$=���<v=4����R<�q�`__�ڻ����*���-�V�C�Q:�W*�<��B��X�E��o48��d�:E��<N�*)P=fYܼ�N��Ǩ=�L=jAE=�ž�:��H��	�i<`��:􄯼<}<33<�$B�G#'��8W���Z��Q/=
��1�{����<oT��5� m��vS=���v�%�����A��%�<Y=�ꃼ5/�<�k�=�3z=��<N�W���<şG�rڈ�j��9�7=��Z=goϼ]f�;mG�;�!�<��D=�;<
��Ք ����3��O�(=eX�;D?ż�����=�<��?==���︼U�<PA�q�~=}����V�S=�'H=P�i<K�I=�|��k�=Y�Ǽ(5&=��l��6$�#�;��U�<r����;<	�V=�%V=F�<�����<��:=Kz��<�kz=�튻��ʼ}�<�.=�<ּq�`��=�C�<Մ]�\���;��=���<�*8=1rƼ(����^=��<杬<��<��ۼ �X<���<����;4C��=��j�,&�;��:�m�R=ɼ�O�J� �������=l��<��7���;<ͳ<�:���;�un<�;0�8jQ���<=���_�N��o8��=��f:�=|�0<'ڿ����<]r���<��(=�I[��_s��yy�Å���\��Mof���?�O���N�9?�<o�|=J<=�9��N=���<or=R���)<y;=��=H�=��_���6�R�o<�U�����v<Ӓ�<�ϑ:���;ҲR<L����9O=��P�̼�<�i���<g�;T�ȼ��]<���<V=w��<D�%��_�� =�[8�\.<'�?�յ>�Oe=�D�<��<�n<&����ۻ_I���z��S3��g��n��:U�6=#kK=.ؽ�'�'=C�^���@��p�T�7=�a<m�7=(e��tl=������/��G��&�K�c<g�3=��:�*;�%=��+�O���=h2;���˼`��<���<��=� k��%����r=S���I�4��<�> �����'ϼ�
+=q�F=����)=�Τ<y�m=��[��Y�z����K=�=Bk+=};�pM�3֜=A��<b���������:��Z��N=x�V�� =\�A=�|<-��<ob��d>8=;�*;��=yF�;�G=����C=�3=��<b�<�=���}�=��.=hC=���9�����ᗮ��;���[��]�<x@k�I>��ʖ�<t =��"=�bq����<'ي=w�=cx(=�͑�M(1�3�<)�_�Ԧb=t+$=A�:�B��j:=9�E����<�����A�L�v��զ��_�J3;�<�<�p=|6�r�<R��&�b<
L=BZ���)��Mv=y�X<�c���'���ջ�B�����NͼD<S�0��<\}<,�6=>��6oJ,�۰{<N�=c���F=�U��vm׼u�;��v7O=2�7=ّu�(�=��==��=d���<�	�[�"=��=�b=�%���b����Ҽؔ�;dX������4�"��
]�������;gn�n��<K��"�����<_�"G�;HP�~v1�_�=s��;hy�<���@h)=I<�<�1i=��U<���<'l=rHż��1��(:����x�^���ͼf?<��<��Y��T�{��<��<��=e#<3�j=Q�޼Ӑ��]?<�o;�?&=�;o=�e���dȼi.p=�v���i-:u���0y�z����=��=�aB=�=���<�x��m:E��?<����<+�z<e��=Dlr�u� =���;��$=�]=���<)\�L���YF�Btf=�E=�!�<�钼�PƼ�!�}y�W�</�H�<
\��L�=��<�z���6<m�<?�&� � =�i3=�� �,�<Lt-�3�[��z<�+=LļCF�W?(=@{���J=�=�fH;��ϼ�n��!���q���&��i��{<<� b��ꔻ��-�#���_��4��2��*��R��<���:�����`:��N=�o(=>!2=5d"�j�:	�(�2��ƨP�~�=��L�O}üI�$�%�-=�K��U�9u$8=�P�~0=���<g�Ѽ������r=� ���=\JD���I����<��F=с�<P��q>�Q��<3o��b�b���9�d����<)���z�t��+=��=�8�<`0<=:Z�<z̷<���=D�C�:U�<T<�:J��d�:��$�:�/�-7ܼ���<#��;ǻ�@���=i'��l����]=��.�B�yxҼ����@�{]N���J=j�պ0�,�R&�<$�=v^��_��;k�
<�t�<�����=79<=c���B�P=�1�<hi =86���0�N��<�$6�3�<1IC<Fd<=����Ǚ����P|�;m�= <�<q����B���2�;���^J�ze*=�@"=��<~��Ѐ�/@��H|<�g�;���$>��O_��ZP�ʥ	<Xdv�r��<�ē��d=�i��=<-�<��=��5=���<��>�eGL=���<�y*�P��; ���p�<1Q=tlg�K���O��|�;h�.���s=ɘ<��R���(<�X6��.��\�B_=�<=�]L����ڍ<����2m�<9>v�lEV��K%�[�<��A=���<�4=�&e=*�&��\�=ͦ�<��,< `K;_�����=rA9<��92؟<�3;J���|���C��o��<S+�(3�<�;=�!r<����=�;��O=4�O=ߨ�]n˺��=��� �<{�1ռ�Xc=k@�<f���L� =������<7����2�.��<s$g�1pU��h����O��h�=�&9=!�<~�6��D=�Z=o[%=Iw�<nb=p@q=�)�e+b='q���,d�]��<h<�&c#=\�a����<�n����ᄼ����2�;��<��<>Y=�o<�V��)�;��
����<��1=�V޼�I�1]���˼�z}�&w7=l���Y<2�ӻ���� !�ߩ�;�H���@*=m�i=X�j=ھ�|��<��<ϼ�<n�<z����=Kݕ�����w1�;���<�����<�b�<zn �����7]=�	5=�SD<V9��t=iRs�tDm=]&���u-��]��Ί\=p7�<��=�<�7,� ���&=<�|=�<�<�cF�R����L<d�v�>7]=mAO=$������`�0<��=�%�K����鼨���R�<��-=�Z�F����j�<.�5��Z7=��s�5�Qd'=�3W�P�����)�E=�F�X2�iT�9	���NA=���A�M�����8(����<;�<�A�c�E���V=1�X<h!�<��@<m�a<_ =)R��P�<B�l�q*4=] P<:i�df�4<��+��]���-���)=�4=�]&��s7��>�<�%O�uc��&w�VlY=$蚼s�z=�
�BFt�.�<�;�`@�BGD�����#��<�n�<j�G=�Y�<��׼V���^�n�;=�6>=��9tS�<��n=#=��C<H��;��,�6#:=DH[�Q�<��e=YHW=���;�@=�?�ϵ<�y <7�<:�5</�骙�j�m�s�b`9�E'V��n"�Ɉ����3=�d��l�;#ー/�V=�+<��5=9�<�LA=�\�m�<)�f��E���Ƽ&����� =m�ͻ�#�<�|��0<�3=xxb:�0�<��<O>�7=���<�=A�:�<ܼ9�=ou=�H�<���;���!����&�;�o����<lǀ�O�;p�U�o�W��Ӗ<P��<��(�<N���A=�0=�GI=�Y=gG>�o�ܼ~�)=>�$=i��<�t^��*�<�B<TY�����;m��;�sp�;Fּ�^!���J��=RM�<],=��'����<��P=g��������~4�&��<q��<G����R=>O*=}n[���s�Ǖ�;��b=*@�_&=��<��x���0��~<�07:��<�4ü��\���@�@BD=�(�<�Z���ļ��=���T�<x3��n��C<�̢�nn�<�/�<w�<'8+=[��<���<�<�E�<��2�"4�=�N;H�#���
���]=���<N<��D�� ��z�)�������{IA���g�G�e
;��E=^<=�MN<���<�Q�:Y����S�z$�<�J=G)x<��=��<��=Y��<!4r��zL=F�<���"�<�1�P;�M�=��B���=����(|;̄�<�*���=��*=��U=�4�d�e�������+=Qp=�_Ļ�<�;�H��＇�ļƉ!�
S�<0t#=*_C�,=�}�\j����<*��<6�A=�4�;��;6A�`�4��iS�x�=��e����<׻P="��!��;+���}��9��^���E�<Q	f������j
=�.4<G�?A1=���<r�X(<s�<��=R�ʼy`K=L?;I������;���Pl=,�<h,=�Y�q���y<��<KqS=}j?=u�|=�缼1�<�F��@�-��O�<&�F�3�<`q5=�=Op�GG!�f��:�b<�"�<��<��=�u$=�_��i=H8)<X<A�����&���<���F�G��A����;Rh�8��E&N��;\�6�R_T:�KA<�ew<���H=��<L^�<�J;���;r��<� �=�@���!;{eY;��=1z�=F�<IdY��xK<L�<���<Ǭ�3��<�����<6�ټp��<J��<�=�����J������3���<1n=.�$�<�m	=�J�<4���O�T=ڹ�;��!��=P��aT��O����=��=���4��Yy�;1�y<�\G��>>�Ӿ�:��ʼ_P�<��=!��<��'���P=C4�<�w3<����?=I���i=�}{�fl�Ok
���*�V|<AQ-�������`ؼ%��<9��<Ӯ�<��g=m26<*F6���.=򶔼��R<L��Y�t���^<�G�<3��;���<� _=ݏO�`{�<ÕP=��u�f���ʅ<�D��+N\;�EN����<¡m���|=�Zw<��2=	�=���<�鼤n����=Q<��V=w?;���ֻ�AY�,�5���6=�<�j�<KżJ�ż3	��<?�����}Y���1�;�-=j�)��,��64b��:�:s%�,�e=e��;K߼�̼�
+�*�k� M5�li���2=֗���V��A�J�<���<�Pj=�@���B=�G��GN=��P<�e��ģȻ_��<2(ؼT�7�n�`����<su-���������F����{��<��"���̻%���#�=�(/�|bR�+��C�<�<��%��i*�<g<={�<�I=�ˊ����PP:�~����#:x3=���Q=�H�<�����<�j{�k{P==����,=1y�<"=�t<�K�<7΍<��Y��ΐ<q U��/ܼ"��<�l�=�[*��嫼�U=>��<̘�<��
�l��9=0���<��P<�q4�t3=F�=���<~ӼxQo<4����<~w����>��p�v><��b��E����<K.����1<}��; �o=݂��C�e��(	�y�3��/M<����0G=�b6=���;[��<�0l����p����< �*�BT��!2��
�<�T����<Wu�<�֢��H���-�;�<�
���G�0\a=ʳ<c�e��X�=k=�ؼ��i<��$=����9�<�)��S�u�$-=��1��� =�)޼��X<q�g�㺅=�8�κ;߼V�B=MU
=P��<=S���d���<=H
p=������-���b�=�/=�:ռT+<�!u�ar�ٌ=�M�i�=S�=��	=�[=`ț<��i�OB=H�v=(b=�,=�wN=�u�<"�:=rh�<��^=H=}=耄<�=�<�_�#���+7=�U��@/=�Wȼ�p�o?�O#�+�8���u��#�H߈�jGȼ�w�<�b���s=N�<� ���Ȧ;�s�;�0=GJ�l�I��W(=��G=�(X=�ӕ����83���<��<�|/��(�o�}��p=9J=V�1:���<���<ᜳ���d�bzX���D=��5�N7r=��e<�k<]$=���<4=�.ļ'y�!�-=��s�C!]�7_�uռ��<�R���F=]0�<Gu\�TD���E�t=��b����g=Ő4=n�\���1�W5S<��#<���(4�<-�1=
Ʒ��؇8f=���<�8���E�_fq���`�w��l	�2==���js�X"�<�_E=Ye8�y�<��ƼA5\���1='Dv�{6���=��=��Q<��S����:X�;��w<��o=,���?=y$c�g<@��D=��"�������9�3�8�PR3��D=�F����N=u}=�r=hLV<�4=J6$=��e�:=���<�"�e)���%N=�tX�T�2<�w2��b<n��<?$F���O����<:�-�2�"���j<��8=;޷<�6��=�b�8�����-�6�.�c�M<5=LF	=��$����<��;�}B=�t��e�¼��Y=���H��!�Ӽp�#�-��}�n=�$=�꼞sU=�/<��<��j=�A=<I,���d=��[�o�"=a� =������;Q	��p=H�<��<�8=P(,=�;+�"�<Ϥ���1�O�M=Ewg=�\=+N�;λ&��M;�겼�ډ�иN��/��^Y� ů<�6=W�S��#���F=�e+���s;`Y�Jp"��X�<�E;C��aN,�E�$���<���<��E=�?�����;e�<��;Z�T=�ȼB�?=|���s�P<�
=ӧ=Ҳ�<��"={v��M�tE�����:���<==�O<��J-��9K���=�K	M�pq����<$�m=��!��H=]���&N�>���ȥ<��;$����9
;�E�<�><`�<J��<w��<U]2��*8��T�H��<�������<g;��\<h� �Ӑ�[�^=��<��a=]V�=؝/�����ݏ��!=B9<�v弼��Uh=�A�iB�u�;����$m<H���WT�<�8S=��<�R��h=<�O=#A�4��<��X�D�#=�f�<�3�K��=�3t�2=;6�<��˼%�꼣�I��O�=f�
s��{|=*�7��m=y�<�u�<���
Lb<��K=��;g����<d��H�ܻ�R�<��a;�Uj�_��;IE9�����5�����x�<g4<ԗ+=bŘ� $��ѻo<��/�>$=t<�;OE�;�Y��{��<�L�<�8:�Ȕ���<̒=^�<��ϻjpi�z�1�;�T�;� ;C?�< �;o�1�h�=���,��;�U޼�z�76+[�
a��ɉW=��I|0���c����zS��ES��Uӻ��<P.����V=����j�;=�d纁9=Q&=��K��:(�:�<w!_=|?c����;v�8=ɜ7=	����<��<=S�L<I�=��g���ټӊh���:=��H�yJ[=+�ֻ�W=�~�<5E=�*?��4/=gc��<�z1<$vO:����mn��J�<<8=�/~�"��t�J�
ў;�L��f8�B�5=U�ѻ0<]餽M�=��*=6�)�b�	<��1O0<�x[=��J�ڞ�<�9�r�<U`;�J2<8�*�R9m=}Y�����w<2h\��g�<;r�߾<�HC�n�F��(� �B<��q���ָ��|�LW���B�50��F�V�A��/V<f;�'�M=j���
��� [=%����Ҽ��
\����<{V6;�I=�#=�M�`'=���  ��i��'���?��bB�Di�n=�@[=|U=0�p=����(� ���(�xǈ<�t�<�����;���漊�=�;_�
��"":�&=TR=�u;u�=��?�w��<�Ś�D�t=�d���Ky=�P+�*]<Q���ẽ=������A����5�&=+l=Dk,��#˻�Dq=��<��%<)Y��C ��&n=����s���~>'=�}<��=y7r=G=���[=p�ݼ�1=��=7�����=W�=�9��S;UD��������k�s��t~;�`�ڡ����"�'eV�_�V��o�u��;a�B=��S��M��+J�yQ=�K�<�����[=ß:��3g����8,�*�=3z���;��`�J�������{�輫�F={&�<���<��=�� �4�
�2�>2�/P��0=�z`<9�S���}�z
��9O<��s=���<���Rj����)�k�6
Q=�`��0<@i*���<۵μ��<ޏp=> :3�ڼ���<��Y=Vf�<�,ٻ)*=='7m;�Lͼ�*C��Pz<k��;�N=���E<���<1C=B����������NT=d��<��=��)�fe������!OS=��<������;�-�<�z;#=�$-�a��oǼ�-���(<cĦ<�9=���N2�]}|<&�=��
=�x=+p����<Fћ<���U�D��,(=�[��+�<�y= �&=,I8=�u��X��ZKK=�Q?=1V�<o����w��;�u��'��<{?�M�Q��A*=%ٻ�������]��5H=��5��L�<����<��ƅ�xZ�<��_=2
�	J8='c&��l����Mx<P��)��<U��;G�N��K>:�<;�Y
=<5=b�뼗W˺n�޻:�	=P%=bh���=�:*���<ϯ�<�%ͻ����g`J;�"��8=� F=��+���N�>g�<(
�7?��/�<�̪:��=Cd	=�j=D�������K��<�%Y;c6��A�Q��lc�P� ����W�;=��m��Q�p�/�U=ƌ�<"P<���C�2<�C�8��3b����<�+�<�hP=�ӵ<[=+��/_���h��H<s�/=jx��
��������`�7�.cc��_��y�c;�?��z�n�%=d�N=�<sg�=���<���Z�!�1��<��J=0��<�ݥ������}_=k]�w�==C�s=wg���_���:�A<�F>�4�=}W=h�
=��E�N;<+j�i�-<;d��3k���A~�y&W�Mo��D�<�˟9�:8��ʼ{��<t�v�`�U=A(���<a�c<� �<�-=R3�<�.�sm��s�%�A�B�=�&�<Օ�1W	�{W=F�<de��ԏ�<qY���<a= �'=��$���ܼJ=��=�8�"]<���@S�|��<AF1�u�����;_�l<�­;��s�so�"M#��H�
=RRC�}\߼>kj�V��@S�<�M<��P�K�輷7Q=�0Q;��O=��ϼ-�:��3=�n= �N=:ŋ<�
/�c��;y��F��<.�
���-a�<�E;��z<�:���I=8��Y�\=�3�<�_&��O��=�`'=�M-����<hDA������n=�����
�P|�<�=�=�^<��ȼ��<���:A����a`���x<r�L<�G��F�(li�v�����<����<��<�@��wr���ػ�悽�F�8��7�d��ё�;�\/=��N����<����븏<]l��߁Z���(<�g�ט���i��H�%�Ϯ�P=�ּF{;��;��</��;�<�Q�:P�.�ζ;�����@=4ؘ<D�t=�G��dʹ<څȼ�Ƽ�*�<��D�-Pk:T��<3��;�H˼4,��N����[=2%�<�[=+G&=�i=M`<cÈ�(6�<#6��|HK;��R<��<�4 ��HH��|F=��;B:�=��<��o=�1�).=�,j="��<�K�VB���)=~�e���¼�7�Q�u=�s<�Y�ϊ�=Y=V=,=@���=Xml<�;T�,=aG=��3��>�C����]=��`9��Q=�}�i_7=l<��0��o[���+=�m���X�|�Q=A��US^����<>��<��<�=�?�i�����9��2��o J<%;�4h=%�_=�T=*O�=O���ֻJV;;��=pX=$.<`9<9�ܼ!eF�S���&�!=�_)=?^��N@��>;Q�N�O�|�F�>��;���;������;ܿg��;ۼ�(鼀�{����<����7�<�eH<{���+"=�5�S#�h?(=f��<D)1=�������i�B��� �/<:<��� ���?3=��<|�p=�a�'6���n>�	����M����<1[H=�䅽�$<��<;E��C
3�x����%����3��d=�==�Ϗ=R8��d=���;q��:�)-��-ۻ��=fv�=�x�=$����{k�G;�<�Hͼ�\��#�<���z��K� ����<D[�����S�<u=���<��N=G�b<�<�E=�=�z�� =+�=<Y�;�<�6<�=8ټ٩����Ӽbo��+N`��W�<݈`��׼���J5���.��,F��^
=�z�<�4�<Q�@=W#�+��y�<� �=�	����*j �'q`=.;E�ͼR�ٻ%]<��7��(�<�g=�s�~c�3��<�(:<���!��s���=�A�<�+D��-o<1=s�<��=#Z�/a<F��;��:K�$��|5���.�iy}:�5r<���;ʂW=��)�.*=�=�2�#`=o3�=P�5=ܸ�=+���
g�Мϼ�l<_��< �<�G#=�>�.<���@�6iZ=��<�	0��!޻\(/��"w�f�:`C�;�#`=�� =�����0�<pY��}�A����<� <� =���N��Ҽx=�E=`�J;Tu�R������:e�=H=��ͼX�:�*=|��<:���8�{��<�
�<XD=_�+��==H(z�H��:�?5;�e=���kζ�f�L�(�	��<�fʼ�Ii<5���<g6�=պ9=MWv��<Wp�<�fw�R�=K§�F��%	<�xU����K<�t-=h��=��;"����]�u��<��;��!=^E��w�<u��<�<d�����I��R;�#��ʫ<���L<SJ:��!=H���]��#R���a��t<dRE�b=ڠ�<���Di@=�ƺb�ڼ��=�/�3�<�z<���<oE��n��;JQ;A~=��C����<��K=숽h&,=�旻!��=�<���<�)���<�-.��u�м���� _=m�m�v9�֊L;�3?=�'�"���s��h�E��<m	< T����#Tj<��q��<#a����:JE�	Dl;�@7�h2 �˝<��g���_<tp�<j�I�[i=;�t=�h�������Y�=-�<�g<�d?<4S'���&�Z��� {��U�<��=�g;^��;Fh�;cMr��Ħ���/��O'=�C���
f���=F��^�;o�F=��s=�C<([�<^���<-=Ȕ�<�+<|��;j@2�T�?<�_���rN�
 ��[��>��;a�4=�>=/�N=��Ժ%Lt�S��<�B��NL������E<���g��]%������|=Dū<���:�_=�8<��P�F@�#��s����<	W�гN<��o=��.=o�$<����W93�9֌���;j�x=���8��<i%�<7��<Vt.;�<��V� \�����Ƽ.d=T��˶;�a5�h)=2�H=�;<�鼾$=��׼f1O���J�6��恽fA�<]wȻg|�<�쵼z�<���#r=$�e��A3=��J���F<�5�<bw߼�'7=[���W=1�.�_��4�f���]C�<��`=o+��P=�WV=/�< �<� 8=1`P=��<$M=���I�&=��=F;t�^� x��R�����;$�.��Jc<R�`��-�<I�B���s�=�"K����-�=�
��k,=��=/��<I^A=�
8=޼E<ޗ(<��<2ǻ�%=jDd<M��<Ti^�1��<R�м9Z0�}�;�t@=���;,��. =v,;0I?=�F;G=�\�<�AO=���+uR�|2���<L*/=��=I�e���=d�<ξ����S�K<�����5��������;]�ʼoF=^)A=J����4=P'm��NO�+��;�t�;�=�:�U=�D�=sTR�m9��sQ=<8<v���Ug��*]�
���d���Y�<� [�4j.=��u=��MR=�X�<�"4=�󄼋E�oS��e���� ��B떼9Rn�j�s=�$�I{�<�{t<ؠ9�y�=T�C���U;4��<-h����=@:���~ļ�
��H��ܮ<���;�g@��c0�4��ے��ca;.=��_<!k=����:.���"0�=3=՜��=�
������<��G�b���=�t�3���)��f$9��sr=/��34�A��<�)*=*��~6V����;0'8��̻q�I�����м���<��Լ���t�켇�N�h=#�=�kۼeu�;�?l�y�b��v�;G�=��=h�j=yY=��<~=|F��z��r��;]y=|"/���<�	��E"H�8�"�R^�;�Q�;��2��=�E��)A���M;D�;Tj=`�h�DS-�\��<r�P����j�0=�����"�M%=L���6<<[m�I(��,�_=
�m=#�ݼ�?μ@����<D�=�)̻Ǫ��|=�V�ܢp=T<==f�R��H��gl�r�.�-I��<��e=��?=j~̼8�6�v����^��E���DG�ޛJ=�~߻6�E<OEI=0;=�x�����Z��<�%��Mi�r���ٻr�����<]"���������G�=o =Ⱦ�-��<s"�"3T�ӓ=-w=���=��˼K�o94��F���ԻTku�@��<kr��.��O��L=�7=�7o=��;<*h8<fDK=|bC�r�ѼԊ
�V
�<B^=�)=�r$���U=!�(=C�;��=�mk�2�=Y�ټ�[=��R��z�<���<�s�<L�x<�gȻu�3���V<5f,��7�B�˼rT��h�����"��,=�O�@�(�7mB�5�O�:�7=!��W&�<�-��P�;��=�v
�o;	=x[5��c=&,�<��=K�<�a�<l�%=i�ͻ���o��n�;�=$T��3�@=�E� M��_&=�
s�L�;M'�k{�<Vƻ<��?���s=��s����b��,�<c!�<���=�E��=��;Ժ&=Ս�J�q�/h(�W�5={M����=��⼗g=D�==�8
=S�J#��ύ(�%9��F���Q�T=� =�;O=V���=�=�H=���;l�;⻯���=ae�iDh��j,=lH <cN<W�'=,R=$���=8p#=*�#=�H
�g�8�x���Z=���6=[Dz<]1������3��e��=���3|��M8�0"=�n �:A��<��:������w=���<싸;�+����asq=p��X`a�{��۞�<���<L�'���C=��d=�Et=z�k=�a���M<B07=ɿo��L�<G��y���<�>%�G��w�V��!� /�<�uH=�촼G�~���<��x��2;뽯<�K<��G<`Bڻ�wF�dn���[=�+�;} ��L���(p<���)|m=��!<�0&=N*�M���ޚ�� ��<<�F=�<����{޼�E�=bI�$�\=6�G=Bf<�ŘF�p�U�z>F=`�<6J6<���s��<e�i��=v�T<H��̙_<�,=�J]��h��`��� ��}�;P��1��n�h=S�t=C>�{�Ҽi>�=�����=�<�G:�E=�+==Z�=���<<�c�/B=>���46	�]�I=?�=�'S=�g��[3��2K=ً+��w1���;��f=�!=�kh=D�<e��<��
=.W+=3q�<��A��_=?T�;P��<��=�E=@�;���Z�`=,��;IG�3�<8Yu��|u���	;�1�<�+�0j�9��A=�\Ҽ,jJ= 3<��	��K��[]=��<"ؕ���=ۃ��:�	=�
(=�i�U�����<�J�4��;Q��<J�[=H!�;~��;�A<��]<��+C~�Ip`�Դ)��s�<P��<�m�<U�|�<���;yw=�
=(*=��F��a=O�5<�A���=�=��Q=}0�<L�=����P��<����M�1=����(O(=[�=�h��#<7>�<
�n�(����d=�;Lʼ�U��{\=��%�.�ϼ
�+=m�4=�M<~r~�y[q���?�KmL��H�ץ��i���=Α�:��n�6� =���<��o��q�<��6;)I<��=��i=0�[�q[�<d�#��~�<{)���P=�Wc<�Hl:�TJ=�@:=Z9=�\��.�=4]S�BX�;&���N�<>�<V��Zԙ<H�^<_(���I={�ʼ١,=��<���}��(=��O=>�<��:�;!�<<5;�R\���;7E=O�<�벼e,�<�{���"$���=����
 =�3/�x�h=|�ͼF�==p=�������%�<�PA=��6���h;GE'=�������<��<0�69�[���R<�;�<���9��їz��l4�����r�=È�<r���ɂ��T�:`=�-=��A��<������<O�=���:��>&�e�����=�X�;W3=��<��@#=M+=D��;��<0Ж<<ˮ�
�8<F�`�a+H=[X=�qg��*��JO <�^�;ӧ��d<�,�<� |=��E=�7;�w��<���z,��
�����+/< �I��{O���]��K;��<��z=���<kc�<��;�u%=�=zo���*�WB�<��L=ك=��H���<t�,=HF_��˼�jc�.K=]�=4�/���y<J�%�sFX�
1�@�=j鈻�L;=��=,�=)�����	H?��=�AF<+0=v�`��z.�ˀ=��=�%�<��#(��d���F��\�;��G<yI���43=���<潢;�#�x�m��q=�{�^�K=92n���[���;�HQ=7��<��B<W·��M������f*=
��r��[-�;P�<�ml�ʂ ������ˣ�\pt=Wq=�L�k�<X��q&=,<��t�� ���<�!�#�MG=k��<�߼��-=ܣ��һ����;вB�Iq3�!��<��ߐ=��N��üۛ�;�X�<�ho=ܰK�0�<8]f=�xo<H�=b��b�4������_~��twS�|6��X��<z=��Z=�!�:~u�<���<��i�Zj'���;���~Em=}�p=�Du�<ʼ��<|ܻ�#<�`c�����r_��;������%�<�fW=.�j��μ'�3�N}<��<����.H����<�tF�Z(��,��1�	��B=[Zx�
苻ƿ�<�,�<�M=�kY�� T=�Ì�ԻV��7���%=�Z;<���<�/<��M�?�C=0�ռ�IX�8%=oɼ�a>=�b$={� �)y!=�}����2�Yy��IB�_��<D9�<!<*=2$��<a=�Ze��z�<	�r��e�<��b�e��m�Z=萇;�Y<?N0=��:	�B==��t-���{<J/�=L�Y��J�3PT=�8<ǅ鼈V<g�<3|�<D�<Tt�<�̦����=~ꄼ��+����
�N��إ<�b�:�ol�l���=Cl<�eg=!�f�z	�:�r=�[��|<�8��E����;sJ���.��Sܻ�%=�=��k=��~<+L�9<S��w��歼��=ؔ�����=�3�O ��2=�5i�J*f=^�=�������vУ�)���@=#g�E��;(���{h�pY�<X�^�u9<'��<�4�;��c�;C�9=��y�%Q�<}���B݁��a�C�;)1�]+=�p=�4��E*=�w�dA���YL� Ao<'�I<ԦA����O,��ٵ�$�<rE��A��j��<�F=r�f<X�=,�μ9�f���
=e�����<:(�= �;��0�7Q@=U��<'`=�;1=A��=�L=��	�o��<0������^��Ay<�i���=��Kr=P�c��g��䡘�y\�<���9$�-�q�Z<��=�踼SS�O-�:oJԻk��&�:=���<(�<�*�<���<�L���j)=:s�<Z#�<C��<�E=�������<��)�q�+=G�>=�?���Y=��G�,)2�2�b=�A=Ӵ�=�
�K�=�^�<h14�ǿ����;��D=�1=��\�yYx�R|�<Yyj��<=��<�N��Tn2<@$=��)=��<�zC=}3�25��H8
=W���>��/=���<�c	�6��<5���%�=�P�<E�=u�'�*������kx��
���O+�g=��=6���V��mƻ��=qR=�>��ݱ<e�7=�ۼ�j!=�R�;T�ûV��<�Ɨ;�(>��k�<"pL<���<;�<��̼�	��_tü��:=��=;�<����dY<a>O;���<5�A�4��;� F=_8����$�Yb;<Xh(=�0��鼫�Ƽp}J=�d�<�m�|ᔼ-�~=W���\	�	İ���b�,�<��c��[U<�@g;Q;��ʻ�`�<E�滗�<0�N�Ņ�� S#=���$�<�XN�%�L=ĐC����k�;7TY=�=<,�¼:�L�t�'�G^�t��<���&�R��S���&<�1]��x�;��<�،=�6�^,�<V�L�;�߼�2Ҽ�%�;M)������$=���<��2�I(�0`Ӽi��0s�<��!=��<N��=��(��%q<��^=���<��I=�_v��@i����&�.�9�C��8�[*�<_�H�Js=r6<�*�<���<̼w=�H=���;VF�:Y;��*���<��C<�������M=<�>������B3�աu��:黣�N=4�=K��K�;e�=�_Q<�Y��Nu�/���c��<E34=`5�jGJ=�<����:C3���R�<�fۼ&~9='m=�z�Åv;,K;;��R=��:��q����OP�=��4���<�W_:h�p=p��6�aY@�����]��<K7��Nq�gp<��T=Ǜu=��J<��:T5��0��&yC=C����d;��o�2)�<h��<�u���yq�;PK���"��1�;#R=�I~<k&+���<�J=���9�d<>�i�,�I=��;$�p;�9�l�l=B9H=���F=N<�'=�G���r-�ӫ7�2�߼x^^<�=�O�ol���J�ɣd=h8=;L����;:_<�
ƺ=M�������&��<~��"�Z<��:�|�����;�����r��$\'=�z�<�Ǔ��>=y�<�N�<��
=g������U�:����}���;=S:�<�H5�M�Q�K�����Ի��=��<v*E����<��;Iؼ9 ��b=l��!!<��\<�����ܽ��nI���4=<�H���5�$�<S�,��3 � �u=�
�;S5ȼ�߼��)2�*�p��ݾ;b��;ri�<�����E�<.y;m�<F'�<PR<K�=��O��^�\=��=&P#=����A���R�j<�r���s���V���%=~<<�'=��+�o/�;i>��F�:A=2NF=��&=����<��=��)=��<�u	=L�S=urH=��|�C=��ݼxC�9�D�;�6<���Th��؃��j�I�<b��<.�; �=]Β:)�O=��Ӽ�i�r���n�����ú�3=ٹQ<f۳<��=/�����2��;!��\�;���r�*=}(�`�!=�\=B�<�_	�^�ּ�z=�y�<ף�<�XK=F�5=��9�X�f��rf=����
䆻��I=|�=a�G=-��<E�H���c=���=��<��*�p��e,����=4e�<Ӭ�<Z�����n��[=Θ�<C�@�7�R=̈ =����v �<-vg;�c��z�:��*0�+�����<�^=�� �D�ؼD�˼�3׼n'=@��;�㜺t=^6=_Jm�e�<�Y='�6=QP��� (�?��YfX�[ m<�;R����;�ߖ<��-=��<
W�yh��q��F(���@������u��'�� N���<a�;bG�t�x�1u=2�M=�=8�T=;�v�����<qmռBf@:ma�P��� =/ =J8�<Q�=+R�jk��|=���%����=��L;��,����λ$�L=r�:�@�g0)����;�/<
��<���:"�`���3�-��$<<Z� ��Ll��~=��<x%��=�<���<�;��>=ڇ��q]��
Z9=ڡ��xi��<K�$=&�6��H�㞎��� ��!�<-�׼�4�<��V=2=�]\=KL=�F��4���o�,;�-�nI&�{�<<6z��	?��^a<�掽�\@��pb<~_=�N}��QL<ٲ��ܠ�=z��<�N =z�s<��<WJ�*�<��=[R�<�u��6����CS=t��<�SU=��d"=o5*=,��U�:p�;!w�:(�b=E�;CD=
Ǡ<T�gH(�0�9=V�X�uoT���!�L�\��<{|\:S2�<Uļ*�g�:ɼ�@���,:��g��޼'���ѻ^�*�tOӼ�=�g��,Z<��!��{Y==��=��:��<��E=]�]=������1;.=�w=4rP=�)��p�2m=���O�<InV�_q<=�T�*f"�<g���+��T��ӗ���ɼ1�B�����:&��!X=��q�G��Dwq���8<	5_=\�����å<��&=�g�<�r<�e=l�=�剼�:t����������;�ۼ��=p0�<�m�O���<A=C*�;2��<��==X�=ԩ���<�t<R�:0�B:��A=j�<������Q�E�;=�0j��Ba=�ļ�4z��:j=@��Q��<Rs������IZ=C�e���Ud��<-��<si�ɼJ��4=:Pt=�3��=@��<�� =�v�;e�����;ݚF=Dx�K�Z=7 ��f�W=ظ!��?����hn�6z =���<T�<Zֆ�M�;�V"�		�~p9k�<}j<��ļˍ�<Eq�*�l�E�o��C�Q���ʼ�����4�`��<�B=�*�=���<��/=��4�	�����r��<��)=|l|�{_漿TZ=���;��o=NT�<�+��d��<�O�<%AF<�P@������;��	=�=xu�{㾼���U��;�Ur=�<���ݗ��P?<t��<�W;��6=b����j�?��<3�h������?�X$=u�m�cY=yd�<[O=+���{�B��]��l�F=�L�m��	��FC��r�0�=KO�)=�9�a�<��=7$=ϻ� ���
=U!w<�jB=Q8�LE߼A�^=	���>���!X�c8�<` �+M�Gؖ<B)?<�4�<��=�Œ��H#���u=��9����<\�U�lm�d,p;&���C����E3/=%m>=��O{d;�f�=S�9n���������=� =�E�0�km.=��/=n8t=�=0v6�A4<�]üBG3=��<�&=}f\��na9;�<�F=��7=u��D����;����b<=�>f<K=��D�=����Z��<�`�<���<�:Q="�:=��D=G,���=q��<[�9�CH=^��<d"�'��;B7`��t=�0�<��⼬*�s��O��<��^<�L�<�����;��D	=$�<�ly�3�w�#D='��=�ȼp��=s���a`=c�S��� <�o �+�'���${�&q=��0=1�����"=�ZV=�&=^|�W>������}Y,�v�P=q�<��w</����J
<Ｙ;Vي�x���>6<�1=�4�<��`��4��qi�04O�	]�;������aE&����<��.=R4�<�
��|𼕗n=�qA�b�6�/$�<zmO��t��i�<�\���:=l;��"=��L=�ͼr�<z�.=�`���}��ݫ<�.��ex���f�w�Px=��=��޼�b����6=
��+W��!�2��=@�
="i��=<�&!�k�Z:��
=N�����=��߇]��g��j �=�@I���<�	�U�x�Иf<�@
=��μ���%=�����'����J���=�Ǘ<F�G=}i�i�B<�PƼ�c���k̼����� �Ø�<��J�D<��3�"=K6��/�n`�<ʏ<a�;	n_���F�A[��҆<b�/�|c����]��׬<��=��7=�%��/B���(;f|߼�>=�Fm��u��=0����=�:+=��o=$�ڼg�=tl�<t:-��mv=|� =�<=��;�34�7�<}?�Sj4=�Nn<v�<8�R�V�ۼ�e������<y��<�޼Uf=�.�y�<�������<>�=�U"<ZJ8��V���.<�$�<�X@���p=o�^=�����]�;S�`=�ڻ��>=��=�/���9��\=��ź�8���==@r׻_M�<��?�.,꼨f^�[��͆&=љ:�=�F��=�B�����׎6���<��a=�>��G���Y=!�wrX=�m=;�=�W<� u=��F�>��Q�!B%=�_���Ƽ|���;;8\��g�<�;=�m:;\�:��{��!\=jK�</v<X6ܻ�=�vc�
�'��1E�S�;�5l=&w=�������E@�<��4�+�d��9���T8���X=��X7�d�9��*\<���F<c��;U0�^ʹ<g�;��<���:2U0�L�{���ͼQ�M=�g7=�D:�;h<<���;�ʼ)CG=�r���<	�<��`��c<k�N=J�=EX��Z*i<a<o=e�<Am=�T<�ɵ���c;T�<�Q=R	:<N<��`=�p=ֿS=���R p�zm��5y:=A�T�Џ
�s�K=iC��:;����:�p<p�M�����N<L��J��<��`=�y�`��<��H�W�"�����n<���=��,�N�j�kP��z;�K�h��JR=��n���.=M�+��H��BB=��={j�;jS=�a���</���M���u�ZF�<�L=gv��[���Y<8����9�h=<����5=���<}1H<+�;�.F�C����"M¼��~<���<4�üF�n���G���n�B��sG��5�)<�����缂
F�D�2��=��5��I����J��e]=��R���4��b`�.=�V:�>2��*�]'=h��<{V����;�N����<v>�U�#�?�Ɩ`=��<;^?�=��;��<8�i�&!�<��=�Fd�%�����g5��V=�NT�����x�<��(=CG�A�Ἳ5�<��8��;��7=��	�{�#���R;%�T�[`;<Mo<��8=��<3��C����[�/�==�E<rVY��� �L��<8�N�_�X���^=	<��E��/#=��.=���L9���I=V�T=�<TQ'=XC�F1���Z�&<�q��:���d�'�=����<�O==��Ҽ��8��]��׵a�ݮ<�q�<��U���<=�O<��;���7��n=9⋻ފ;SU=�*Ǽd-H���n�==%+�:^9�Q�4q#�!�ܼ��'�o�e�W;�n�����u=�=ϙ_�{�3=�証%jw<���<Ą�<s��ڕ��O���aa=�T#=$���گ=u�=7�{=|�`� ѧ����<��w��
�<��w�}��<4�=6U��R�ƻs�(=7k=m�=�7^=���J��<�f��-�`(f<�8c<'fW������7�=�s=�&�<6-<��~}�<2��<A5�<=YW���"=B��Oߜ<\���=�c<4��<v�h�C;��^=�ch��r��L>{<�L��x�Q�hL]=�V�jH=��Y= [��C;�NzY<�,=��B=F�<�{T=�p�������<<��Or=���q=�dż�"l��4���=��+=&c=sR���R=y��������û�v��:u�xY��.�<�V<��;��;��\|<iԵ;(��<�w�<�Z�<�G�F��<!�켇g�9i���X�M���=�7	<�ۏ<�1�s�w=��>�T��e7-=�D�)ܗ�%L�=�lJ=q�O�>�)�3Aɼbo��D]x<��	<3g��,=��g<�m�<�5M��=xK�;Q�7�>��;+�=��r=c<{h ��FM��ۼh��<�-�<:@=]�H=?����)=�9Ѽ�c=j`f�lR��J�;����IC�LS[;�O�<�[��zG='E4;��'=����QV)��h=cg�<�����a<��<!S��d]�<��Z=4�G�6YL��k����<ɤ�7]���=:��Z�$�H��=x:2��;!�⻆G��R=uN==�]��q0=���<�V�<)%���N=3�f�Ϲ�c|A<��=:^�<�����18="?<�+��H��<��0��q0��M����<��r<����s�k=�,���8	�X=��5��l$�Z�H=�0�J�u���E�s�=��(=�0�;�><SEh<���<�}�v ����G��U=ڃ�<����I����J=�k%�k�F<�W�<�oC��#+:��<6�_=�<c��:�K^<d�=k�f���n�v�)��'���1�2�<�A����I���߄=�=��(<��E�ꂼ�8��'׻�=�;�<��T�i�=�W�;]�ռl\�<��<�z=��v
��Q'>�_��;F��<:�<��Լ}�j;�Hx=5��<�(��*φ<)�	�E��;�WM�9*�<�-4��3!��NI=�8�	0ϼ�pݼ"����IT����.=����_� ��T9�Nx=���p�ya=5]�<�I'<�7=z%0�q~�9��n�Em�����+�P��"��Զ;�53=⍈��S=̷=�"q<Ә1���U�9= �g:�J�<���:��5���=�k�@���v=N�ںQ�h���$�=����<���n�(=u[�<�e޼�[h��,=�� =�U�<�<�[���<��"=�U���n�Ҿ5=�D�:��=�L =4�E���<�(=�yc<�=����|�.=�6�CϹ��� ��.��4^=��<ݩ��Ӵ��z��%=]	)���-�S�p�d�"E�;��D���G���O=cd�;&��<��l�HSY��,=^5�,v3�)=ɗ�<���;�-=��<�T�<�wK����%��I�����i����=7c�<�=^���r�r��C���LZ=;D,�Js�s=�+�<����B�8�E=f��o�v�	H�f>
��A=ă=1����u)��9x�%@b=������D���켋��<\Z/<l{%<�z�;��L�<lvټ]�4��|ɼ(�<���<��ܼ `={��;Q����1s<�D�<�<��T���<^�@=�o��Zn<2�]��:���: R"�m�;3"�</F޼x�d;N]=j�R=��Q�p�=��J;�"1<��[V�<<v=꩟��c)=��D�ABO���3� ��m�稼�8��w|߻{2�ts������M=��߼L���仾��;���P�:U��;�#�W%=��9��<�㼇@Ǻ�!]���b�\��<��~��_B=8a�<)U8��9L=V�5��(=�s`�������<[�K�/�\�f=�<�E���V�<�}�< �Y�-�E������u�L(=��$<��n<yg�<Z~��r�s=�A+��;M�f��/=ֻR=R�<_,@�|���CP=��<�1=���α�;'P=�~\=��t����<�n�<������e�ۤ2=�-<;�0B=�FS�,��<i�=U=l+�e�n�Z'�<,���?�B�CGϼ� ,=J��<�z�<I�m=q`<h=ﹷ<��M=qO�<��D=O��L�����<��<߄��v�0;�U=X�X��7��=�v�<��O�:+�)��8�$�<����1��؜U=՞(����<=i����<"���==8���<\��;m��<*�z��ʥ��('<��S=C���F�B�(h�̵=�j~</�H��[&=���9�X<
M=��<�^=��L�-�ͼ���</>I=U\.�T�ͼ����?�ּ�ZR��=��F=<�N_�,.<�]�����:���<F�����<���0k���7=a^	;���<�Z��X�<�:=��<��u���w<5M=�"=�p��AL$�l�,=?�Z��?�<I=�:��)6=��T��k�<Q�Y=��=��|��	�S��+������ �=s?#=�TD=���,�<�6�
�@�����)�=�b����<)RL<���<��=�Q`���k��<g[�<I��<�M@� L"�*�1��F��n=K�*،;W-��<rͻ��
;����ب:�06�T�;={H<=~dj�'[=�[��@pY�(ź���<IC��^J<�c<�];u�<��<�=�ަ<e�8=Bb=�$=E>l����<��	��/%=S��<��<M@=Y}�<�r���=׀0=�V<irB=:M49d��<��c��P;I%=O	5=.<@�J4O=KC���<^�G=n=˼�=:H���ݼϏZ=pG%=���'.%=@�=�6R�(�.=��TM=n|/=5�$=?��< �j=va�<{t�j,'=��Y=]�=/(�<�y`��w����0��<j15/b�;�҃=�y��j=���;�ϼi����%��MT�7�0=z����<�=�/9=մn=k�W=iH6=�@�dW4��>�<�&����j�_���u=ݠ8�E�����=y��< (�<�q�<���<���<�6=<��X=�bx; {C����� .=-��ǁ�<�S���/=��<t�;����<�<ڼ9��"�=��˼7I�<k��<c�ȻJ2w�f�=ʼ��U=@]=�U�V�^;��0=�����}=iCs�Y*�;�Y�<k智!7;���<��sF�<��<e4�(2<[}��/-�yT�<%�=�\q�X�=x#��{�;�u�<y��<�a	��<�%f���g��̼�c=�»���<��=3�(�EL6<�+b�1�<���d=�d�=v�=�x=��ǻ*�����$<�y��O��<�K�&�1��*�~�:;Tx�ޚ=��3�u�0� H��I0=�C�'=�V =j���Q��w;�nw�{���D�t=��r���O���<��={�<� �<_\���6�P�r�>��P�J=XO�e�I=y;="GZ<���;����\=���<�t5<>3=�=��E��f"=ϻ�S=��;����^i���4V�6�)<_�<mk��b�<�Ӌ<�
�EC����h����;�ݼ��2���<U�ϼi�����C=~O=�n�<�4��U=� �<x=�C;̕1��?=���;���<3R�<@h}��=&���}�7�7;̲i��kU�0=���3���o55��fF=�r�m-%=�_��tM<b�<p$����5��'����<e�-=�l<<ã���;�:=�ҺB�=����Z=ͽ��T��F�<��==¼"�B�dO4��h}<Ȅ�lx,�a�E�+�'=���<�K�_��=�X<�B�����f	��O�z����	���W(=&H�<T�F=��6=^G4=H`d��@I=l?0���1=�J=eJλX����缛���C��������<�N�tS*�=p�*=�=;�� �B=�R=��A;���l< ����f��;��t�c<$㒼j�F=���<N5K=l��<���:i@��޻�3J���n���N<�ϻa"=��	;�����=}�"���<X���4ͼ�<�`�<��4�4����=��p��n�<L�=��D=>�*=���u�=�Lf<�(}�`3=-����F��sx��z=nꃽ��=p�p=�R='�A==ü��Q=�|�}=�f< �=��P�1��<���<r���Ζ�j�1�>T��O�%=��<t��<�-J=�T95e<�B=�4L�[����]=X;��ΎH<��n=c�Y��i=���A�<YNU=�x	�ڏ<�g
��m<3kr��Ԏ<���<Y�0<��	�ƣ�2�r���=����A:=DDo�MD��=͔K��=����A�;����$���B�<�I�ظ;�@�S���U=��<�{��k_=��(<���=�]@=g-�;�ng<~V�:7
�;T�<f�U=�u�����c�;85�<mPk��߆<�,�R�ؼ�=xw�<r��;Ec�<��u�h>n�ѺP<Z9X�o��,V����)<_�x�����5�I��^�LC��l3�|�=Sh�NuD=,�=��$<& �o�� 6;c5 =��u��Z
=��\=��C=��;�;q=�Ջ;(�q<�!�<V� �(�ܦ�<�V�����/I;=�J��"��I<D&7<*�[��@'�5�C<3�����</�=x@7=Ê��k=	<u�r5�or����:N;<�ϻE�$�"�����V��`��C5��a/�M�c�md�<�Y�< �{= v�=T�N~i�WD�t�F�"@{;��/<��h=!��<'2i�B�d5=Qdһ{��c�v�$w�=��*=�!=���;�
Y\=�U_<$�[�THM�1p���;�� >�=੼Z�N<(=���5��(�[�S=V|=�n߼8�#��@1�p7��EO=�):;/$�<Q_�:�\�l����� ����;G���?�0�<!y<��	Z�����<���Be'�3O@=�Ā��e%��gY=V�N��B=���<oQ4��,	=1�;���=K/D�MM�[�Y=�� �����R�����۬�����_�r��=-,�>�ּ*AW�����k�=$gG;�Fp�"���D���s;Kۢ:F�-=&��K�b��"�3z�n�=)�i=?�N=��0�Χ�Nd��DPk=\���� �/�&�r;�R�<�gy� F�<�=g�1=��6=MT�>�*���<��v�ѩ=.#�<�o|���e�jƸ<I6�MR���C==�D��;�,���z��<h�a�����`@��<�}�-��<ݬ�n	=f.=nhI�Zx ��
�޺<� �:Ҿ�<�+껏�9<#�4��?�=~�ϼ���c'ż!��N�p��oO�jN�������:�����
���1=�3໤��<���;8y鼡�!����;t��<����򐼶����;W���b=h�=�ʼƦ6�\f;����5�=�a�z���=^��s�P=��<���<Y�=��[=U��<�K`=U޼H1A=�]�:4ق;�|�CD5���#����<���<	�<-5=:������0����b�p<X�<�&������R��=��?;[�;��\<ML�!ܺ<~9K�bI��\.#=9��f�s=�HE��[�<������D��~�pL(=�H���@=��=�_
��Rv====bD�<ؙe=g�;�I�8=a��C��<�z'�b�|�l��;3=X�M=1��'�m=;�R=$��I:R���x�b=b�5<u����|���Q�$㷼���<׮<L��:Kx0�7#�<��x=|�M<����e"<$V�<?T�<X��;E+�=h�$<��=n/A���)Ć<&���,�D��<�I��==��0=3l��p�Z=��L=�Y#����k�C���������P����;�B==Q:��i.< =ۗ�<D�μ5L=>&;�憽�����@�a�]����;��M=�w�<�/?�-U=��.=�x
=M]��Vw�P�:gL�<�o)�r�<w����@�<I I=8U>����<��:�l�;>8�'��;,�y<�a:�=�"=�:�
�;��=q_n=��;��ͼ�]����ټ3R�<2�;���IO��e��<S��;��=��ct�&�<��&��<w~=p�0��AἚm3������'<=0/.�6�Ѽ�yF=����`]=T��e�~<�� =�h�=��V� "=�i����=�Qm�\�w<a�,6=��d=�Ig��z��+=��=0AL=�3<���<�rz�P a=�ef9²^=��'<�0�Hh�c�(yR= �~��	I;eA2=�OU=v�:<��>=��Q=��.�{=;�M;� ~�����	.�ٕn<��<��ȼ�&�qک�X��2)��*�x�"�:��7�;3�L=��ü��8=	�=���<l�滩�=��
��
7����w���u<�za�7��FWT<��z<�M;�1�z1	�IB/�#�<��I<���<�ɜ���/���1���μ�+z=�E�<ݹ8������'=>/'�<4K��B)��s\���<�`�==�l=�K�<�|4��'���);����<��=c#=ē)��c��Vy_=�֌��o�<֍��~�R��f���ǉ;_:�W�=�E==	�hw���<I	\<4��/T1=�^�;f༬(�<���:�F�9s�0�4 =�V(�B!=˒���\>��仔'�<�3���c=�[�<��<���<"�^��|x=j�<�Q��� =�0��6��<�Nͼ1G�4?=��0=�ŝ< y=n�^=�
@=3I@=��$7�<��!=�gj=�%X�?9�;��.=醯�֧"=E�f�H1�<�;�=4��K�5�)I{<�L�:���4H߼+3]�Q��<<��<�]�n	�<t,���vG=����>:�u�B�X��<k�:f�w�)��$-=9���4�+<�>A�.�S=�4<Ҩ3�N�=#����D�\���{=�L��e=Pa�$��h�j�l<W��<�چ=��=�����_?��Ϸ�=t60���#�\��<���"=>Q�;�*=�K��=����W��'l)�1�>X����C�>�!F=xb'�L�:=v�<�;�{+=[3<�^m=�Lr�kT�9�o"=������;��z��6O=�O�<�?�<ԙQ=1�����<p>8;9�5=����H� =H-"=�f+=�wb���=��&��$^=$)�$��<�`+=�E:=��=N���_�<Q��<��c�k�	�`5��6�;u�@�\����S;���(�<���<�b=ש=�H�����<g�);�L�!*=á#=ݣ��#�^���,��P;=�Y=�S�<�2�B�Z�D�W��:�]T#=-Z�;�
�<��)�2o=鿸�H��<�m�p�;Bf�t�X=�!;i��9Z�<��;�p<#�c�z�Q�Ԛ�<�O�;�鹼�����ɘ<�
*�bN�<[!��v)==3B+��iZ=oI�<%�;=E�D<1�:��.<����E�<*�<�&�՛���=����6��K8=n2@��<�C����<g꫼���<��Y=���U�<��[=گƼ�=p�ԼAu��Ò��3ռe_�;��=d�B�̀ƻcW�;`ƃ<�@ ��*� T(=~�o�>�?=VC`<5B�DE�D��<;�M=d�0�������<�Z���/=bv��;5=��6�Θ���G��ps<&tF=U����$?��w)���E<�o�q�<V|%=�>��D=�o=��=�=�tB�&w�<+)@=i��<�X6��~*��v8��,�<���>�开\<l���C-#=*��:!=
PҼNX<�L��&��˼w=�v�"��.m:,�?:��"��.=!�=�81=�1=��!��=Ɋ<p�F��"=-��<����k��J�҇p�q=���5��l�Ҽ�A���NͼϹ �c�5=l�X���:<����x��;߀=k��< j2=�� <��%��k�� =묂�Of�:�1L=�?�)�����x=�5,��<������0�<�?���uY=#t.=@y.���Ǧ�:��}���`�k���E=�k=�A�<6�P��/�R�Y;�NüD�v=LGW=�F�&c��Xؼ���=��H='�MV�:F�<;��<�~'<}A�kAP=�V���LY=$�n��1<�����V=L�;��$�C=/`H=� ����p=Y�P=&򖼥8%�wO&=�� ���<�<q=�v#;O�<oz���{=��=�RL=�x�:��v;��P=~n=�['={���<,�� =<�M<4��<��(�QA����=� �<�p� Ox�`��<ieκ.�;�u4=��5�(E1���u��Z!=�=R=��U��G=��%=���X���x�����#����ח��Mr�;ϡ<m�z<�&=F��eQ��.�Q;[=�DF��ѻm�,=��H��<����˃�X�:�-P=�
�t2*���{�<����\��L�t<V�,<9�<��P���=Is-���������r�R
<��;�<��
=N���a<,m=�e:�0���/�X�3=Ǟ=M�Rb�;w�Z=>�J���<� <�և�B*�=`�<b)m<�wk:����w\0=8w=�w���J�<�r��'V=y�n��c�z�<E���\X=Lz�<zvY��8Y�����h=�qu=}1�;�>��sU=�Q����%�a�~�2T4=�%���O��>�;�I��ĸ�����h���{��(�%�b<Z�ʼ�~�<9G��#�;ߛ�<.�D=F�<��{=��o�.�!��OS�� ,=�J��e�<���;��9=��R=�eX��~�<�	�H���ټ��R��ρ=^��<?�0Al���:�=�>)=D�8=��7���==���v2=P�'=4�7����AT����<,�p��K <5���#����L>���@<�2�zDɼ��<��
��B	<�0�{���H�Q=</=�}���J��0 U��p�tU=%7,;���w5�c�<��缇��<^�o�d��<�	:�	��`�3=��<!TR<�B�<'׼�!L�����V��3�<�(k=��<� +�$'<�C�=K�̼��<��K����o���� G����<� �;ĕF<P�:��R������4���[=�#�[z8=3�)=˨D�i�����<��	=����Dr=�8��)\�_���h��)�=S�4=g�*=�H�B��<W�>�G���	;�g���?E<�E;=%+�<=�t�.-��M=Q���6f)���M=o�e=��<�V�H��<��m=o��<�s��q=E5�<?� =�܇�S��<�R�	<�<9�<1n�;���;���c��?!ļ���=�x�<��K�ԡJ���<�矼�i��Vż=��2=_�k��l����<�;!,n=d���b�<w���A�ق|�@�;� =o�=�J�<�
<�Jr����<gjA��<[=������%<��<�@����<���l�<��;���<��=��Q<�Xn�Y5=�%<.<9�X3=Rk��x<�KD��A̼S @=n3=��<i��:&!E=$H<`R3=��K��莽f�»}���{�Z�M�T:��W�J�<F�v<�)�U1�m�=�B��1��F��X�3=��;�S<�F��<'k����S<�$��V`�0U=gV�=���Q_#=�[1<]ep�Jn<:'x��%��4G�FHw=p�»C`7��x<��
�Y�W���[<���ͯN=�UM<�	#=�J�����<�B7�
�G<i��<��k��?�.r{��h��{*=�s/��5	�?W]=��K<q<NS�<�Sx���%<8X�<U�r<��}<�-�<��7=����z�2=^��������+�FC=��h<��=1�;��J�Yd<E~=�v���\�<�sS���!=�6,=�Uؼ����j����g�[Dֺ���(kƺ>�	<���<��="㪼�A�<!�==���'f<�$T=e(�퓼���_�h����Zo�Z���=*?`=!>%=N����l�Ƕ9�C�==ɼW=��
�[�%<�~=�2F<��>�zo��y	=jGC=�=� 5=��;nq�<g� �yi�����YF=��%�9���eü��=j���H�nɨ���<��K;�C���>_���E�!=�WK=�E�;�9��ujD�w�ռ�����O=�^���/�*��:k�ռ�э=��<�=��:�]Rg�O`̼]6�<1�j;,�=��P=�<���)G�<��/;�Č�+t<�o��ৼAW=˗�<Jp������1=-�T=:�w�y%�;$,�<�Q=��ƼJ�<W8V=�W=G2=�3� _a=��ټ��B���K=�g�̺u=�#v=��<�r�<_�=�>ƻ�K���V� �z�_�P��<\�>f��&�n���f/��,�_�=�.�}����<`^�<�X>= ��<��&��k`���`;S=�=�>=�<?�Q=GJ���{�<�t���+3=���<��l=Q�F=MX����a���=�U��V`���b=6�;��$�
�Ƽ��5�����tFs<�q�}; =$��
G�<x<A�"=��v<�b	����<�Gż���_BV<'�(A=;�x=v/8�+��<�k�̊=H��=������X�<����~<��(�b���{=�/=W�O=y6J���Ӽ���<[�B����<W�5�gQQ�2�����i
y<�^=p��}A�<���;�s�'(C�.e7�X�޼�{�.�C=���՜2=.̼��<y7���)=a��/m�D�<=`<(=uS�;��>���ʼK��#H=�滻y�=*�;g���+=�����Yu���EF���$<�;����>�N=.;��_��\$}=�3D=�ҷ�z�<�b<�(<�4ƻ�Aq=I8�4���Ĺ���/���+<EK��̄�r��<�g�(���/E���	=�W=f�;Զ޼.<�<SP��"�n�0!��<�l�;	ۻ�q=.q�,M#��ȇ��:�=Z�/���=~����Z�{e���v>=̻�عZ=��v=^z��,I<�]=���<]Q�<������_��߶<�� $<�,=@�l�{�!��*M=xN�Iͳ<X�������=٪��AwT8��}��;µӼ8��<J�#��3t�k��;�:=���&���!=�ǳ<k�=A����ۺ���N��<c%�;�%=8C�<잼��<z���(<ͻ=&
<�;��ú�Af�׫%=�F:���[�X=�Y�:� �;�M=iM�1�=43ں�=|�;�"&=�R��������b�<
U<G�=0d�O�=w����f�<�H=ٲ��A����)<�~�=����:��a=`�(=�J=xE=���Inʻ_�=k�<7o��_l�_��<�;x<��B=��?;Zb=샽��W��9=��y=�|�;K"��h�Y��Q�9�N�; 	����<��=�{�;�
.=�G;�#�<�G����{?� /�[�������T��5X��~���̝�F��<�l�9�el;Ԧ=��@=-�q<�/=�z���:�#=� .���;c�=h_T=���9Ho�<Y�/�/=��C;��)�ͬ
=?�S<!^���;��J.?��s"=�Q=G�p<.S=��9�z�U����<y�O=h�<�-���B���%;�1�<`)�:d�ؼ�F�(�;�t!����<���+�t�s􎼁.����<�(�<��4�W.C�wG=�*�I���|�<��*���ͼ, ����*��=v<U����+;���<�μzX<����/	=L|�z�l�V=��"�: ������H=���<�h�<a۝<5� =�>���޺;���=ͦ7��q����Q���?=�3�l�^��.#�l�=Q�2�,�;��K��ֳ=Z�ڻd^����p;�z��T�@=�,=�T=ɚ&�m�6�y��)=�)�e�A=��=��
��?�<Ő3�g�4��"���X�?<��/�̕�<�d<�7���c<;�W���ح=˂>=�=���gD�2=�,o<9M:;k���W����9`�릇;~��Ҳ�"Qi�v�"���:F��<��
�ѳ==b�����n�;���~�B=b�Ｗg�;�q���C<5�w�B�:=Q��<G-<�xI�ᕊ��4=�}�[j�<��~=a�7=���<��|<ғN���Y;��<���;��ռ�(�v��;�=wG�<���<^#��o��mT�>�e��Gӻи���_��hR��x%�4�g�\����^=!t=��?<=C�s·�J[s��x=#��<r��@��\-��3R<DμX}�</��<O@��4&F:\c,��IռN���c:���,��u��ܼo��<#07�[eZ;:/^=�t$;S��5>N=��3����Pu0�<�}��5O;b��<ϫ =�n����<�Dܼ�J��AT=��F��,K<N��1�<B�G�
�w��K����;4����s=&�d�:82=x>���I=�*�;��=.&�<��;��=k7�<4h$=8���$C={�ow�<>����y�)�;>Y�<�0g�Õo��<���<���k-�<7_=��; !K=�ܛ���=���s����Ç<lI-;��j�}�R=���7���f�;:%=���<�-��J�<1;|�;�,�.P�<�/y<J�4���<����8�;5� ��=��A�t&��_���Z;Qvμ �<=;���mr�<�F�S���̼<����b=�4-i�M Y=�K��L�e���6̞<7мP�;�-=a�)��4�-�R;��?��ȹ��'f��A9�Q��<HdX:��b���*�s`Q�+`a=�1|=�i��Y<jŰ�X@���i�<I��<�)�Q"�,t��#"=��&=���?Co�͝%��Yܼ;�W;|[��f�<�Y�<\��<H))�ʭ�w/�<��<�r�;����.�����89�=�Q�|#�;b"s�>�%=H'�v��c�O=�s=����2~�<_�1�GS�<c���pB=�v��8<�=��P�#��<tl�<�;�,?=�x=h*8�5�<�I4=H=W=�w���y�;�)?=��@5;B�H�~�������z<�Z=�JH=JL=Y^	�Bl��u����l=�>c<�I�<�W�<��=��;1��<8:"=x����<��P=L�K=Yga�����Z4*�@�ɞ*�v��1s��ွ0gI=�<���]�U=�t<��=��A��6=����o��<�Dؼ��f�8`<��X=�=��f�I�&��i�<�ͨ�a���@=�I7���U=J�<�,�=�Wݼ
�<ͳ>�Xż31��g�<G��H{��:!�K�m;������Q=g�N�.��m�c��k-���X�0ؙ<x�����H==�="����#L
=2�i<0�<��q�[!<�I��~����E���Z�A��'�<]I=����¹�_�������]]��Tq=A�	=���y�,;==�IϜ:��=P2"�5{F=����!=����;Lr�<��&<�=���<6��F/=�<�'��)o< 4����U��s�<�<$X=�==V������<��;jb����(�P�J=Í�ׂT=n^M���8=Yzs��F<�3����<@���'����%ڻ^4Z�De<�x�%:8��û��A�LU��ru�<��<�*,=jXټ�P=W/�K��<��8�x�=��U<y�/��v4=iqż�����N=�j;T��;���#<���a~��@�^=0w��3Zܼ�j��\7ͼ�=�={�=�3`=��^=�3G=�i8=��Q�Ȟz����;x>�5Y�""=/�<����:��^�T8Q<;�h�=�+ռ�8�<U�><��T=�h�z�_�C-|=�"�;ǎ�j}��_�"�FM=�Q�:�*Ǽ)�5��x�D)7=F=��<=n��s�=l�0���{�c�<'73=��=y�~=��`=��=5��<n;~=�l<
�I�s�=A[=����Y�b=v?<F��4��~_��Q�R�n��m5)��n<��?<I����)�<}��T?��c=�����V =#�j;��L=��"��fK�#��=�kȻ�"}���H��L�<�	v���<I�=@��e=[�+<�q��g��H=������1=���<
�=� M=@�ϼ���*/4=��b=��O�P[#����<.(��Yt�ײe�F�ne=�Q�^3=o���<|���=�d��K�<��%<d�(��#=[8=���<��= ��FC�<w�����t��<m�=qg'=���gӅ<�@-=#0���w��=�q�C�ӺB��#y�ջ@=-=ʇD�?��<��k��#U=t
<�
/=q�V�p(
<�L�<#�
=�v^�+�>��	?�g%1=�9�#��<�Z��qQ�-�d=��=*x=��}��B3� 1=��=_�I=�wü���<�/�9�;�+=����Rc����/=�z=�;�,"��!r=(<�=q=1�x<�.;�� <N��<�M;�;�;��8��Xb�J��<�a`=1l�'� ��>�<��V�^����=��*��Dz=$��;��f<�e�=�t<���=�f=���<�L=�6=��W=�x#��)�<�<���;���<��P=6=N�\Q��fM=���K�=.�<�G�<�Q�A[A=��4��L�$�E=-�W� ҇<]�=����j�>�=h%�r�'<B�8=1K�H0-��3s9n��Hf�]=9��D��?=K�i=N�<�@<x��<8D���2#��ʹQ��<��}<�����\=J ��"����k�(d =����<A�9:K<DԿ�ȴV�rIj<�;=@Ǹ���"��
�<���<���:�2�pG�<�Y>=R?=�P�<D'�)4��c|<D����^�<9�<+	�Wع�����4%=bf��(�<8���=�H��{<�=z[i=}�&=�~=�
ܼQU��`1=Z��<m\O=	m:�,=�@=Է���= K��L�ӥ<�|=�'��	Y=�>R;��$=���	��<T��x��I=�:��R=$�ۼ��7��4>�P�Y=
��oi=���<m�=6]=I]=�O���T=t$`��d<e@5=W��<�`�w	,��c=
���@=N��K�˺C��<��X���z� MR=���<�'��c<�f�=8�;m"d=��=�]^<9W��P+�<���<�H�U =��㼤�1�㿂��ֻ��=�];��=���=������=��<Z-=����A=�q3��y(=��U��D����H�b������>l=� C���0=��7:�E(=����B��jM=>T'��#f�+�=�ϸ�A;�.�k�R9�խ=�<�<�z��%�l=6�ڼʎh�q���m�=��~��0ü���3�<��=��Z��<<��F=�G�:ƚA=~�=+Ƴ;�u�9&���c�1�޼f�!=e�$=�W<�-2=鍆�=�6<���<���<���=��<g�"=\&�<%b��>�<1��<l��<�D	=G�P��c7=�Ӽ/�`���|<Ƀ:�s=3<ZT=�q�;Fr���>'���%��b�<��*���d�}%�<�z�<�Y;-��B6�:��:Ĭ�<�b������C�b%�rK@�\W<��w
=��=!�e�,U=��<p�=�.�<��{<�)��A?L=SQ��t�<C#-:$� ��bɻ|�r<�J���d<¸�<o/��a'�~�<�V�N�q=�6=@ M����<�<��׻�Kb<��P=!��� �y�a=`��<��A�ʀ��y�<�N�*�!<��s�?�K=�3��л=q=5����@=��(���=� =���[ ���(�k�~���{�Q$}�F�4=@/ۺ��+=��<�UT=��I�:S��F=�$@=�uT����<*|�K��<����.c���H�=5�q��;=�P�:�ȩ;��<}~0=X��;;�o�]����E���nL�f_�=������Y<:H<!�+�ctX���2��9�;�i� <�!�h� =1ջ�u7�U���dg<�eιȎ�bpC=]k����<�D=��)=a]U=��9=�����6"=��P�ʹ�<�q輾�;=<i���+���=���z=�)���q��qA��)��T|�[�#vʼ���|��t�����<��;�0�;V��@Eg=�z�;N�<�H�<�=�'�<�6�E.=����U`�<���;P\���5=5=p:=���	=�� �&�5�P��;���z=Q��;����[������n<l=�0�<��¼2g"��-�<�`?����; t���}D=^�5=���4<�
+=��K�(��{�<j7.�* ���\�]��=�\�-FL=�:=��t={�����<��J���=�[��v�@M����v��Ł�Ŭ?�>�y=�lS���=�l=X&��V]=��v=��׼� �<T�A��֤<+�żV���$p =>���� ���<�7.=p�<ŀ��Z��=E:1=�;Ի�F`=id=R�P���мl3��L��<&ă=Y�j��Z5���l=��/�#�⼑�y�W]��,�=�H��7<���t(���F-=p���I�<��t��Ů<���%�2��w:=�/���<��^=��g���<�(g�m���Y�<s�<>�P=�\��B<}2�:���<�[��\5���_$�u]��������������j��6���<6N<��a����<Y��<�=���@?�<�6��3n=���<�)�<�b?=��y��@H�᥁�G�=�x�(��'�<�=d�x<r�`�0��(�<��n��WG<���<��伺[��5*=���<��H��<X�����<鼣Ā�+���<�Z�;t��{�����l<n��;\D�ę	=�	c�.˥<�j��47='��##�;��e=�y�G�t</�=O݉�HJl=ސ�<�Z=�=q��<��<7 ��b＀�M�2�=N=��(=�F��@���BZ����<T׼E?ټ��<�|-:��;5O�=���<Ԩ�;�Z=��
��D�<7OG��*�x�)=�6"�><3�G���/$5=A��<Sb�;��2��;%=d4�����9���=��i�;i03=�p<>g<�G!=�c<�	CK=�Y� �S��Á=�YS�da.=;��}��v����<O��֋�K_�<O�:����#U�<~&B���<���<gmû�v�<��V=#�����H�;UF���� =>�G	ļ�q����U=O�3=@#�0d���?�e���Fj=w4]���F=�=YS�<Pȼ^��;[������9;c]<螺>>�<\|<tIH�Ý��y�;��<W����F=��ػC�=a�Ѽ/�<��=,֊<���n�<�¬<��*��
=��^=������g��<< �<�q�t���Fш=㌮;��J���=o+=4_:�.�;nA�n��,�}���:����)�<�l7=2�ߺָ�<��<q<��==����>��^��
BJ=������=�/6�!��nf2��V�<��=�A�<W�:�ʙ==�ـ�3�q<oN�=T�����<z���z�;]U_==�R�<�P=�G⼱N��p�<��U=p~�0G <�����=�/ɼ�"�<�i<Q�[=+%"=8�=����ax��b_�:����(=���<�>�W�D>j�+��=~�<��>=�f/=�V��u6_=��<�V�����<���:0p�<<=�oJ�7Z<1�<��<<���o��L=�k=�<��Q���O=��=�.(=�ȳ���{<�m<_⃽W�=�=�U�:~Ԭ<W<l:��� ǻf�~�����~y=zL��SY�@���n�A���z��q�ޤR=0��<�=L�μ��^=���o��$�<�[_��h<�_��b��<�s0=�v=��5;�����R=�g=`�����*�M= �.���0=�.f<\��V�e=�G:�^F�͇V=��X={!r���=�����<�@�� �<�K���4��64
=V<�(��n��,���=�+���?����:-�:��B��ޫ��k��k-=�D�����<J:=��#���ֻ�H=�|=�<q;���<�P���,�y|6=�b=�<y<�Jr�;[�;��<E�������<�Q<��)��A�;P>=��8_=(>%=�t=z�'��=-'�;ܪ��D��<?��<�u�<�4H=��[:n��D�<��@v�$7��ad��0X=����G=�%=H�==��;Tߩ<������&<��o=9�6���-<`j =O��;H�'=��+=�e�<�H��΂]=b�=��V����ǖ���=p��H��W`=LH���1=�%D=��<Z���as�<���:y�=�N��t���4�*=��;u=u��<�Y���{;�z|;�����U�<�Ӌ���<L*=�b=y�<�o�yz�<K�m�k=ɤ�<Hw�������y;Ӽ,�$��-.<pJ =5��vH:<��N��h��)fW=���<�uȻn =���}T;Rf�;Q���-d�y�ӻŏ��/��<}�z��=o�z<�U<�yv<زR�e`��d3'=���<�=3=*�'="a=�$�<�����û�2R�oj/������>=f9�;֐@���y<���<4QA=�X�:ZO��v��N�==��;������<�<��7��<'Aռ���;9�󼸓�<|d���y=�#6<s)y�h<�"<��I=��6�<}=>� =dD<�ռt?<�GR��a��cq<l^Լr�/=Ų���!���|<����|==�$c=��>��'�=q�(�Y'�<j�R�'8���8��_�<S��χ=�ϼ��9�Hn(=�2z;�����*D���.��$̺Fz�<|7�����r�E=��<��:����[�Z=���ѼF�<Ah���'�e0���]]=	�
�[&���|�~�<��<GW6�#)#=C�����'�gS=�<�<���<��=8)(=�&�<r�<�^-=�Te=i?7<�P�<O�S���<��ﻱN���Dq�A����9���*=�C*
=������<���ڦ;Dff�l�<�>�a�k=s5<=�=�� <��� �/=��#��*t�����6ͼj����=����"�.�R=}D���D��i�;U=�<YV� �<���<E����4���1=�Pp=�*T�GA���0="�» �U���.�<<�C�;b�9<���=���e�lI�<^7�� ���s=��<��(��[c=O/�dؼŶs:���<TF;��<�(���Z=���<��<��
;ѳQ=��;<}%=k��H/&=��%=GE���m�2*�<�ѿ����3�:E�����p?g<�5=�$X���\�ѕ_�\�y=_< P<��Y=o�=��0=�����\�O�!��2=b�=��"��y��A��X�����<G&�<ir�hH:=�3*�K�<�����8��~�T�>� ��BżN�m<a��;}��e�;����j�u���|��,6��B���x����xм+��V �;����=�1�?���q9{�������������<�!����<���<֩i���z�6*��k�Ӽ�cA=`�|;ͭ��֠�����<]����k���ɖ�"�;L'����O=��c='S<Q�<�	W�E?N=��=���V��F>����;@M`=�c=X�a=�\�b+��p����+��4
<F��������ʼ��=���<�%����;"=�K�VS=�j)��85���<R�7�[Wm���h=qr���S=�:D<�c�<V.�<C<�<k�)=��==&⪻�F�[*^=�����Ҽ��&�����U�<��c<[�<�{y.="������<1�<���R徼��;k��<q���̎=��
=D<=�q���f5=ý�GM�<.�m=��\k1����\�V�8��<�3C�Rr�:4� =�U�-o=��<�ߍ���J���k=�y=���5T=�
Y�ƃ�<��_��Z=�?g�������ȼ���A�<`��;�X�=]��/S\< 	=@�]=� ����%3=!��Up{��u1;
[�����yG����<є�<��(�CU�B�J=��<���<�FW�ǥ
�73�<9�M<�^A���4=�ޓ<&f~�/�e=#ƃ������;�%W<	z�x�A=|C�<�#t���<��=�y
��T==��=ށ�<���;�W~�GB�<3��,v=O��;5����x<��;�cX8<�ጼ����?�,@=<�WR<{��;ܭػ�{��Ύ���;Ș/��R2�b,�<c�#;����[=ҽ���Ӽ���%y�<fv=��u=5�G���	�oZ�<��<�@=H/(�'����I���=dT�<�v\=z/��y�<E �<[ꂽ�ɷ��H=L+�O_��tѺ��<�)=�s8=��'b�<�m�:�C���'t�at�6ȼ�����^��i����7�����Y<�=S��;�n�{o
=�N��!����Tϻ���<s*��e�=MMX��b���+�="����9�
I]�b�e���2=T�;��)=�`��c�H=u(K< �k=�< �¼l��9� r��._�K�K܎<�����:=�ἆ�;U��<�7���A=8���Z%<ͻ�<��^�'�b=`�<�:����;M�U���U=?�z���C;6<�D=������<W��<y�<�����w@=ha@�R�<��1�Dv<�0=����;������r=�ߕ;�>&<�>	=�I�Y�K=8�@���8��H�'9����<J�{��ut��]�����m��%\�X����P����å��;���'󍼥�5=����iS�<��n�s=x$N=4���3��=8�;e鍼�2k��+<(I/=�/�:�*C�"r����	��z�<�(�k@=���<���<��<d������Z�)<o)�hlb����,<_o-=�R�<͔�<�P�<|_��|�<U~�;�)O����<m��;�w*�����u�0�'"��R��)�=eB7=����:�<�V=��<:_�<��;=0�<v˼<W2�;.m�<['���6[������+���k<�Ț�<2��5�<c�<z�<�ב�Gݼ��gH{<� >=��!=໗����dSN=��|�1�&A�<J�<e�!9�4=^�Q�>B��A�<�9<�g���6�p�-���=0^	��_7<��g���;�=��c�MS<tC�tO�<H?=���͑���o�;g�t<^mD�|���G�ŝ;�W�<8�����<A���R =w1=V=��=�+�<ʼ<6:�
�;]߼�'=K�%=��<�zL��s'�Y�=�'������eL�|�=���<jgf=&yD�b�]=M>лH=��G<4�<~h:��9=|y2=ꦋ<u8ڼ���<H�z�s-+��:k=ޗj=6�S==������Xck�A�_�%r:;��y�j�}�&���jٻ�Br��ۨ��A=Ɍ�<Q=�TԼP�<&&��.�FG��@�=y�O�ڈ�<�#�S�u���!�2�<�XJ;�9ü *�<Lr���Y�����<��$���!��
;= zK���<�,>=g��<���<��;�nR�@�<�:=?AD=��;=��#<�H�����y*�7%�<ǫ0��~��R+��
8=�uV=l�/�,X�`p�E�H��G&�`"V=��<���<�����$�<��=�m꼩zD=�h�}��}�=U��<�;,:{&:=���<5d<�#,<�T��+�<�pI<�n2=�d������W<�Q༩�G��=�U�<	.<톑<=���D	�m���_/�<�4(=�$м�/Y<R�Y<ߡ��O�8�C�Xd�Cw�<c���t�2=�� =�:�=+��t)=��?��`�<�1ܼ2.<U���� :=ˇ�k�+=�м<1�z�,�<���<;9��QW��E$<UN=?�!<���Xܼ`3��0�v(B�q�;��=��I=��_�79=>�+=�s� z���9A��=�ȼ����/x��,�;�6���{t<|c���;�<�ۍ=��$=�ƀ=�#�<dXP�z	�WR:=e6=:==�8=v~���8�18�<�ԛ<��*��ռ6�N=��J��.����</M������`@H�\�6=�2ͻ$��=��;`�B=�W��W�;wk����;$�<P��ud|�,��zj,=�q[���:<�%�#�d=dTt��(��m"<�� =�A��7#<�u�<��;�Cu�<h~���q'�R�N��e�ȫ�f�_:}�n�y:�9�/��]�;;�ֻ�n�.rm���=��=)��f�r<�#Z��2;<���V)8�<�+=�kB:�$Լ�N�;ت=��2<M=�F�<ޘ����<���<ʍ�<�=��=o*=?8<�x�
����<fм��ټEo�<����و�=��_���!�d<q�=�<��!=�V*���=��c<5UG�נ=�S7����<Xqg<�����G<������h=�o�ܲ3<���0��u�W;g�<ƹ=D�¼Bxy=fH=8�=�7A=���<k/:�z����ay=!�<�"@�d ��c0�%�=�o(;�L=B5�=����~' </EL��,�]Q={$û��� �<�Ax�:�J=?>=`*=�g9=�ʇ=��Xώ�AJ����s�Q��u=��<����[=���Bsh=-Q�q�<�/=�B�q���B=ֲ � PH����g;`�C�;����pUӼ��E=y^���Ҽ��y=�m)=�*_��bB<AO(�5K�d������F�x�=��=��]��}1=6�2���<=*A��=�w�����+�&��1���QF��2��4���p�>h=,+��D=V��<л<:�<B�x<G9���^<�z-<����<"��i;������9<IVQ=�y�-pF=��X��4=�Gq�;B���Ľ<�U���~H��+=��o<��)=�$`�́����ػ�����="Mw<8}�<�^�j%q���1=,-=�*=�Ǟ;��=g�b�˱
��$<��|��1�;��4�]X�����<�O<0g�<뢆=�}�<�#�'	U���=�[�;��r��z%<��Q��b��~D�5��˘������I��	�=Br�<*�=`K����;�w_=��_���!��3=�{Q<��L=�A�<g��<b�[=d��<d%���W�wN=e��<�K���/�����H�<�!6<�q%;/�=Y =�ˌ�ٳ;P���0�漉(x=�fQ<q�;� ^�L��yЊ���P=�CU���l��q�U�0=�wx���I=Ң;c��;�������뻇[=���������8=:%W=�KZ�{^=g<��?��������f}�</�=����z�$<�~�����<άb���<d������D��=gU!���<j�=.��<$�.��	7�d	����<�
3=<G�<�
b�����h+�R5�;D���tݼKd��f<6�;9�<����p��<��P=�6�A�c�n	c=���.6�:��=�=(��;�Y�%E���x�:<�=ö9<T�V<�W�<���6�;8�E��U��o���I=�����j����<	�9�����v�����y�=
rB=8�-<حQ�x�<���;��i=�=�*r�A�#<W��$�|=���;6<�*�B���A��71=�+ͻq"�;�~o����T�~=r��<=jм�����-�C3�?yQ<S?A��4=/��h����2���)��(��r'1=�������(�&�#���bU&�8i*=th�-��<o�N��!B=O]�Ȍ;`.�<c.��������<\&/=��Ժr�=�qU=�mR�� �>?X�������=6 g�']�/�:='�=�#=P%Z��,G=Y�1�V0=��<�n<y^=��x=�>s<.h��Q�]=g�<[��<0aL���>=������<�܄��؆=��N=0Z�h{-�D���K�]����Ԣ�;��]���=�j�;��<�:��6��<,��<ҫ3=!	=�=��G��|���͝<}B��-���0(�53ڼ)�,�lo�<2=9<���<M}�xg^���ü��<n�<��=�!b�<Ji<�6m=�u:��+R=�X�<q,/=PC�=�!=�~^�5����C=~ ;� \=�1R�] �q/������N�Hr=��<�(ʼl虽�=>�=5a���Af�������=��D<S�=%��<dϡ��ّ<r�w��m�Ib�<z�B;'&�;/м����ɘ_�	}<��~����;	�<�oݼ_��<;q���<_�47f��em=i =࣠�}�:3Kr=����3���S5=���<��z= =0=n�`<����H=�ߗ<��<�j�<	�2�|�d=-G=u��<�`b<	������9�U1�X&��[W��|�P�n��b=䊦�a�M�f�<���=W��o�G�x]�<��W��-�2V��X��3F���X<N������f��s�:=^F����¼"O
��%l=E���"<�QO�:-���O�٩i����;9r<o=�58<<�=]
l;��Y��G�y��=CP�M�y��
=�+��3�5˾<�<4��<�<f���X�LJ����B<����IA�sf =�)�<j���zh	=��/=g;��ߋ�<���߰��!��gI`= �9O�缤��<o��;[�����<�����"=O�3�:�2���1�FUJ<���.= �E=�$�K�<�L��q&���<���1~;�蜼IZH�O&3<0��`�j��D0�y6A=�==}=��.=k�<S��<��ļS��;�dl�����:�<[�5=�'��:D�;�_Y���P����A���=�B]����3�ʼ��*=Y�T�vRT�uk̻-ļ��d=?w=��	���?����<$��;K=�=�v�=��,��ۼV��<�����1�(��;���bH����ݼ&=�c=k@�<�<�c�<d g=�`=��+��;�S=�0�<����<v�H<(�<�~���X�<�
=�>�e<B=W[C����<���<?p�<��W�]8N=��<��1�P_�<f=���F#<&����Z�;w<�B=�6=�e�S�2��{'�c�,�L���%�����:Q3H<i�<��f�II�=�
�;���;����6��<F���^R<��ռ8�2��d���<7�ۼhS����ѼE(��Ŧ<�<+�ɻ���-�c=�?0=�+D�[m�<����K�N-���Q���&��k=�>=�z�{�N<�(k=�9f����<��<�U=�������-={�=�L���e���<Tz�<�֡<=��ļ�k��k��;��g�3�m��<�,�'���ml��E�<����F���$=�N<3^=o�W�2�o<��;�K�<�lK�jL���!H=���թ��Y$<}�<�����~��Eќ: �e�R��(�޼��q�u�,=E�<#��;���<o��L���R�a��P�5��U�w*��W;3<l�J�q;�<�M�<�"��E)�����@σ�|��GAN=F�98|���']��)��i�S�=C�=��<=(ռd"߻_F@��B=��Z�i��:���e�<E�����<�G;=c(j���:=��z��!#�����b�K�=Sv"=��<7���;�C=���uB��"��Hw��:��`(����P��=C�o:�M������ �<�J���<���<�6B<�;�=e���A�<�{���B��`�����=}�=����;9�u���B�)��;�l� -���ӓ;�����^�;�:���U�t�8���G��i��w�0=�_B��=�+�2=^1�<�&ټ���<�j�<�n�<��:��$����m� =���:��~9!���,�w��<�2<*�v��Nq<O@D���T=mIV=cb
��������\������<9�<��,��v=�b*�$��;�@+<Y6=��e=�B`<SО<ҽ=��=��G<϶Q�0=*E��AA=�� =0�;;EF<�&<��o<�渄,���V���S�	D����S��?O=1�i��@��Z������5�<��;��,��R߼PT��dr�<Jn=Or�َ9�=���<�9�:���@��<�6=�/"�c��;x~0�JK=Q�=�̸��G;='{;=�2�<\�=���k+6��;�𾼇�<�&�tb�I��Z�<����L]�<P��(��g�<m��<��;Ҽ?5.=h�<%�(��U��R�W��8����<�a=r�<��;�K���{=J�</��<���J��;��b=}�<����v�(��<]<r@3=)5��	>���>=��<6<d�iN =�Kp��+�x���Uu��=��=_�<2ټ� =�=�<~�ż!��<��ѼA<��"�~<�M^=~8?��}=|���/�M�#�[=�L��+��T�<�bW�9	�<nv2=7�H� =�	M��\=yL_;��J��?"=�r��l=!Z�<i;�9=u� ��EȻ_p7����;Xѓ��M=ZZ���X=�ͼB�)�ȁ�<PR^�U���{�/=J=�7ȼ���^{��W���<� ^�[<�����<[:������XT�<C�ؼ.p��-oO=�<�2��dQؼ���;�^�<�Go��~��Y���໻��m=l�8�ݮ�^�<xv�=JRG��<����!��<�>�<��<"?=5!&=��=�����:!����<�;�;GP����=�7�<8lE�7͔<���;S�%=�h<<�o9���P=ר:=����݁<�N�=��[=Vx�������n=�:�<��'����7�^=#�m<̾L��_=�U�M�^M>=�G����ZY�<���J.�,| ��J�<-`=���<]��_*����;꣘��z=g��<\[<�ߚ<�<�=v=�G�܊)=�$�:�����;��\�;6'(<.���b�������(n����{�2==d�<](���U�z��֔<L={|��L�g����=�����2=X╼�q=�p�4:/�f����"=���<N��<P���dO<�6Z��e2��B=��;�]=���<�<Y���!HK<��y<i�輠���2�^�^A"=�z}���;�+=�=�Y>=p8=A�U��򧼺=E������-=9μ54�<��=)kؼX��G���8ּ�[@=Xg=)4�ȿ!��1=s}g<]ݶ��TF:&"�<�{�<�6	�f�μ���<�����Q����漎*,=․:7��;K�=�u =Q��5�J���\�>`@<���<M:<�=�<@-,���Լ6.��`����h�^�� �<>�!;z<����<�^<4�a�Dz�)�t��f�0�T���]o������\O]�!�(=1�t�t<��;2�><� ��R�<%|���)0�V����+&=40/=��(��9�?p�<�O2=
E����=�e=Z��<F������<鼰�Gf<��鼔��.�=���<�V��n��-=ms"=��q�����9D�6��<rN�<�� <��ϻ*��z`��w��Mm3=�6=l�<�7�9F6�;��L��S�/&3��.W=�t�^L�<1`Q���N=0��=�C!��޼�fA����P�=:�{�E%d=�!��C��؛=��g�k<B��d��ř��]=U+=��o� =�sV�+O�s��Ӱ6=�ƶ����<�O�<�!��0i�%�.=�@=,�ڼ�o�:�*���'�<�1�;���<��x��|��EB�&}ļ�wL:���<��ƻ��<=���b��<�7�<��;Q	�
[�<x�����<3�b���>=�=B��eK��jJ����<n�=	����X�2���=�F̼��^�V�<�d:31�=%+�~#=X1���(���L�;���<�}<�;��F=�h;<L�xҘ�2�y=�<��}(�;SH���%�O�P��'��L:�ڰ�e��<
��<عMvC��aȼ�=���wһ�,=�=�<֣�;_����~�z�=@G��S<�>���Ei�+ۊ�uZe=�Rh�5;?�]
n��f=�VQ���V���<0�姚:.U!=]�<�r�<s��<�&�؃��hb�]?1=�Q0:Q����C=T�/=���;�=e�@=�>μ������@�����,<���<����nF�<W���8��<�a��+=�`=r��/� =(/��N�X<�ݍ<`e!=\=h�<M�X�ڨA��[�<I��<��H�ڻ��i
=��=� ��4=���9�=o��J� = �J�=�B;�1�<��'����<q�Z���-�M��< �1=5s;=��'�U����<�9@�'��<.��c��<{�u�Q�<��(��7�T <�=��C="�ƻ��jZ=|��<�G���_��=D<�G��"=�3�Fe.<cv���j��GJ�M2b=x�6���=�(<F%�<��A=�i���=٢�x�!=�a=�Y=�e=�]y�����]=��6<+w;77����Y�
��<�^3�?�c1 ������j��*�ּR�V=��w1=��,=^ ڼ�l��%��;mЖ�@�M=��6;L�J�xo��[�Z�p<oK	��"=9�<J�<>�1�DY>���=!Yּ�猽�ٔ:k0@=�x=�Z�����<t༃�O�3 ��J=�N�:י]<E��;��C�E�!<ݡ�<d��Z��a?ۼ:�<���:MB���y=@9�eмb6j=yۋ=��>=�K�!=,<�x�;X�庭yP=DK*<�c�<��#=T�"=y��<��&<B��S���~�<ͽ�<PQ=X�;��ݻ���<��1=�߿��m@=���;����"<�D�<}�)������K����7=��4��I �\zu����=�C�<���;����&��:`��|X�<��;�$��m�<�)=����<޵��a=���<H�<��<Xp����(n=m��;N?�<t�:��f�NtQ=�3(=��J��M=�oV=a��K�<�-ݻ̈�Bk2���/:w�%�� :=O�:cd����<��<P5$���L���z;6�D�S���$��Ę<[x��H+���������(���#�<ҵ�;U�g��ϊ�{�u�g�t���Y=-���c=��˼IX=b���/K�M]Ǽ�͆<� �<K�����<�䊼�;=���;�� ���=gw=������9��<{Wg�b哼��@���;=?�:�l"=��W7=��H�vbԼ5j|<����O�!��ĭ<kI;`�Z��F	=@Aؼ��6���� @=�@9�;�<�� ��n%���i<:ü����;([=��V��m�xt"��B����4<y���@=�(��E#=b����F��k���S=*.�I��<�S�T�;�Jd�:j��2��<6_~<B$�d���&D���<��}r=�!$=�a,���wNg��r;�U=�����3=��.��n-=z�1=���:3<� ���9�vy�w%!;�͜�~�=OT�<c�Y<2�<�
(��F��`h=�ц<f�,O�$�k���"	�	��1A�<3 򻤸Q�ܯ�;��:�۱;w��:��ü�k�<�?�<`t̻^�.<��<���<fV �N:=�ǂ�u��L��=�T>;��$=GL��;q�<|֜;If;�zɼ�:=��<��<�=�:=��;�;=`=Hfe<��м-�<�	�kۣ;�$�<�_�j� ��)��@�<[�<[��5D��E=�IF�2��<���=�s"�x�<�����*=j�I<\t@�R��?�<��̼��o=��R�~gڼB�"�.8�=N=���Q<\�9M�=�8˼aG.<&q@� ��d��.����:�=�B=N-8�W]�<UK=OC�n�߼vy����;�iA� `=���nB�?Z�u�	=����:�t�$<��G=B��~ڻ3z�<�z>=��<�3;�V[=�	=0�I=�,�NfQ=C�7��Hb=����}+�O�����Ǆ��^�8���l<׬<�[`=�R=����L�%<�F=�Rg=�B<^��<�L�<Le=
�<9%R=�,?=�|���V=�a�;#�L=]�"U���;���<̻�<O-����<�r�<�����#=�9=��2=�&���\���.=p�7��X�fR�<Gn�<��<���=5��;¢��%�< F��#q;�ۭ1=0bN=/�<G�m���(�H��R�<T[�<��j�wؑ<Q|Ѽ�lݼʄ=�-��N2=wO��S��̻e��W�
;Y�H=���;�� ��.g���<ϓ�</�K��`f<_��_~~����;���<��M�=���<��x<Y)';&�=�@=��=Y_μ�|B�&c`=�t���x)=�h&=`�x=yj��/<>G;Z}�=���,y�X�
�����@�/�d�Y�ݼa�=:�<�7=�z]<��^[*= ��p��<�><3[�<ߊ5���4=C�ڡ;(�k�mn8�7�<~lN<�j<�W<G3F���=	<�Z���+�����l�2�;=��;������	=*�<t5=j>=�<�#=.�<�y�<Ѧ����4�F�b
=���:6B����B�e�< <���-=~���;�3k=)37��]��;༏v���4<?��<��=U��<�W�z��1�<��<F7�^T���=�
�-� =�.<|��;p���R�<C�ۢ=#$�5˭<�yk��,=�d=�^H�F�>�[H��
N=ϟ��|�<)-\�=�^;S+���z=)�{�PN�����>�uUL≠��Bj��Z�M��
xL=ȃ��S�$< ��<�o)=�<�<����{	�g�=+%�<WF'=z�B=곧�g,���:��=�#�=��_=*L��Mؼ���;�QT=fA�x'�mo��0p=x�;�u�漊������Q=��==4��&���Q4�Se=#�L= m6;�b�<���$0=B>��?�g<�E�����<̬B��O�<@/̼4�$�
� <�

���n�ӣ�;��d<Hcj�����M"=%�k� =V��<z,��뼼�S	=�#0�Si���<�r@=�0Ǽw�N)�q��I�<���BC�j�L<nJo=y_@=��/=;x'<�3R=M�<>`!�����#���(;�qR<-�c]�<.��"��Q��y�мn0U�9=�w�;{��<���<}�B���>=�5�XBO<��=�r��=%9���A=��B<0T�<~ ռH"�;��*��T��5V=���<�3=.��<�9�}Lx=[bG=�f=�����"���3���j�<��<�|Ļ���*�ź(�ۻ�=�o�:>�`=%�V�ρ<�8�<�S=�ۊ<��J�<Zٺ�]�<_���d���`=�n����P=���`�����<��3<\�٭�J��<�<�R=85/���=�_d�ۻ�<��&=�Q�,�};��<֟��Q��{� ;V7����M
���<�r2�	9ͼyUm=�o< �)�3=.�{=�#y;&x�<�(&�/�A�$s!�!��;n��;D�d=��ͼ�p�!�=r=BCz���8=G�< y��|�=p��ּk F�(�;<a��%e���F<̰�<p
��~�;+W]=�,=5 #�����;�,׼��=i��<X�o��B=�JQ�����=�O=4xw�7�w��XH�s� �B� ��dl���H���U=�R��7<\�ռ��b=ZF	=]Ay=�k<�=�XR�ʇ�<7�W��M�;�~
��c$=A��W�<,ـ��eȼuͣ<T�<ۃ=&C�nID=#ӽ���8=�>��dQG=Qr7��/�~�<�?�9��U��� �}�b=.\�<D����oU���%������$�<k<_N�9��>�Ẋ���<��:�� ��C����~�p��w����a@�;0�`=#!�<G�==�2=TU�:�ڋ����[Q�:'�Q=;�e=X,=�"R<4��<�M=�����W=1N3=���<�f=��E=���<:"
��b�;�A�<^UH�e�<�;r��|�<��+��=����W='�n�����r-3=���M4J�e�-=��k<=�(�;;�<D\=���;K�p�߰ �&�X�_�Q=�c$���N��c'$;��<#�;)�(=Pj�:bW�;߮V�=�;hZ�O��C��n=/2�@q�<<�)<w�(��t*���-�r=J����;�U�Ț#==���L��<Ӗ�X�"�OO�<?��p��<tMB�͐�4�"=��S=�/���̼m =]P-="{���»	�b<�*�<͹$<C<Ue�i�=P�?��Kq=�C&��e<'����=�y>���W<T�<�cZ��}N=�C6<�{��nw�Y���s�E�QB=�#W����<��d���=$�h=g|<-�=8B��J�E=E=Kͯ<RQ�<� Q����:^�ټ��<�o,X�&�=����Nt<B�C��H�:� =\B���ջ�<�Vu�s�?�U1@�0ꝼ�v���\$;�Q=��<I�)��RX��lR�1� ���2��ׯ�sQ�<�6:�f�<��=��.���<=���<���.��<�s`�~ά�P�D=�C�<6ǰ<-���H���;�N=����W�ػ���;�F3=��=�j��<�:Yּ��5��*=" ���}�*y=�<-�.=k���ń<rK<n����$=P��_�=��#��f)�͑�MN���}=s)<g�:��b3=f!=�V�<������;̑;~��<C�n<���<��=uR�J�O�,�R���4�q�E4<<�N��������3w���T=)Fi��M=�Vż�ʁ�׀'��Ã<R����=�l<�<I�1=�T=��?=���=�>�_LY�cf=њ�:�'��Y(�;���wj2=~�Q��Ù<��=��=V :��&���[�yz�	�r=�oo�d﫻�o����S&=M�ɼ���Z�<_��<��I�<�g���<��a����m<M=c=��D���;P�L=�zq��p�&��',J�,)=yr���X ��8+��=���;+ ���,�<�e�<��<�C����<�r
=�/�7hx�w����t=12���c�=���]Ri=�u<��="���q =�z)="i���P�x�8��F���茼�`<=-R��x�&=�0<������嗼�����7���Q�J�-��w[�I��� G=��'�������м�	��N�081=jT����b�5���f�����1=�2�%�yX����.���d��9��<0M=�.%�t^�e�<�9��e=8�J���0����<B=\�?=�0���:�;x���m�9�3������u�������<��R�t������r�<A�h=PM_;hLU�Tn9=�=�$N�k��<����!�j����<������{Yd=�K<�Ó���d���<�K<�iZ��K����]=����t�f��u^���ۼQܽ;H�=/�<�M=k�"�T=�e<��f�q����<�Q=g�<��ļ$"�<��B=(k�<	�k����<:~=�6<��c���H�xE�� c���N<��V=7�=>a�6��N��<��1�QcV�Z��.@/������:8},�b,v�E?����;
�<e��<��K=����� �L=�(�Ҧ׼�S<�A�<\�=�;���`=v_=HJ�wGP�%��<�a���$�u+A=��.=��==����s�<��L=�S��;J���&�P��\���I�]|4��8:��<[�
=�=�yf���<uT�<���-=�e��eP�����:#���V=I9=եӼ0�T<�4�<�zL=��;��̼Do7���켝�	<�)�JG#=Ȩ�������=�ˤ���ü�d=E�=�!=Q�<�� ��q�<|�R���B;��P��8F=�B�F"�;@(=R=�׻*uۼB�<kX����&�ܻ;�]�����M��<�b�:N�<�ڃ=p�ʼ�b
<|]=�Y,=�x�\�T�^��<l���9T�;x�!���<�b9еj����������>�Dˋ<�3o='-`��O�Y��<*�?=%	���:���$��c<�\�$�H�"iɻn�x�^;*=�&=Pf�}-b=e?
=��5�q��,ń;]=r}9�R)-��=�-=�7=�kh= �<��<�����B=w=|�����μ�D;�3;��K���m<�$�ʜ�;IoF<�,�Y輎]��,�#*=5
�<���<d(ػ��W�k_	���'=��v=4�;���;�p==���;@奼�і���K<4	]��>���4/=��9��,=�0����(=���<�=���<|H�;3���(h*=uJ̻O�Z���=/�0=؁*=#�<��8=z�w��Lؼw�7�7>�z�+�9�D;��M���5={�$=�*i<Y�=[�:��=p=��[=6�=�i'=$� f|�7oD��+=(-=��;Ts�s�`���
=��6�!�e��9�=�e<����k/=0���V�<�X5;�Y���.= �R<}׼��K=����Pt��F:=�w=	�C;�K<��<=��0=�(N����;h0�r�8���j4���@<@�G=�<�X��}��;��=�(���b=w��<�JY=��s�'�)_��|9Ӹ�<e�^=ILP={�=~<�<�w���l����:�$����fK�<�����T <�[�<<�c=�S"=}���2$���<��1`�<���=��<���@!����<g��<	9=]OF�v$O�'Yu=��(g�:��<#�<:S��l�%��=y�)����;^G�<K�n��G�.�92��<�<t/E�jLo�F�-�5�<���Bp=�N�A��<6:�<�f ��K<�����/=��<v
;��l<�=}��ۼ/���X��2�<��o=��3-�<��%���L�<�`���!=
�;��<��]<,�<���<�m����d�=�-�<����������<w:{��
⼌��N�C=��=��F��Ht�$' =j�@=N��x�4�R}B��f���ؼ�i_�禎�t?=��n<�^E<��"=��k�<2Y�����<�+-<$�Q�Tt <a<="N�R�=Ŝ����<c"==o5��T=���<*��"=1F��a<� 8��M9�����+�����</���ܴ�<��<�e�-�=ԅ��0� =F+=?=v`漻ټ�~�;�'_�Q=���mXJ=�����:3�=�<�&|���=2Z>��3D�d+�|�N��=�������;\T5�=,�i�^���������~��'���K1=�L�<mټ�����3=�~&���=ܻ�
&=��:�¨W�`��s"�;>��;�����=\�S&����e=U|,��QջK��<(M��l�r<4);�[a���ݺ�¹���<l=�G���y�wi�<	�=��<�$>=�(K��׾<I�< ���*����<�PO�U6�R��������h�9���yN�Ԫ���:=����(��*�?����@t=�N��)���I�<��8���?<CRռM�<�@=��{��x�Y򦼷qM�1R���T�� `=��;��v�v��������<�8 =>M�D���:<���sM=ZU=z�w<��H��@伋{�<�;��F=|�D=�t�-Q;=�"1=��M=�<�������<�]�qC��>�������<?��zzO�!�=Vn�<S���x`<	�==U��<Ye�u�==���(����j�$�ȼy��<��X=&D=:�:D.�Z�t=f;*�v��w<�5?�����8Y<�r'�[�*=;���#���n�ǻ��<
W!�3�2=�.���	�� L=a�<7!"=��G=GVC��n�&Fr���:�:���'=�t(=4O?��%C�kO��{=�����V���=\A���v<�8�# :�,A=���؈=�0�<O:�o��<M)=�a^���y;��=X(�;�ez�TtP=�!_<Gp�<���M��7:��\�<�m=��Y�rᠼ�,4<6��;>#�<v�b�LQ1���;��5=?�=�%~����<b���������'�>��;{�:=*9F=�:�<>��'=8��<ڍe���<cْ��żq��h��:)@;B_3=���<$&=��=M<KH�<ky�Qx7<�8,<ZJ�q3%���<<�5����&$<�:Ѽ��O��:%=�-�;�6=-�G<V�1=�n^:wT��3=���H4�lvļ;3�<��=5>���ab��W��<y���� ��Añ<f�n=�	�s�<W{^��j�<6�"=-VA���`�c{=-I2��'̼c��J�&=w��x�g<z�J��j=r�==�L[<$+�<�_ļc?��	E���+���<O.=�=r'=���f��<;���ڼ�7X=݄=*�����F�F���S<x~�����9�<ћ�:�?�<��л�7=έ=�1�C�G�����ƻ�0ǼPW���G�3�==�%m<s�=Y�=9k�����<#mR=��>=@����<��C��k_<L_=�DƼ�&*=$�V�����	=U#=�Tq����95rx=��#��)=��R�Ʒ���{=�A�<�BD��N�<��<ί/�p��:��+=�üYt����_<wÀ�J�>��(`<��ݼ����=�Ji=�n5<ー���<4�)����YR4�e�=a�>=���]�;�e~;-R�<!���C;�\�"����(`<��<v�U:���<Az5����M�@��8��
�S�<�%׼O�P= ��i=��>�1� �;=�Ur�Z5�t����U<F�L=��<N�<�Jʼz_��x��h��7D�|���{��<4�H�	���t����<����{���R�<���?/;F}��	����"q;_cb=eWb��#��߰����=+�T���ۼ� �;:&μ���yƻA7=䒇=������<ǔֻ|�(<�\�<v�=D��<�=.o�<��ڼ��<߻�:d�w흺��?=ѽ<�i�S�L;	�S=n��<(�=f\�lL<CM=��<;ǠI<�hp�ʘN�2�VǼ=�$�j=l��<��7�T˼��R=�O��]�/����,2�+�D<tu��lJ=�#=�7�;x��Os�<� ��)EǼi�����a��3o=��@=#�<��C=�'=,I�;$+!�����_M���=�
���a�Ky"��E=�`T=��~=�ì<��bc$;�
=�m̻`����=֜����<ҁ���L6=y�=P�{=�O��p1�<��=�On�sX���=�B�?�<�j�μ��ڼ�O`�%A��x�<?�$�`G�;m��<뭎<ˠg<^�m<!�0=��W<i/��	J�Lwv<�<<6J���P=5Ck���{��S=CU��$���k�:9ge=� 4�ږ�<��=�=���<�=Z��<�*J� J�.�={~<J��ZY=����`F�1A��*.=��=+ӻ��=Oy���:@`��|��x=\����H��������yQ�Y��<�^A�\�d�v3����<k[�_D=��;�ǻ��Y<D%(=�!=���<�=t�����x�P�L�=��ۼZZc�n�<�'�����q�߼�.���j�"�;�α<�?�1* <�S�k6=w����8�<�i��N$=q���I��}�<辡;,��i�M�?��:%�<٠�?�)���N;p챻���3=ղ�;�]ܼCP�<)a�<~�����j;nu��3i�� L�U�;�fǼV���@�C;��<g"��(���=dݞ<6�9�H_=�D���⚼��=G��<kN<�k&<�MI=�B����/����<����o*ټ13�8���<�Sp=w	H�~s*��p<����l3�菭�3j�,2���I����|;܈�? �L�I�L=;���~�b��
=H�==�I=�&c=�<}jy:��;=/�<�7�kK��=k"�<uR5�L=2�f��A=�?;K;�P3��3=�M��w�]=f�ۼ�6��{:=7���̻H��W$z� �;p�=O�����;b�>;��#=�9=�aN��`�������<Je�z��<�,=iN2=LV�<��=�A[=v��4�h��,ɼ�]+=J� ���G=xƼ�F�<䱼����UDi=kE�;������c���<;�m�<�^�<��=Nݗ�U=�z=nR=)��<z�Z=n��ڼB�M��u8��Z켕N =�	=�D�<�oi���9=�mh���<��J<hgJ=�W=��.��_ȼ'�W*x�n94=����uP=p;@�(=��>=�Xm��b=��'�Lֻ�J�K��n�<n@μP�4�q^�<U��<�����=4��o��;�<�P�����!��<~=��,��z=�:�:;4Ӽ�)=���<�3	=q� ��)��ԫ$=��<Ӫ�=tn���
��(<�P�=�=|��E�8���<�C=���<=�)<�F�g�>�7�3=%
��U�<I�e=���;]VM�g'5;�y�<|붼^�h<�EǼ���=Q���=�;�-w��R�<��ؼ�j<�H=
K���"�08��&���(�<��漪4�ގ�=���U�X�hn����;�@e����	�^�B�G��	=����.�<��Y<Pn�<�d.:��<��[�;R�=�ټY�9��V�[��<ըA���c<ێS��A�;ڦ�;*�;=P��<��V=�6m��K�;ݒ[=�(Ƽ�L��="��飼z.<9':=�^I<~w̺��<b7<�G���='М����<B;���%��;��w�eZS�_�8=�d}�>�Q=D��A�k=�J�<;�1=��+=�3=�G�;���<M�>��B�;Gd���p�J��; `?�e9:��<��_<{)p=be߻�e=&c�<�}L=���<݁����k����<h�<ۣW�i�,������=��!<�Y=4A�%��<LO=qP;U�N=`	�<�%��		=��<u4I����Xz<�p���Z����<������;���bt�۴e=�4a==fp�<T�3=�E��F0==��.�f��� �f(��aQ<3�'=k�<�f��VS���<̨=GVq�!N<�̼rs=��<��;z�����?=^[�K�%����	�<R�~=�yE�g��A{�̘���w�[�����g�U��B�<�˽< �Z�xrO= ~	�sj���6���żD�{=�����<E�=�]h=�$�sD�<C%=pػc�׼r��;(��<߷.��z�����Kl�J����_���0��@�<��[=���:�K��f=������i3G=��g=��c=F�=~����J=R�����k�>�d�7{<�2�=���ǹF=��1����%��5�?�]�����ϼ�rP�ϟ㼕�=|�輻�=�=�?Z��4+4��Q��S�L<�q='�=�f!=�V�<�����x:�U,�5v�<��B<l�:=��:-"=@e4�/�T�$�2<�-��ӽ�,p�<#��؇=��;�u�.hk�Xl<�9�<lʅ�R���4"�+a��^�=����^Ӏ�xN���ɻ�7��"�LS=Ǘ>���;��˼KW�R�<���!<~���<��+��ټܟ�/T��-=	]�<�۷�<��-=�K׼�Fb=7�<��M=fU�<R�𻖛$='<�њ�\k4��rA��Q����D<!-�� ����<^����p���]$<Ȉ<��g��-���U�9��$[=Ď���8�<���*�I/�<�=�)�<�<������:=H�C<3C=TA<?�_�^�=�*�<|cL���\=m�<��<)��<��4��+�Sw=,�<>��<�z/=K�K=H7�&��<��k��=�Y���(=�T=A���y�=��<�D��x6=M�Z�ڏ/=a�K�6N�;gQ��i#����;,��W?��yK�d:;t�X=PJ��R^=�u�<Y�x���,=�����k=���<�U<=�I=��'�V�=`����;<=-��<x<�:|=B���~�N�����|�<@&�<��k��!9<�=Q_��>	�����<�;(=,;���8�<h���<��n�֦O=�=PL��=����:��;�?<��V={`�<�"�<x�J��]C�o��e��<-��<H�u���n=�3��w=���|��<܏�<fP�G����&���<+�0=�@�<|p=�@�s�����%+��l��'߀���.�#ϒ�Ey<,>)< �N�aY=yZ#�@��o���:��^~�:.=�&�x�"�=ɄڼE�9�NM������D=��;�hF�B��Bɳ�wT=� <��[���<�O=J��<�n=K�0=���}�n<�Ձ��yp<öf<�2b��R�:===30߼CYB�����ڼ,��<1����OU�Zlq�p}!=�D�<�k���K���t���)���Z=f�<'"=x]u��Me��˼�v��O�<OVu�3c*=�9��c
<��;���;��N=c�k��f=��<����s���Y��M���7ü]�[�wr�����;�~�<�O&=܊O=�͋<�7=�5����X=C}�\�P���C<�AT:O����,=n)��E��=  S��;o���Y=�D��#oѼr�=�~b:�4��|�m=��9=O�p��j��������&��������<zv��	�w<�0=$�*�!p=�:Z�Q>)�d�<�%�!��<��\<�;�<�N=���<��8;p9m��m/���J=}��_�i���i��#��;=üO	=R& �:g����<C���F/���[;� �<�k�Cu=�� �!�=S҇=e%q��<=�Bi��]6=w$��H��x�<˳�?EN=�ґ;P��<`��@=K <^�a<��v=��@=#�<*�n�3<��ϼ����T�,z�<;�7<u8=zY=�X�<�I=�^�;5=*��;�X���W�<� B�j�¼Azi��z=�W�<�c<��<�-�<
�.=�<��7��`=3���S�M=��뼍�5�$�?���<����]H=��<(�+�.@+=� <�j�6Q@=ŕw�9;b�1z �p»<D,=� =	*��NY=��+��E�fC�<����J�xe=���lӰ�y�T��SG���`=T�s�P�;���;��B;�E=�D=2� ��h�<�=u�p��0��'K�m���#<�F=���<�,�@�-��,H�V�ؼW�<��/=p���0=F�L;Q?���]�<��n=�xr�V\6=�	R�#<3��z�0s���Ah=���;��M=��~�x#���\=���<��=<�6����E=b�S�`9�<�� <&ܼ�����%�<�=�<n�<��*�[o^=t}=�C����=��oI���e=vڐ��4���:�|��<��G��7=�k
<f���yJ��B�����{���a=��K<�e1�\l�o��䑼�<=�܅n<�aU�a���c����;y����E���E<�|J=�'�\w�<�=]�I=j0���<�m���6�mY�S�=I�5<�4I���!�8ot
=��;=K�O�sRI��`�<Z�<��4;� ����%�w=6Wj��
�<Y#(=ȏB<�%�<�1=�kS=��:�ě�=B�m=��_8S=��<%f�K� |���<��=��Ѽ�q6;�=�(�=ɽO��!����<L��ڙ�<t#c;�r�<��3�yGN=�m�<��l�	�V=`�$��w*���D���幻�Z���"=���<}@ =���.8=���;ZS|��0�BO>=M��<�!.�y�o<�B�DKD�0�<ڴ̼.��)=&�������7=���ݪ�k��j"=��<&m=HںZI=���<��_;������X�N�?����<"�_=^$e�&(Z=\K��&���^#J=Z= 8������A��=-��<~$���=D==�$�<�[o<W�S�����3��;��;<�x�<�2���*4=�O<�0�<(�=�i��;�F�<̪H�ۆ���� =<ᶼ*�ϻ2Ӯ��:a=�Q����<Y�=Bg@<*X=u�ͻ��'���/=� �;/�%=���83�`=�X�/��wd��'<��V����LbB�� =�������:�A�+�<������=L`��mG�T��<`;<s�t=�
=� =�"�;�1����<��<2��;x1�<R�>;�%=L��\+=���D�<l��<�a�G=Rb�<��;��U<��<�WG<|��:{���G=-iҼͮQ��=�I��ON=�3�<r<����6=���S[�%Z8=�=q`żC�<'w��$B��4=�I(=B�=Y�<����<�����=8�yr=��"�$�dW������ ����s���	<m��;�N=���<6zἔ�</a4��sѼ�"�:�F���a=♑�s*�<���<9;цz=��8c��?��z�S�z����I=��[��!:<�s���5��<�=I��<�G��a�K=��X�'�=�Vɼ�d@��J]=Dup=X�ż�� =F_< ��[�N��Ŏ��(=	k=��<�J�W�,=g�=W��<��F��O=z�=��N`G=���:�6C=�[���e��;��.=0�K=��=u�<<�a=�>����=��V�-�����<�i�<+0�<�_;��γ<3���h�;$�=���<\�r=�/�qh#=�pT<�-=�J�=e�<
2����V=cO���<ôU�-l��Ds�7�ޚ<P)��Ӑ��竻i�.��=�< i?=�7N��ɼ�ͼN�)=[��<��<gyH=�dH�ָI=��d����eB=�R��T=���;�Þ;QȔ;�F|;�t��q=��<6�^��T;]Yd=6��<�x�<K!(�K	=`���#==7�'<��8<��<z�^=�LR=���;�R�<�:�mQr=h��qX$=?j*���f�b�b��;�bM="�}��t�����<V�<畹<	;�<�#��m	=Ө#���,<�VZ;��=6O=��m�q��<
%���c�G��<.m�T=�N-���<���<�=.tn=AҌ���<�$r��g{�Kp��~$=��<�v<�vK��`غ�[5��C��h�<�!<�H��78e�sּ��<"�	=�)'���F� ���[����?=c�!���=k��<�8<��3=%�=������\=�=G.�R�\�Jш<J(e=Ĕ�8��˺��`�����?=t��|�j;	�]==�<��'��;s<s���=+RV��=w�Q�HPU=��u=,�<
��/���g�ؼ� m�#�~=�=aSt�iSs<�)<=�l ��x�=6�=�I(��\���
Q�<-��;ino��m�<��rk�<�C�4<���֎�G7�m�g=A0V=�]=[�:d�N���%=��><��g;�V&���<�6�z5�Z���*�5=9qk���<
���o���uv0=�*J�l�=��7:HYW�9�[�4Է��;F=�k��r�@���	���H�f�2���=vw,��Pڼ�݉�5�e=�
��.xf�_L�=6";���<f������
#�<�l�<+++=TY໩�;�8���1�<�(��f\�8\�� ~���k�<��;P>Z��q�F�=���Q���*=oT=�\�UC��l$��1<=�p==.���J�5=@'��ߋȻ��<
T��lnR�^�P=�Ty��۱<�6���V=�v���z=�(���ռ^�I;F�.�&�<�ȼ~�ɼq��o���۸,=@�	��Y��^��<Rh�?�=q9�<^�+=$�E�4��v�r����<޽�<�=��n��<���<�A�9��U;K�<"]��� =�N�<R�<i�l��8߼c =Pta=e�<jn��O/=����W�=,D��wO�G����,=�@=�==7N
��`(<T�d�d�J<�R�9�)=H��;� >���=o�N��;]4�<�-��e��A���lӼ��<D.j�Pv9=@�<ſ��$���;��{�+~ټP <o{z<1�=��2�<�.;Ku�}�C�KU-=ٴ9=Cc=Btؼ$q<|O=���=�6�<�\��B�����^�#�<��;z&K=g�=@|�<��Q��c�.*�rCs<��/��q9=Ύ;�3���ⱼT=Q�XRV�߹=��3=�h2;;�Q���Z=�T<�R#<
�.� WS�NdW���\���.�%��;@N��b�>��Ov�+9�?��<����S$�~�e���7�Y�ϼ>Pw;��Z=(,9=�q�����Y=�XW�<��<1�e�*��V�W�Y�$;���M�<��h�6�E�����m'=:L=��<�N#����<l+�>�Y<9�u��t����<8n^<�>=Xc���%�<��;��f<����i=K*=�4����]K��;`x�]�Ҽ�D*<�#v<���H�ټǠ=4�,�d��
l�ץ(=��n�&F��q�<�
�5=�U�<g��<�7>;��u=		��ϺU=��Z;�VS��#=\AC<(�T�f<�<p�,=�𼫚ͼRQ<l�<��N;H�-=;�1=�!3=���d�f.ȼ�!��H�H����<��R�e@��,�В<��l�[�]���\<bW�mTg=��(�3R=���<�L��N�ؼ[f�FS=�r<q�T��9���<��l����G-��������$Sͼ��c�"%^=���� u=:ZǼT.�<��<�����CV<�F��c�Z�!8}�t[�<�hE=މ=C�t=���;�	<�x�<���aN�Ъ��~�<���;e����?=�N��X�<]��X�o�zAP�T=6�ar�<�uh��2;99���C=5�Ƽ���<=$�;�����=7*��@,=����r���G{���޻��]=l�]����U�;��F��d���[	=Q��<ǈ7=��������(=�<%���3=�g<, ���Q=�w�<��D��뼊}��E+=3JK<�݈�Qӯ����_m)��1=񷼽����nH�W�<x=���tN�<�F =Z�4�s��;�%L�Z=�XG=��
=�T���!��=�ꌽ(�N=�A�;�z=^�vJ=&c��R�s�l��<aD��]��<�rD=���<�G]�Zw!��9�<	�S�Ӣ�<�;�fS<�ܱ��B�<ϖ+���=�0=!����_<�j=��<=��ӻ�-\�;�<GM�<��=6���)���g3=�g��p�/P�<�i�<� F<`T�;w/<�G(=��ֻ�*V�#-O�j�V=נx�۟_=�z=���<g�ƻ��e=�׼�b+=���g��3��p�<���;�ܼ�'���G��=��u���="7�<ƙ{����<	�$ �����<i/=�ɼ�=� ��!-?����<$�
=��A=��@�h�<6���g�:���,�a=�*<#G���)=��G=�ĥ��qg=T�2=Z*�j_=��7=ȥX�˫�<�ļ�R=��=�J�� �������4k/�'�<A���Z�;�?�׼�<E�8���I��;y�A=ŝb��1����=zT@��Dּ�4���$�0[�2kN��[�=��<���<ha<^��p7M���m<�c��X����=(��<0����<�W<x���d� g����<Y�����`:=N=@bW=/�C�(�f<w.��	~�{���^�T���<�^�=��E�X��<1zZ=-�༹j�V�`g;�P[=�ȼ�#���y=d�5;���)!=X���Q�<���Mx=�h�<��=��:"���;��H��8�1��nΘ�HDl=�)8=F:8=�๸��6��4=V\�"i#=rc¼Cէ��b�3ڑ�t1K=��=p�_�ڎ��B8#=ӳc9{���UO�<��~=�0r<sƐ<���<�O(�J4�;`}(<
~E=O4l=��=�8{;6��<'�;�` =xA�U-=X=n�P�h�<��<�LL<��<��:�*=L:=��Ѽ�@N<oH=<���;=�@��\�*�n�ϼ�y=ы���T�a=��r���*<*Nܻ��=T��.=5�V���
=�B��r	�g��|;�f\
�?ؾ�U��<H\�b�=�<˰��8><���*�<U+�P)����<�:�<~�8��j4=d�<�@�<X�d:��n�.P���T�ֿ����7L�	`l:�)(���<߯�<P�S=��I<�Y3<�����7<m[�<�EH����;d[�t�@�|Z�\���[�����:�9B=��=��O��_�<b�t<��<�~=K0f����<���<ԯ%��0��7=$�L=��2=��R<)n�<�= <�`;=�C:���= ��F�<��ռ�Y'��0#=�0�����=F�2EC=��~=zv ��Y�<� ��G>=��:=���<�?3=�]��_�< ���[�;	<Q�F�P}�%��@���N=nZX��/�;�B�<'L�η-��I=M��<:���\6B<:��M|�;+}�<��6<=:�<(o���f;��U=&�<�qV='=�x=����fA=D�<����o���a��*i=N
�<�T=7^T=̨<]�ɼ�=�-�.�I����<�N���<9�i�^���K�
��}�P�v���1��-���7���Y<A`s���S=!��<9^=�ɬ1�������ɼ9� ���^L����]=�<�>��I;�`�<��׼�`ջ�������< _%<�d�<�O��k��<N�F=~��ٻ�\�<��,�!K�;H�N:H�>�CO���3�?�v�����e�<�N<7��;�n�<�\/��B����E<�V��"\<�}�<c�<+�Ѽ,b��t�ܚ9�5�+�ޣ�<�i��wZ�����<��!��
�1�"�A��<�ռ�r�<M��7H�<I�=:�S<���)=���<0���/
>=S�;�#�{U7�X=��=�X�;�Ћ��B<�9�ǘ=���<#������<#��;����j<�Y,)�	=��M=|��;w:w�� "��S��(c�i�=ٴ�<��=Fu0������;�r�<ɀ���س<.��Ω<�E��2�U�U�-=�hk��2 ���:q旼��ʻ��C<�V�$HR���7�Fu�<��<3��� ";��
=0�y6�6l�<�#�[<����r�!=8�=a�<�µ<z2,�3vټs�<��=1�ʼ�
Q��d��|�G;"jԻ1T�Rq="�#<t�?�k�1=#N� =wo��===^�ӼX̓<�3G��h`���=-:N=�CT=)�<=}T�*�=�#�����ӥ���*<�H<N��a1���<��m<�C�;"�=��<���<{�2=ʓ�=K`��z;w��
=܅=�F;G���PQ�90H�i�=��R���ϼ/�ټhj��<�5ż�_C=�`�<gq�<�B�1)=��߻�`8=��:FW�1�<�vļ#�$��<����N[E�A�?��bN��a/�LTR�= ~�7���c<��)=|�.<*���==��Ӽq;R��܋�����:<��=�;B;N�:�p�&=��X�=A�f=j
�Q�a=@=�&>�t��<���;��-��A���l�<`�����H��}���6�<��<��s��=d��<�G�t�>�U|.=6o=w¼)��<�w�r�+=��G�m�~;��=ϊ�C�=�.=�b����= `�;�8A<>=��wn�&�����<�ȻD� �[���0M�<�=r�<v{�<Jpּ4}S�_c�I�	=4'�<��<wE~�Qz<yd�m6f��.J<zǧ<�6;�!�;�<�)=�!��8&����:����N%��d��媪;&I�<S.�<',��Q�x��
 �ںk��O���*=�:=@g��}L�a�O=嘄����<{�p=;$t�}'?�u���F��:����W;�I=�U�?��޼#����i�<�L0�nj��oG=��B����<�L:F�]���<X������G|=��X��i9=|�&<:AĻp�{�~����$��x=a����=��z�8ϼ�	�9����<e<�܊��7A��Y;��E_|=�����x��/K׼W���$����<`=�S#<ԫ��i/=DL4���z�M=*c���#�`/=�q��K��<��Q�榼Jˎ��L6=�Ѽx%��~=��5=��=���<�<�=���X��ՔD���r=�xQ�J��<��<�_:��B޼Y�ټ>9��-��7��d՟��ʄ��F�����~X=&�ڼ�劻��c<Y�<tZ*=���<�
������-�؂�/���4�<��:�L�=�GY;�q;=;�\����;�X>�Һ?=��%=��k<1�=	�[�#����5C���==�f�<�h�f<�S ��x�<�l{�Wf�N~<�R!������Xջj�<])�F�!�LN�<A#�3�K<���+G3��=�sݼY�^���V�HZ=�:d=uQĺ�}ùU]=p���8=��<O*�<`�������=o�<���<y��Ȱ!���)�N� ��@<���:t�;�N.���4��O�;�	b�C�!=�C<�/=E���L��v��5"�< ���޴<IU��ao0<��=/`�����<Ge$���L=��;�[;�29=��鼙�&<�m��~�/����|��J�<��7<LcS�*� ��퍻�pW�1�:H=7�L����;L�=���<J�8=�
�<��d���.=}�i�f�ȼ�:��h�<�k)�B���g=�q���=�u�l��<
�O=`���!ɼ�H���k=�+ �x���o� �Fg=�]O=\�o�u%�9:5=�,�<��X�	��;hR�=e�B=�$/=���y�"�n�D�w4¼�c��I�;3��<��Q=������"<R�4=��=j�Z=r�a=v��;��W�k@�2�<U�#�8o ��1F=
=�2��ƅ�<�G�;��<.e��k��\����E=�ձ�pPN=T+�<�M���J=��a=kN㼜���uT�e*]��l�7n�<?!Z<��<E웼����n������ù�79\����<�r�<�&;{���730<3�Ȼ/ز;yw��?s����<��U���h���a�4}H��)Ƽ��<=��.8;<!1�;����1��R9���<f0=s�q;t��12�;D*���D=�@D�\�w<o�<��4=,m�;8�+���4=�˲: �<��,� �ü�of<�F�1Jf=>�����D*z=�ʷ<���<8�ռe�T��%����<7;=)ī<�:<���C^�;S|���nV�a=�w!�����i	=��M�i:�=���pȼ��A��A��[�;�=0��<m����=��s�=���<�sۼE��<p=��&�w�=�a�<�<�$K��&8�̅^=�=1G��|N=ʙ�<ȳn�WNa��� �L�I=��N:T��<�yf����<�0=�{�:�22�S�<�! <q43=YY�:��;�9m=�>�<���&zL�(=>�ټ�-��2�`���!�;���<��<`�=�l7;��A���-��U�\	.<\Eb��O�TU=��Ҽ�^P�7�>��ɻ�:�<�]�z����9<T|ּ+=�L<=p��B�)x��<`a=�(���>:՜,�`]�<�
;AJN��}x<��></����8�9R�FO=���!j=�O����<����=RǼ���<�7o��pY=w�5��M=W)໣�/;���:IB0<���<�Z�<�E�lͼ�0�e�.<�:J<�N�X7�<*����|~;I�+�=r�
�N=}e%=`!y�j[�L��<�7<2+=	Y���Y�`�z�ȉc=�0����t3�-��DqS= �#�ơ׼ǼZ���Fr<�RB=]MB=/���7d�̿!=�?�;�<37=���<�QY���'<����\�2��z�ܵJ���ȼ�&�<��:=��/=�D=2 L=��=� ��%#�_mռ�l	=mi =�x�<N��<ZK��<cj��:쑽�2: e�<��A=�̶���<���ɼZ-V<�vF��<��a=��T���9<b�X=�1=_�D;u=���<�(�<f�{ Q���Z�ϼ��<$�<�~E�k�ռ�^�<��ۖi;�Cl��/=u�޼�$�<ׁ༶�=+������SX=�l=��f=���<�}'�E7K=�g���ZN=L/=QW��;";� �;v|ؼ3Fi�c�<�o�:��B���_��g.�6��<U(�}��<X�=��=;��`�r@�	�;8~I���<�*}���<m�5�R�z=J�=�;<���'\#�I�F�#)��U*<;���CS=~]��/_�\���/z�	h�n�:��B�uua�Z�[^B���;�28�"=s�T{'���x�c����<hn'=���<@�ݺ���$ں<�,�2l2�%���pKt=�=K�l�c����=X><������f�.df�5�뼓y���2�;��M���ϼD��<RV��[= t�<9�=����&OM�R�Ĝ�<0�9�ԕ�=7��~���B.�p��o��<!�<!\={A�<0����o=eI�'���0�<���<sdg��ڇ��%��R��8��0�A�������S��u���I�-���>=�o5=��ͼLv�<v�h�~m�<*x��sc=\e����/�C<� ;=W]���58=A�纅[=��4=0�v<Ӧ�<H��<���<+DH��,���'(�<B=��0=�r`<Bs��^ ���\=GS�;܇����U�A�­�<,=�?�<���<�&�<�J�<G��<F}S;��C=k ��Z�A=���kG^�`9�<*�<9?P�%D;=3j=�^ؼPH$<R�<=��=Y�ӻ�U=u�%��8
=}�������	&=9�+�8=�}=BU���G=K�(=��R���S=�q�;�C�<��S���.���<�������#�E�Ɋ׼�_a=4�q=L�a=|�<m�}�d��<J�:�/=T�R�1<��#�¶�:/��˭��
*������	;�qP��cC=���<m*y��]����W�=���V�<�����?=�-3=H=	��;�ON=[:T��䍼�G��J���i��ժ�{p���<�E�<�nR�C�	�C��<5��F�*�޼�T=��&=�n�!o;��<��<0�#=U�K<���.=�&K=#jܻ �=�x�<(����������=���= ��Ր<�
�Y�6�'7== ��Rq��̔=@�o=�z3��(=c�����.���I=#�;0x=ѹ���ل<b�@�';S=����gD=i+@;NfD;�l�<<�m<
��d��>��3?�@o��pK}��v�<��0�n�<W7^�;�ϼ�l�:=�=��_<�
�b�;�eA=V�;;�/��E����j���1�������i�|�=�]$=�J�s<ȡ-=^_�<�����$����f��=�<)�ȼQ�'��=�>=PV2=�=�;1�.�b���.�_�����<�=�%��L��=�H�<i/ =�IļL�<yy2=�i��)�<(4X�/���*(��ͦ:�� ;�ؼ�o�<�К�1��x��<�d�<M=��R=k��<I�ۼ���FS=_�e�b��<�bW=;7�;�$C��=�
���$<�T3���2=X=��N3 =�	�<KC'=|ʞ��2�;B�9�iF����<�D	�������$7=��<�+`��פ�2��;�3e<�����<�%�Pͽ<�ȩ<o��=2�8���<��d=L5���D���<G��=��M;;� =m.����\=��i=sم�*@=DAj<z����;=���4�t���d=�D�<��E:����_=�:���;�x|1=��=��F=;׮�;D%=��<g�M�i���q5=��<^p2��h=������
=�}�<W�Y�� �<=o;=��d=�}�A�P������m�� =-�ϼW�a��PP<��~�N�?��Q���/=_p�|��<��<T1<��J=��4=�T=~ݷ�7�	<�U�:�'D��96=�����Ҙ<�gU=�_��":¼7%��f�=@,=���:-���N(��N_=��-���;���L���������@*M<L�='��<\�����1=�O�����t	/��z��Jq��D���5�<��R=$9=BĖ�"��<�zT��?d<�]k<J�<p�ռ\E��Px=^��p�	=h�9=�n3�w�\=�4%�Q�;����o�=�;h<Z����:6=��1=r�3=;����h<�=�S�;�BP���<Ħ/��+���Ӊ�<����[���id ��,s<�7z����;�v%�n�����O�rR8=�@<�� ��<^�I<��%��]��>=m�=������������<��<����/~;�Fv�}F<�	�t.�=޺�W��j�<L�/��V�[�@=(R�<(����/�������9=���<��9��z ��Z�<��]�	=�>ϼ�QN<a��=�rỾ̼+C���
=3i<���<椱����������<��K;��\<�2�x?�������D~<�y)�vЂ��;=-�c�x�/=N�;تм��	�9�=�GY=a�P=W2�<J��gN�=̽�<��S����<4�ܼ���<[�;��/=5�"=E��8=�*7���!� 9=q�= C��P��<�lE<Qc�<� K<��=^л<U��<��=�"y�!��<�]j<�j=�t=��<G��#=��p�.ۧ���G�t��<�{����;U(��E�<*_���=A�B�Lʼ�{Y=wz��r$=o�w��̂�Ӽ�:�sK.�<�6=g$=�N����[�|ֲ�9Ux<�̀=��B=�ϼXHi��1<�29< İ<��<��"<|����lX=�,�<ŏ�=k��EW��N K��UF=ˠK��L=�uM��磼}OC=):!�`��;Hc=�X<�H7��T���M=:kA��[����=��9=���<v=�w�<#r/�6��<���'��<��<�����b򼀵==�����<Ws=�|�,��L��-��$!�����=��)��P���*u=�Wͼ[,�<��J=�z=���k����=�"Z�?��9�����3=��k�y��?�;~7��MT%=��=;I�<x��<+�亵Z���<��<q� ����:/WE��������<;��<�I�c��<`���:M<�x�A#�"*J=�N���=��g�d=ǀ���8�[.=�i=R�C���T�s0�9�;��y�N=�u��p=*��<E�4���=jp+=%.^��b=��h<�p�<�Hb�Dݕ��ny��,s<�G�7�=�bD�+�o.<ߑ�~�i=�_5���<n��<�$�;6�ü-F��R�伩'����=�m�<���<��b���==�<���;5�ؼ�=M�|�J=�����Lb<�+=� >n=/�=}Y�<ʏ��s���y:=]Z=�.�e)�;��f�S�m���߼a��<꛺���<���=� $��p��F:�eK��S�Vż�;*u��{���<��rR;��=k��<�����m��;��<D���ϼ�)��7=9�W�������{�޼ԻP�B��/���A���;�Sͺ��7=M�u�K��<V�Ӽ�F1=-�7:���q��<9c@<.u =׺m��`=�6��Wn=Rl��ݴ;�!�������)|;�阼�]K=�P�C��$k����s=f	���l= #=.�Ѽ�C/���a�����!M<�W~=0*�<���<5=&��<u�<��<]��<��a=j�!�1���i�-��M":�6f=/=��<Tt=u0м�\̺yD������ ;͸b<P�=�3�<�Z��EQȼ��=�C$=�[�;��J��
>���>�����8��[����x=�t'=2΃�R1N=XX	�ѯ]�V�c=������;��x=��<%W= ӝ:l$��4�E;9�<CX3��`��X�<��,�b==v[=H�ͼ[iZ��� �� �<3��<�E<��;;JA=� 5<���<	�d���U�k� �%=����4̈́<��ڻ_4�:4���a�J��\� @ �b����=(��<,n����="�����;�SԼ�*�<���<%]���5=�H=[�j��V);T�<Y��bżP<aڀ;�uw=f{2���:=W���2���zg=��ɼ�Y;RDw���0�E)=iB:����x��x<�1=	���l=N�3��У�=|&=+��;g�=3(<�i'�K%b=u��1��<��R��	i�6a���(<G�V�[#h=�����\=�I<,�8��ꉼ@[=Q�$=P�l0��O<���: sw<�yQ=�NM��zO���Z��M{�0���,�:�R�rz��O_�I=Ƨ?=�^Y=#���a�o�~=�D�h�k���9�Vm%�c-��[�I�ڼ��,�����Î<(*Լ�~;&/��s�<�f*��c=��ͼѷ��t��_�;2=��|��-<DT='�<���c:���;�sN�[��31��`T��jb��2�<Ê'�m�[=�����;= <�SE=���<8u�<Ơ?=���o5$���$����<��l=Qq�<�;�C�<F�����q���$�=�;w<	Y�vb���I��h��!�Ѻ�d���=�`0<(U���*��`9�(V=�c��w��<��=��=��$=,���؂A=��R<�z(=�T=��=��M�E=��&<V�<;m�=Gȭ�s��ɔ1�M��<C����A���]<�H���&m:ˌO������k�ʼޠ�<�=��޼Lh��=�<���h�+*���<nv��(�]���!=	*�v���V=��	=�ڻ��;��2�-:�<�a<�/I=0߃���^=�1�T����R��2<�%=�}W=Z�R=���C޼q>��ZQ=L �<���<��=�&"==$W=��켪֠�2k==_�Ӽ* =���<С=���<Ҷļ�"�G4>=Z�<�t�<m�����s<����Vw=̍c=�ֵ<��
�>�"<�짼�_��� =Tj7=Τ�����y-=��.=B�u��m!=��;l9��Z缕��<o��LI��&Y�/����j'��t���<j�=p�=��,<�J=[ͼ<�%�<�o�<!D�<��F�����a2���C<�f=6f���)}��YH�W�	=����#0=L�)=he=���f�J=Z(�<*���^�f�ټ�n�=	�(�ڻ0�����=�/D�/����p�,ſ<��<+4|=��Ҽ�0�{�ټ'e�<\�<l�{�Nm7<� 2;ɹ6=�عU/=ҫ�;�v���w�z�6=��~<��=�_:`�,�	=�9;�A6=��1:&��=�i=�"�"��<��V=��9=��<WG�;�U4=�W���EѼ�r7������c=ͳ�;�=���;U}<*��Js�;�o�pf=���I;ҳ���f����+G=��c=&�?<@m[�G�v=� *=�_�;_T�1
=��#�`(:�|���=|�"<C�۹�Z=�����<��=F�+�D��]�<�����T�;&�q=۝�;��L=x.���_���{ؼ�c=��Z=R������]!V�ՐJ=��R;H%Q����<�)�<�s|=�ɇ����=�M�
�-:�FS<$om�ln�<�z���]�q�<�i6�?�������9Z�+��̈́ =�Z���;=���;;���` ��_=ޔ9<!x.=_~��T5=0!P���̼ڵ;��K=#p <��'���3�Js�<A�� �P<;[w���<ͲH;�Y��~����د�Ww�ZO��o.���=��]��ؠ<"�~=��<���EWH�n.=#\�[�*��L��V��/�<���<ξ<iU�<
9<��)=C�X�l�;�*�<����<q�u<�Iw���,��<=\:�|����ړ�<: N=2I<�W5=.���pE=���<��1=�`y�f�=��&�r�<)!n�9/3���<O���7�<�Q<���<Z狽p���]0<#�b=֣�<�(V<��q<�FG�|�<��F����;�H�z�=���<�. ��J��� �3�X=kl�����^=/P9=�Ѽ}x#�^1�o���6#=�k����:Sp&�t�i�.=�`��G��<t2=�k;4�=�e<��S=�;�~D=!"�<�M=�>���:�J=�c7=�3%=r_�N�t=	|==�ͼ�BZ�a�4<K����x��Ec��)=_=����=&�<d+,<R�<�$���ͻt�i;���R�;�]���=�r@�{�=���_�o<m$=��L=]�/=o��B�l��"���B��`���кA�=�P=�8=�<�<u�Y�����
�?=�4q=RoV��m�<>^�:��T<�ڴ��{=�[��>�;n�u���f=P��<�Wϼ�+Z��o��,�<y����0=��N=�HC��n����U"s��/¼>���]�<�`�<���<�s�<�A�:�=L5�<-O�;�n���0�EV=ej(��=�;A�!A��G��׉��z����L]μؼ���*p9�9�a*B=Ķe�_�;A�
��}�Hke�%�żd��]�Y���;�\��9a���==f7��<��5��<M�;=_==���������<J`�h����S=z�:=m:a=E�V;Y��<�B.<)��n�x;v�һ�N%;���<��$�O�Z=F;ܺS;/x�;N�D=P��<%=���Xx=�����)=.O�<�P;��]=���<Ѐ��]�<XTa�gV=Z�=���F�=���k�e�$�"ļ�N/�ц6��O���\m=z'Һp�.=w�=���^��\~������=zW�$d;Jt
�O�1=��$=�A=�AI=�x	����<���<+�����r=�<�Y���YӼ5��"vI=V��<��+=�VZ=N=mD=��G�#n<Jƺ��$|;|���8�b�P=n �<F��<R�+='��<�h=�<�<�:T��T�;����SA=��{<�A����<��=,�0=�o���*=��=N�^���h=��/���u�X=��</F=_ӼOL&��P^=.W6�|��������<�=3�5�%�#<�0=J���=�q�:��<oL�<v�t=6�aK�;��9�{�<��<n(=c�<�>)=�*�����<�м[T=<�������<�i��X;�j)<�d5=�=-#�n�[���<[�q<}n=\�k=��e<�>���V�y܀�#�`<���<����G;�j��E��<�bS�K�<�w"=��b: �ټ�/ռ����t�<"���(�<$��d��<e�������\T=�0���潼���;!	�O�-<���=I�`��v=��X��9c�?W�:n���y=�Nμ��Ѽ��r=WG =��Z=�"��^?=����P<�%,=���+=�ꢸ�'�~�+=��;��=��[&l�A'W�Pݘ���#��P����ɼo-�<�锻ѧ1��*��'��̸�<gU�<��9Q;���;:�����ɼP��W�E�����[:���<��Ի2Nj<WL�J�<�B=�$=�A<�Z�7`M�~#�<�=(x�Ĕ;\]=>U= �=L��<oe�<j_=�=�[=�7�<sN&�ўy��<���?�w�W=��^�L=��1��V="�l�H�=�a&=(��<��̹yx����p<�$�;dP{<~�<>�C�e�(�{�=X�^=Cd����<�(�<'�<�=\�����<�-S<NzI<b[N=\��</d�jv�<a���HϼP��<"N5=
��p�=�=w�ļ�h�� ��<h��mt�)N߼��<P���LB��i<��	=�Z�<���؏8�٤�<@��<��;��<��=���97=р�:�Ȼh6���f_<��ɻ��;%��~� <�R ��X<a�<k��ek��$B=wjG��s��g8��g�<��;��μ�A{��*`�G=x��;����|�;.�:����e!o=$��bR=��P����<y�)=��n=wu|�WΗ�|W<�b���/���a*��C=��%=�z\=ì<F=��s?��+üm���<���<� м���<�\��ѻ� ��.x�'��,�}=�0,=f=PEμ���_=��N=#K(=�.�� �=�T��ji8=wqG�D����1���[��<
�3��U�<�5=�pN�8(�<o��<�v�<��U<<�}��缈�'�'6'�Ѵ�<j?;=������<� =�.�^F=欁�A5��"�<����N=ŔR�\��<�I�<�y�U�k#
�p������HW=�L[�q�=��3�wA7�r
C:˾��co�[�9<�+k���Q�������1���=�M��i��ۻQ<	F"���=Y-<5AE=�[���-<=9�<=��7=.	S=�]=Y7�<`[P�IS=2��1���7���C=��<@A�
 6�JUq��ѻWdO=�f�<��Լ~{@=��ѷ�bu�;Z�$���7�x��qѲ�|�c�]q&<ȿ��P̼w�$=����L�V=f
�5g=V�u=�<=rۺG�=n�;��<�8=�8���&=������'=�Cf=�?�<l2>�,dQ�����=�
=��=@05���+��㥼dw*=�u$=|ܶ<� ~�b-=��L�<���Qa=����<u�t���G�Ƽ�N-=joY�]�V<ϵżp�̼+XK=9p#=��=sgb�h �*A��X!;c�O�x;=�����K=
;y;ER7=c`=�00������鹼׷g�D�q�Yh<�&) � �@���h�M�==��<k�==��b�s�����><@���<[�v=�CA� V�ϕm��X�<nXܼT�J<тg=*��<q�~=�pT�9�M=%�[=7H��:�m߼g��<6�p=�L�������溽)�c�=��'=��l�Sh&�Mg=�* =)=��=�J�D��~��q<���<�J��,R�����۽��Q%�Q��V<�м���<|�W={���<�-=���=sWȼ�xK�!�B=~WQ��_�;�M��t �5=�r<_�J=Q7�=�N���<u���Z�Ҽaǚ�� �%F�"V�< �_�h0s��Zl<ZD2�m��0�$8zo9<0M=K������@�����<BQ=$�k=�Y���N��J��]d�y��<|^�<��,�4���:<lY�;�=�/=n�s���y��-�r�=I��<φ@=�*�<���%�<���\�L=�q$<ˡ�9�� ��V�<�H=�4s���T�bng�'2�]0�.p���\<p��<$<�<��<�l=�%���><2&*<��j�<����~�
=��u��?��'�=�+#=ۘ#�5�4=��2��9�<x�HE��=��_��2<�f�<ї���U�3dA=����a�:)�λ���S��7B�<<�W=׽8��j��x�<Z��<�n8==^c��P��or�L�ռ$�<�V>��3�<��v��U�<���<�TӼE�F;�	>=��d<�=`����B�*�`��а<��>=�K=8N���&=q�h=���<+�D=B��.�>�qhK=�vD=��=2$=�d:��<�1�q	$=3B��h�<�7����&�FE���<M=����)� �@��<�R��|T���7<���E�=�\�y	8�7�<��F<W�"��<�Y&=���;�#=Ů>=��M=>��<3��b#=��;�`�:�)s��<%=�+�<O=���-�<X��� X:;�=�n��پ��Z�s�^y�<n �=�&J=�7�<[�*�a�J=���ި�<s&�=[}&�h`=��@=**n���4=4�%��g�	�F=v�92�=�1�<B����+���v�j�;�v�;�3v=6P�v	=i���/U<ǔ�J��$�g�e��"��a]��i��=���;���;ۻ��^�%=�Z{<�-��� ��0c=�W�j��;���I�缈.\��,�;lK���?�j	Z�_z6=�fL=��;i���ƫ<�4�Ms׼7��;!n�e�<м�Ǻ<h5*=��N�9G=��<�y���<�<g��^��a�׼�$ͻ���vʷ<|��<�}����<�X�<V�=�9������<�%r�U(��O=l�)=�}<������f߼�;be�
��;Y���M=oU1�*�%�}����;��<Ҽ��B�aC�;��<�D\��=�L*=:�����A�%=�,;�Rf��� �#�e�<�V��GB�}�ܼ�D�<�rm����6��<����)�ox<�ހ��0(;��:J�%���i��(<�6n=�B`�э�<�@V��/8=�/:=Ê<���<�=wԂ=�Qq<��y�Gr̻���<�n'=xB���;��=5�<rH���3��s����`����:)���Y�<�X9�>�<��^�R:=lB�<�܀��\+=\�	��X&=�<=7�<���;��=��"��=�%�<"��<W�<��r��{D�{'��n�Dü~SX=�Eo<,��|Bz��ʹ<��B=8֪���Y��
�=;�g������yU���#�ғc<�B=Ʈ1=�� �~�5=v$�<���<+b�T>;�
����q�;�k;��ڽ�~���6��=�N��*-=�!�<��Q��H)�#LB��|/<p���7"=���g"�丕��p=��T=(�;=s�=��s��O�����eR=�{�<$T!��S{=
a�<��*<h[�<6�$=Ad8=�X�<�݁=�ے<�1c�As�:������w�`�b�Z=��L���!<+�(=��:�
e��l���=����r7�\�:p(�<���[��<��,�G�=��;�gh��ԑἪ�ɼ��l�pzB���K���,��T�$�.���u���V�Nu>��i�;��ռ(ȼ�	�;��;�k0���<>�<=d���#��5!<Jp�<�f�=��`=Z%=��j=c=�V��^ɻ"ǵ�dwJ<�M߼�\=��,���K=�d�;�S�<��\<�R��ͻ}�6<�=U�D=���<�dG�'u�;�&<9�V=�U0=`�<?��n0<ƪ#<��S��H;;�CG���ݼT�ּgI��Լ���;�<��������D�<	��:b\5=�ռx�=�4��'�<��<3N��\"=B�i<o�;u��7��<Z�O�a��<߲ؼѠ=��<�(=1�ٻ�l�<Y��<��0��KY�u�;��W<s�t;�J�7a���1�<�5 �ΰ�5I%<��'=���<[��<э �g�;_�<<�(���پ�MZ=#db�UP <�].=s��*��ƥ���?<��<�����-��Iܼ%�C�1�,�Z<�2R~=�S=�8���¼�.�����<p�H�$�ݼ��D�!74��TL=w����+��H�;B��<{���f2��������qۄ�2�z�N�c=���<��z:�H�Ɨ|��hm<ZQB=�漼�*=�����=ᦣ�>��@n�<�w]=y�#�˳=�Q�/�S���A�=_=��s=��2����<>0�<��<���q<��1�*|U��q� �X=�N=�l<s��<���D����=�B����<��#=��˺�lQ��]1<qO��
����x���f;ѥ~=iQ�.f�Du<>^S�$�=�s�� ��Q`L=Ǹ�;^� �j��Eἢ�,=�bY�� �N���x�=`q�;�sN�uJ	�I�;��5�`~X��<L�I�+9�<��=rR<Kt%=9&v���3���3<Zߘ<t�1=�A�Ǖ�B<(�="�H�8�f<��<VC<��Ǽ%�Q���V�p�<�=w�B���{��g��Y�E�@���!���@��DO=
�L=�)�<�3d��o�����xϼ�K=�rJ<��=:��[;3�>=FZ�<l]@�U���Q=�����|���c-=7	=͒� (�LSѻ����s����4����K�L=� �����^|�<���<A��&�=��M=y@��KL��8�g=K�=���<�X<|�N=;JἅoQ:�fp=�P�]���6x��
e�:q��;?v���t[�����<v��p2M��jk��`=�9���$���T=�~@=�'"��&��6=1�\<��<w�;w��y2���GU��J漻��<.�<\�
� ��I�xZ��m?�����Z�k&/=ڼc���J�"=j�R=�<����=�T<���	�E�{�;�l���vǼդl==�h�K�;�>|��w�<��;�&/=]�Ի�'=�sa={�<�5d=�S�t��<���3q=l@��A��qG�<��<϶߼��X��崼Y��<�<6�<�s�HOI=u��9�k���O��K弯P.=fk�
J>�w�<��,=zn��X�;NG��}}�S`=�QW4=�Jj��fU<��W�+/=`Q"��s�<i�6=��ͼ�	�<U���y�����<ϝ��K<���b��WR�=�<����Y�<d7<NH=T�$=�^<=�%=<�߼_�~=�n`=�����;=��R�VT=��u�<���E�R=��� �<[f
��<_\���LO=V���ܪ!��S�;�`�<\ �<f�Ҽ�4==�|X���;=6r�<�4���E=�<ܻ�:V=Q=n<+��&�N��<U�<�#�iu>=�m���e�<�Ӣ<qt�<�%��2:�'@l����;ѷ�<��<`Z�[S��m�*<���<q�?�7���E��R���-=���iD<lSV;�"&=LVp�?�<|�5�Gv��^<���V�W=���;�»9�u��D)�<\�<�5j;s=?��<
��L׺z\��p=��E=��J�8�=W
��%=��>�>��pW <�"<�M�;�ZJ��nڼ�n¼#�=\�#< ƻ�f��)�<`Y�<�"�1$<�ۉ���:�u�<×�����<47K=�=˼�<l����.�j�)=�U�g�;�ݚ��wS�o�o�?0,�,g=7
����<�W�<�^D��UE<x�c<�X�<;�=������'�ZM�<�
:9�B�xW��Q9<���8�;<0��ى�97�=�H�<�p�T���W��:�@��Իp�b=�|?���༉O���u-=隇����:�8�<��J=�	��A5=�p�<�\��u�<_Բ������<4�<�|=�<ܻ���<�w��ff=.�Z�r��Ўx��K=dQ��b �Y���=:;���4+=�M�<~���$����-n�<��f=��<ד~;��M<�ܟ;�/`=<yA���<���
<LN=T��;���;�o�ReU=?��2�����_<��޼[ؗ<@M�J0|<���P3��� =�5������<Ѡ"=O�5�D�����6�y���@|=_!{<�E���ld=�<���<v?=܊���w�����M��=ﵢ������g<J�Y=�A�7B��5	<�Ƽ��H�H��4'���ܼ�>��]H����<��={uG=<�;*��<�5Y<��><MD4=v�s=��Q��D�<Y��EȪ<k=<��<]�U�c�=4�<����7A<� =�� =��&�p]}<�e=�Q5��F��F`"<�=�s�2�=���3=��n<7g=���<�y�<�Q�:�(�-i���ؼjơ��r���QM=Y#�bNѼ�<�ٍ�R��;�iN��S��X�<��E�[�D��.����o�<��ջ[��<T�=	L^�	5E����i�< +�<�f;)h0��',=�]=+��Uf��Ds=�N�<G�Ӽ�B]=r>O=F���Gy���W<��q�/X]�-=�?����-���g�+�"�ܯ<֯8=���,��<{XU�ALN=��=�#=S�f=A��CI����;z���������=!:�9$���+�=K]=�T����=2����k<b~�<��;)��Mg�:,?u���=U*h=K�O<���6�'=�?<�W�8O�<e;!=r��<���;��39���;�$="A<{�;�+=��%��؊<£`�kX��7�6=nn<��b<�S=��ǼqK1=��[�!���<�\����<1����ݼ?�6=�:=w�K��<���;x�C����<m�n:˸�<��=/Tw=A.��<=PX��^3���/=}�
�; l�����w�b�^�\<��&;G����l��Â<�k�v=++�;�Ɇ�Ԍ<��+= �'=a���-���J=��޼���K���p<
���F����#=�4��%K=U�м�ٶ�&~��9�s�?��ދ=�.�<�N;^���R=�ڼq��<���~�<*�6�"�u<���}�;�������_��<j0-=�� =�߼90����<�iּ.qB�>�w=���:%IR�X�8���<��l="�Ѽ��\�{��.6=��.��ػ�"=)�O=�U��=8�Ē�<����=ptN=��<��A=f_�;�P�<�q=J��;��3_�\�!=�}��8�����<�nx=4t��� =3��R�W�J��x�<���w��;.~:<�D=�.=ˢ��S]ϼq��:��^=����U����6=V =V<���<�t=،M��k���`�Us����<b�=#�=�꺼�6���b~���#�x=� 3�bY�<I�7�運��!=�v�<��B���6�F�"�:}ڼ{={u��K={�F�N�2�j;XJ�<i43�^��; &��f�k�~�<T�s;�p7=���<�L1=ը5���<g=C���<;]P�N�|=���<�Z���Q�ń�<	��,��yu<�XB��uE=�1P<k�S��a�<f}O��#H=���!�̼�>׼ߔ8=��a�j�V��B�t�H=}�&�i� ��%��;��R�=cvD����<�j9=��<��9=��q��]=�N��yi<Fe�<v>��� ���<Z��=%6�=�G�l����=d+�pB��l0=u��<1�Ѽ�@P����:�X�<U=n 6=���b&=��I=NB=�u�<'v]=7�����&<�q��i��0�<�6������>���}k������m�G=�Ũ�)�5�?�;�q~=D��=<U�����vp=�}=9�F�X�'�&���� ���<B��;6����7�;D�T�O��:��</䖼i����Օ�bW�<�� �&�<Pq=�a=$���P��<eu�G'��(��B�:<Н-��ߖ<�ƻ�jԻ'�#=b�=�v��S�\=9�f���+=j=�rG�*Z3��Z�p�+�4=�8�P®�8P�n�%=Vvk<>�T=�3w=Na�;�e�7����3�8l���a�s"����=m?<����J���J�3û��;�J=���Av=�#<�7�*<(o=H!>��<�Q�=mr5=�L�<�5�<�m�<�PI���<��F=�
.��:�ۍ�<v�2��,=O1:7�Y�I�(<\1伇'�t�L�^�̼l]=*׻'Y��<�;"�`��@�DP���)=O0
���}�^���<���a=�JK=�a��
|����9U$��q%<�<���;Vu��G���m�߼h�=�j�<4�=n��:Ђ�<9�F��w#=���<��x;k*X�h��<R�˼Ĩ���Cּ|�Ȼ����^�<�_�<�W�;c`G<
��<G�=Ɨ;�����=�z����;%~A<������=^���5�׼/�����Cct;V�<gP��S<��=�ټ�5�<��D=�ml<�7d���Z=���=_wl�@��<k���y`�<�Jo:1����P���%�LC�Ys<�.���&q���,<��G=A��:!&�<I&��55�7��DW��o�')C�9޺<z�;6	R<�&M=��J��=�)����"��$�Y�U<�o?�; =_���3��$@��㧻�.�<�=߼U�<�ü��9=a�N<&��B{Z�v�;mK#=��=���<n> ��k���><eX2�V
e=�~+���h���<%���_��F&=���̧��Y?���=~I�<��:�az����<���Ӈ=�� ������l�c��Q���.��(K=��<g-|��+�<Y�ռ2$��[�;��<�rU=P��<Q+=�l�<m��<�1�Ӷ���ގ�lb=4+�("A<8�h=h��<���Si�:��U=uz=�s7�K��s��<�ӫ���==���(�;@�a<�,9=*�/<��,�#�<}�L=kS�Вf<�P=��*��@�� �:�b���=^!X=�8�<Hy����Y�;�c�'�Q�S`�;��=�5�k}<E=��.�<(�;�p8�u�<�u=k24�"�����=H���<�D L=&�����><Y����<�� <]���l=�P��#�6����;#/Լ�T=��3=�]=��4��1K�%�ϼ�l;ȁ>=�X%�����E�Jw�=N��=Ɔ�:(��<le���O���`�<A�,�+�G;߯�N�<~�=�������;�o=AG�<F��<�)#=�.���K��g'�2��G�˼E�S�w�r=�Ӕ=�Ҩ<���<���o�W����F�v���^=�<)����Pm��Q�=9�?�^y�=�yl�i8����=2#K��D(�V`=uv�<�:�XVf=���U�S�ͼ�
"=��l�F�7�m=���;�*��B�=:0 ��=0�<�B6����S)=�@;:�Y�6���W~��R=2'<�<+�����8���<�a=����`=Dv��H=a�=��I<8xX=�=T{� �-�`IX���J���;�a��;n0��ݗ</�j�;,�<L�K=x��<")<=��/��=��~����<�o:<�H=����_7��o��@IY�*n�얀;#�!�+B�zo<t�2��6�<�~d<�ּu3<��Y�U[=��;nx�<�ػ
�s<cJ:I=��=#��<s���ݻ���<�=X.���j%<�[= �F�:�=����/=��?���$���^�r���%=w�F=b7�9��=��^�ш�<=Jm�E=0;<�C=ɫ:=	��8Ct<��7=�#V=I6;�"=�<�<���Y�'�4�S���\�K=�8=$�x</��;���Ə��$�<�����^�d5=[�ͼ~Ҽ����Y�>;P�� ռ,I7��T<Pj��q��xK=FP[�����D������^=�&)<B�<�[��E�;k�=�F���ê<�s2=z;�](����pYݻ�"	� ��<��v��a����0=��<�=3�<�N7=�Qn<��:�d=���n��<^(<��_�g=!ˋ�qq����1=��i=8�?<�>�<U�6<R���Yy=�:/<ɂw��[���"��*o��,ӼvZ=
��Z�ѼVi˻L9��p_�<�h{<gqi�a�n���[�<��a=B���{�\;�.$=L}���7���c��d|<�2<PJ���(=z&��)�:��b<��\=���;b�>=ò"�\�(��i�=��Ȼ��=ͷ)<m��;�{[��&x=��D=庹�6Ҽ��)<v�G;�#�:eL��s�=�P��#;pv��Iǈ<�+-=�%+�e�t=��=�HC=��O�g�<'p��-���O�ƻ[ޡ��Q�E�<�E=������<�V�{ B=Z@�<�VP=�[a=Y5w�D;=��<��(�
�D;�4�<P���f�=�*0=ҿ=O	��6`��#D=m�ټ�,d�ԭ�<6�;j�ջ���;��(=�)�=��0�#�̼.R�;՗<-��<�զ�1��:� 1���-=���;�S�;,�<*��<�(=�.<^���=�����<#@A=�֯�g�x�ޙмT�=��%� ��<XJ=�N�߆�;e��������)=wV=��3�mD�Ʌj���ּ��|��.%��#�-�񼺬#=
�˩q�����)=ln=&W�<Q>�¿���¼`�<�C�$��ī�����<��<��=���<j^D< 
=�]U=�i<=��X<ꫪ<F1�<�C�4�9:�<)��;ɩ�<FO�<?I���|ᠻY�<$�<��#��K�|=u�L<�	=;�x��Z =�C��]@�H ��7Y�v�;�]�;���<5�F�`�4=2p��Y�;��:yl�;�I=T0����=�<P;�K=�H==v=vmԼ��'=tQ =������)���u�m+�������8<��=�G~=���c����<����Nm���ȡ�!x���)=#�~�)}g������<x.�<�Y2=�u=l�E�*Zͻs�O���h=ԟY�e'+=�г�Vn�<V8'=Щ��N=�$=�=N���p�;9��uI����H=$�Y�
��_!�1x=�5�J_&=?�.�HԆ<
9=o�����<T�;�|W���<�ؼ��;�+<�M��=9�==��=���V��:հ���:��<R�>=��=���s�W��d=�􃻢+�<��ϼ�YF;�qؼ��u�@ �<c�=�'N<Z�H;��6=��u�S��<W�8<y*�;WYV<�er=����D=�E=�ك�*_=*/��v�^A�5<�]_=3Dx=�ȼV�3:?i�;ߣ+�����TQn<Iw�j�<�ɼ��B=��G=l�9����z+X=)�5=�8<+?�<���<��H�����3)�ފ�<���7Pb���d��%�R =k�<�.��Z=�x=��~�z=��Z&�N�<�����=�<��U<�����R=�4=!���Ψ����;2!�/J��D4��G�u�'^��8�x���Z���<��������2K�K."=�%R�a�S=�=-2�h�2�l�=�$2�����)�)�<l�"=���<�t4<^��<,U�<��<���<h�6�1E=-
�3� =0�������y��t����eżnTZ�#�6�(S9���4=�xw��UҼ�l��a�;-N=�ܓ;a�Y���ڼ�G�;h8=<���L-=�'��&���<OcF=�<�G1=�o�=aRa<	!�M, ���
��X<�"x=��<;��سʼS/?��R��!�=�-j�=��<sv�6U
< �#=>�p<=,�<�m˼�D]��<���;݊�3=Mw;�q�=ij ��(7�A�<�:=���
�<�I�v\�<<q1<EZ=ki<4|R<��׼��<��;��e=ǃۼ� T�ҥ�<��'=M<�2q`;�eG=Ƨ�<"��<퍼<�[L=q�%<�N<��4=���;��<�|G��^g<����Z=����1����/=�	=s:�v��<��J��4=�EJ��� ����=5<�="^S�C/<O���.\;=��:�W <t�;��=����E�h���,=}0μ��̻d�2=�<�<ui7=..j<3�#��<n���{H<B;��n;l@�<xe���e��;�E<#`3=���jQ=�Wռ[�=�^��� �?���k�<�0`=ӆ����><��='R�;���<\V=��"<���<
b<6Af=�0���T�o���N���ݎ<�僚���j�2<-�.��>��Ä;}���i���t�Z��<��q�q��zU�R�X����;=1E���";��=�G=� ��ng;���<v���K�<�s�<�P ��s�;=���Bފ=�Q���������-Ae���9=���;��B��n��p�=,���b�?���4qY�k����<_^�4�<�~ż� :<�I%��"��=�H=�:�qb�|&a;�J�<��= �.wV���=�C^^=��C;n� =�B\;��F��t)=�`�:���̻�<V[����D=���N��;�;|�V=��<�x���,����<�p�Sg���aw;�����R�Щ<EC�bo�<ox��"�<ݮ�B!��ƿ��6A�]ߢ�h{1���<��<����#����o�K<�m-=����$�m�r�z<W�)=��!=@l(;�=F1�<"�J���2�i��<.0�<��/�'BB=v�"<�@��p������>�=P��I���v3�;�Z�<���H�ͼ�m��gM���@<n弳�D��@�<�̼�zo<)�=�y5���l��\=q����ú���0=�Q[�y��<4K:�f�p��Uf="�Q=�|�<�F(��Z:&��<գ%<m�r��Ю<V��V�<mb�� \��	4�T�<���;��L��a?����#���E���w=�E=���刈��'=�T��$����ܑ�Pz�<���&k=B����=��~�,)�<6NI���d��<���<:x�aٱ�W�w�C{ɼ5��Tۻ<�@7��0%����� �<.r���v=��H=MfM=��Y�62N=T�&=�[�=F7�t�����7<�Z<�Rʼ��8���;���\�<�|w=G31�L�<�&H���O��Xż��|�o~�;wл�2��#� �d�f��f���U�Z�<�p*</½<[�;�`B�>�i=�,q<�S=���<�A��+sR<��T=���<S<=t"=c��<'+��L�4�����W=��i=�b޹��1��<;X���U�v�=��V��4g�x����)�R����h��71���0�ur���=��g=�����0���+��,=>�<��<�I=,�ּ��\<���:@��;��=�;'=�Gм\�<Wp�u�7�ܒ���h�窣��LE���R<:j�;G�����,=�i=<'/��A=�n1<�dq=�
����<�ca�'�o=�=��=�*K/<�D�<�κ�~}¼��P�hk��h=.h=�i��Hc��N% =�@G<5�K<��)=�PC=5�&=��<�T��g���.�<b�= W5=��d�9DG�;�|�ރ�;�^:=�S��=��=3&׼���	�;=�=�`K=gK=�7=���<l��l#q���k<^���޼"R=��(=I'��V�<������;��G��g><��=L_=�W�Α�yXM=�&=L<^^弥�3=�M���Z��(�<�DY�J�Q;0D�<��S����;�g=��*=���<�F�����˿�<��a��U�<b+=7�;�#�V<�갼�"=�<Al\<g@h����a_�Rk�<Tlo=Ў<ǆ�	���d�¼�Rʺ�@ӻ�ü�"�b���L����=�%*<�_'=�mL=y5=< ��;�H�(g�<�C9=�h�3��p	U<*<�<0}T�d~3��o�7� =�M��TU<ջۼ�+�`^�;6�$=�y=��'=H:�K��;�M=H���۾�L�A=�V=�rM���#�4��;��)=jt=(�l=�;1ǋ�Q�O��a���k<��Ѽ��;��f�0�Q�s��<�;x	�<2��	R��j<wͪ;��*=n\}<}v�<'p�8]
=�1�5)�w]%8s�I=��_�A<�_<A�<.���*j:=��N�Ʌ0;�����$�P�v=�X�|��;%�j��������+�b=�H���2F=ǵ0=p�׺PNh;ω��芼Ō"=ٱK�6�v����'r;t��)��&f����֘3=}���^b���V�u����@�bqӼ��;�b�A�h9�H}L<�DY=���n���V����N��q��ز���k���W<��{=�O�܀M=�B�<G���W�����9R���i:כx��O=c9��Ԕ<��c<=�<ǉ�f��;!�¼���@�;�cֻp�[�ｼ(5�٣�<�k<��Q�"6T=y��<�w�<��3�++5<[U,<�J�����А<b��<Ԝ2=-��<9R=3��<�]e=,�b=����@�;n�U��ˉ�1�<��s=s=�#=��<ؘ�b�	�����F��y`�������<B�ټ��!�=�=����-���P�<��;y�d���[=�q�<Ot;���v8=�H=E�˻B�<m�m�n�#H�<��=G	=��	=i$N����:��v=Ao�����<糈���7H�<��;/Z�<Y�=٩Ǽ(�;�h#�:0�;��(�&�]���;>n)=�x#=�B=@j���a�<��+	�/V=+>=�G>=�ߦ�>x�A�ֻ���.'=�O:
O0=O`;��<!L=�0��-��:]�2���q=�X��UT�[=:Z�<.Q���R���L=�;<=LA5=�8uĉ<Ǩ&��&�<��D=oS��Hg<VQ7=�9v;[��,6C=*��dg/=�,'=xXü�y:�� =fܶ�s8�<
:_� �=3�˼�v�= C�<<�8���<��=�ĺ<��<\閻��Y<�V��j�	��i�<�ꐼ�j*=��*\����<�b[<�Eo=�ғ<d�y=?��<ѿ�<��?=Qe�����;�?��W=Mc�7�#��}ټ�1���F<4�=dL�ΪC=7���e>�<��J=LI�<�\��5+<�6c�4��^�:=���<��A=�'h����m��<#�Z�R�9^!ü�)3��/�<2=��o=�L5�E2���7G<��=�PN=DH� �=�S��¸<��<��'<䥻;j�=M&�$T���K=�׻�L��	> <�9�sx��ǔ<.�4��\E���R=Ж�<�/������Hf�V��<��<�\#������^=�����`�;�L~�$�j;jDO=;?=D��/m�=$(��W��?¼�a=�m�<-N/=ў��
=���<�k=i0\<��&�#V�<�p����;�<J�U=NW�6��J����<�큽��弡�]=n�Q���p��M��@��<l�W���U��d��. P��p��<���<�d=<׼s� �v<<__�<��a���8<��&�F(=c�ɼN��9���g�'=���3B��/9�O90���u<^?�<�r/�S�}:B�+=ӕ$��N�/�W=��<7[K=�;U�y�q=�f�c�u��wy<LRR;pi=ɨC=�yҼ^9�Y3=�I=l�!�O	ؼ����M缒	�W=�Ͱ<�=lz���� =�g<�C,��ϧ<��Z����_�/=�;^=��;\�ǻ߳9*�¼��:B=#3H�s��9�V�M�<q���d�Ie�<�Mh=�=7ۻ=,�l<�|;=Sq=�Q5�Z/x�y�<U�P���(<��T�-R/<�*��:� �M�=��\��`=��4�ܿ
=�H(���<*�;�4�<�=}�A�s��<��ʻ'f���=^>��;�(4����=���<9�=��ۼ���]U��=��_�
<8�U��^=1�l<}�ϼ3k�V�/�"<R�zN=�WU�v�f��-5=^�;�ۼ�����(��ܸ��r���<\/�;_�"=����7G=Tby�l��g��F˼d�\<��<ۛZ��0�<��d=��j=F
��o�<��%�$�.=��<�A�5�&=�~H��'��WC=�"�<��s��_��3���E�<9a~;��M;j��<��k�(<�=Dp
�S�ϼ&z�9Hv�G�=�C=�~%<f��KbP<��,��:=c%�������܇<��;;��=b��\�1�YJ/���><�es=�{?��5=��_={TB=�~=�u�<��1�_�<3�H���=XZ�<��<��M�9K=�);�(�-=���;��1�])��#Z���$=Ed/�q�H�>=%'�rl�D�9�؂<��Q=���<]�=3�<��k=��k=Yj~=����a�}z�Z[�<*�&<�O�<��)�9=D�<��<�"Q�<;��;���<�Ʌ��]��}e=�:�<�H��nǼ-af=���;B!`7�y{�=BҼ�$Y=2�_�
W�< N�
B ��t1=Y����<��-�L=��H���I=B�?:D3Ϲ��<>�<�*�kEP��A=�<P������9�v������;� �����:�¼!n����:��)H^;���;�`ؼ��=8�!=̨D=�9=؊���1:ۜI���(=0v6��o����L�ļl��<����ġ<!t'=��<�=��D=�@v=���<|-�<H}��t�!=HF̼U�J������C=d%������%��	���7��ŸD��""=J>��ߝ�8)l��ޣ:�}$�N���ռ�`�f	=&�ټ�F"�0�*<
�λ�Z;�j�@�<0�9|,i9�6�{�x=u�^=`�C=Ok��� ����� ��iA;�A?=�~�� �d�?d��W|D=Th_='Z��������M��;	u=�!\�L��<N��<_�A=��u=� =�ZJ=�C^��bI<N=R���=�<���2<G�=蘦�i��)+���;;o�����&��<��=KM8=�q��c����#�;C�=�5ۻn�2���K=,*�<wH=E�}=��<�m�=W]=��<���}|4�d.=�%m=k;��O=��H;7`�<<ؼ�|�#��;�8�<�N�-���#<\I��<�(��C=�@<�T�j~=g&ۼ��Ԛ�<�r��mK����<��T�G��*�E�
v���g��@�MZV=5�'=ĖT=Ω�<��м�g�<qʼQFz<"y�<d��<�n=�X��lۻ�{�<(v�:�u6��f�<@|�<q	%<���<ݍ<b=��6�><���<�{<���<�����\��/=��<��=G�d=5;+�O�|�w�(�u�<8�<��<��M=A�<R��� �=�8/<<�
=���<Ӽ<�=�c�8 ��)q��:!;�[컉�
�l�L�^��� =���<hz4=Q<G�+��K+=a��<�[�;�"=㹦�G�;�C=q�=� B�Gk�=nҀ�Ƅ.=m��;���&2�u\	<�x=2�d=�;=���<z3=}s>�W����-�'H���t*��8�ޝ߼�W&���i�� �<�b�{g��p��FC=x)j=;bF�^�p<���<���<'�����vO�0�'��=�>h<���9,�H<q
�<
s<��0��U�;�q(��Ry�_pA<������N��;I�e��A(�����7R;=oAt<���<�
���f2=��=��<�K�<ru=Qּ��<�>��=L���![��C�=�d�:�e�<���<ɴb��*�=�r��8�2f9�y���\��x�<u	8=�K�;\\3=��b=G߽�������B��K�:���b��<_+<D��<H λ�G�<hj���<܃3=��H�N�o=V���=lq\�?L�98b�;$7y=h=�#E��&�DL�BE;=la<b���)6<�����7;�I<�䙻NϜ����<Җ�_h,���=���v��8��b��6���ό��p�<x^=r��<�?��U��j��;l1$=��\��=���;7<��w<U��NN9<��r<�g9���;��= 昼<aE=y���5��&n=�G��s��/A�=jϻJ��<܎�<��(�ޥ�� 	���6=.��=$�o���|<Z�ټ�#��|a���<��o=��t���4=ju�<�i:"^"=�uz=�w��o�:�n�rw��NüUI �ɼ��=�ۡ��b/=5��;������_����ng'=o5�<�x0���0���;�I�:�U��+t����a���y�3�=B��.�d=��.=]Ie=`"S<�L@=1��K=����<�h�<�%����)�ap�<M�3<�e6<�]=��<B#s=�Y=���<"<�GJ�������<�O<0Q/��N��=��>�<��:��%=ə�|���>;h��<?8�<�>=�-�Q�q��m�1[)=��S�L �<WG����ur���C=�C�<�����W=G�4���*=�C=1@{����<nBX�ݚ��m��<�r��G��<+M��� <��7=¦.��Pn<��n���;ˮ+��#; dǼ��Q���=@�}��;�<��<�*o�d`^�i0=>e���:�c}<�����<���"<@��bu��#p;��ڹ7=�e5=��ݼ��)���Z���n<`Bp=��p;��'<���k�����]GJ<`Ad<��=��g=�F�<�G=u�<~:=�[=��<�B|��)=qlc=:��<s��<��Q����<�K��Ἐ<��v=Bzf=?�<���6;��<�����m�<	=Ŝ��X<*����;N逽M�<7�:�U=�ھ���<$5=���<��<�OW��́����<�L;=��7�<�2"�}��<�=��Y=Y<3=V[,=^1����	��� ��xz<\5���:�<9E�=�=bT<�
F�<�ͼ�̨<�x�]楼�$k<��ļH0��=��`�Ӛ <V�=n�<N�N�9k���ub�I+��.b<z.=`�<�;(�PJ<��2����T$=�⩼I�;-M�;r!O��k=.ጼ#�?���7=��=G|�<�u=85��5�W6;�O=�C�ɻ�4�l�f�X��;�U	=M�9=}5s�0�vU6�����!=2|���1�ͭ�<?H��"���U=�l�t#6���)=8z�<��=
YN�(�<&)8��9�;�/*�pY=�ߍ==;Z=m"=�*=�OǼ�ݚ�t%=��<���<�=$�w;-T0����$H;	�d��VZ�WC�9�r�VM�<?���1i�����t��8=N3==����;=��m�<�������;�[�<�Z:P�(=�|�<3��<b����f\��h��Q1��k*d��1�p�;<�:�<�Z8=��=T�G����<;��(< <�-�6�k�===p&��q1��~��2X<��<Nln���i1����<�Ҧ<�m=Kt<=�!;Aw���t��5�S[���7��J�������*�86N=@��	�*�=[��$�<�t<Cu#��^���1~��u<Gl�;���<�}�<e��;�/�<����K3��me=O�t�7�
=�I=.��<5�S<���;�;S�O���/��� ��}|<׿�;�=��j=i��?�M�7������/ʉ�!V��
*�N"T=�<@�$=�-=R�>�?_���m��a=�:,�Y�\���=x����=�M/=������i;=�g��33���Ӽv|w�4���Ja���<���s�o= �/�8(Y=�R�;��<��t�7�S=�B�<��A=�\f=Tz�l?��.�9�6�>d%���p=�c��'	�����y����fGJ�3i`;xu�<�rQ=ob�<!p=��\<���AļڋC���^<C�ռ�GҼ��!=�5S= `$=ӱv��YŻb����hD=v��n?<Uٗ�F�*�t�<��W������y�?"=0.�<w�=
iQ=��R<޽�	�2�L��<�����Y���=*��<��<�����0�$S;�[�=�����< s���T=�I�:�h�r�<۩��ِ�<:)=��M�S��;-�<�,�<�Go�ڄ<�ꙺ�]=���;�d<�Q<i5��Qy=�*��[U�
7� ����<�8=�=;�	=��
�E��*�0�=\�A����<��=����e�9=�@g=��N=�\K=�j�<���<�р��K�`=�p�<�	j� �
�؂c�����_q���=ra$='�1=4�5��F�gf=/��<���,����M���8=]�Q�:��<YE=jU=P=���X'C���{=���;H�V�v<z)=���<EC=��
<���<> T��|=�g����Ǻ��J=�M=g�;��=aG=�Sܺ��<��P=�ְ;�]�;�Bϼ�x�
|��i�NqX=��;DW<�w[<��k=��C;ƇI��;3=
��<��<g7 ==>�<��=�T����<��7=��B=���<��<0Xc=�\���l�Z,=\��<{�/�Z��"HS=n�E�������ۼ���<H�M��� �L�j�
��2T�J�F=��꼖�o�d���R}�Ԏ0<�bS=-�;}
,=���<�<B�s=P R�y	(�.��Tc���;򄔼�9�<��;<�5�< =ؒ=B�c;T��Q��<\��}�>=�4M�WD2=�.��LF�������e=NX�<���ꂼ�~�<_^�FP���]d<����b�U�,�<V���D��;�=����W�՗ټ�����<��ټ'gm��[J=�Mo�m��<򼀻���:���]�Z���<P@��ss=� f=��<�D��s�r=A�= �<=��;�vh=��<=K�2 �L�4�V �=����_���Mh=�Y�K߼$a�<l��3V�κ����\�;�� �0�<�a�FZ=�ّ<���E�$�U��<�	=X!�;�2s;�Y�	���c��U����"=FC=�W�,=��<�[߼�6����jћ�y�A=8V�<
�m���d<��t�<M��<HsB=�W;���A������S���R�r]<�����:;��g���ۃ�_.=\
���X�F]|���׻����{dM=5BB�ae��bN���!�r,#=)X=���;at�=VA=�l�<������6	=jA�=���/Ẻݺ��=��/�oF���(=�?���M= ��;��=�<?E1=���~�;��碕;j��;�l�<��9=�=�=��ռR�=���L�׼�e���<��P�;��+�rX��ap�)n=��A�ʬ�<��r���=m��k͡:���<]���:��<䎺�x�<ҿq=C���c��ai����<���<���<�e=iC�w��:l�	�+F$�d���NA=JY�=	��<��<��^�U.�<o݆<��l���<���z�%e�<X5S<Fr[����<Ў�<o���EH�$I�<
��7<����.(�T1�=�G=Y4e�̸A�� =_�7��G�B;p<��<
��;�٨<E\�[��Iu=t�i=;�=��-=�=����Y���I<�+R�݌�;]B�q��<o������X���i��7=�O���� <�M�<�Vm=��=�.���.<�㻬<K<��HpA�#un���=�&:��<���=�$�=F%�W�}=���=�:��#�b:=C,�;Ȇ#=�4=�RR�����Wu�z�r<��񼽹�<�N<�<�������-U=Q�R��¼�k.�x��/[��C������Z��<��<�C=�V<�A�<A ��){K=^>*�|7�2�=��b�z�=�q�;������<�=8t�<������弴�/=���<5{B=4ht;6�'�Bo�<�d��w�[�<[�'=���~Ɓ=4��3��ŧu��o^���V��z�<� �i�L=f�:�r�w+�<oh~=(�=��̼N�G�v�j<�[_�.�t=gy�L�f�=�5=���<��<l�g�ͨ������GA�m
�޷/�Stz�~&�;��<��%<?f�<R�=|"?���˼�@���A��U=��e<:=�6v�O�:;b��;�;<�7<F�Y�)�0�W�C��Ѽ�N��E�n������<a�<f��P8��d�ּ�A�<��;���<>��ca=��S=��Q#]�k~�<&TF������+=�������"�9�A=�.<Nj<��==�==k�<�h=T����`F�i��<UL9��3�<
\�����`=z�߼�g��zq��=����g=��;�($==���X��<y˼�Uͼ��,�cn���t=I�W��=�Aa�T_=��'=���=	D=��8=,_d�"�軁KA<�9�~�J=F���A� X���1g<Hm���
;��=G[<�b=Bei=��=���h	|�hn=h��i�߻�;==&�=O#r=�d4=n�y������׼�]�����C�;m�����"<��F=P"�<h<�!�<�F��6;<�
�����Xs;ȼ<�����,;�%*��/=w>��AO��s&=:"�=�^=�=V�s� A�;s�<�i �����O����H�=oN�'8��`<����M
=���B&���^=P�<O�=`�*���<��=;x/!��)�(m�<N{=W�׼aF=�Q6��
U=��7��h�;#rS=��=ۆ�<�<�O޻G�<C�]��<ἰ0Ⱥ��=��;aY�ʣ\<_
'=���'y2=�k�&��[j���10=�2;�n�N�q�U;S=Y3����;�-�7%�����=���:�>=�8=��<�F"����i�:���u+�(�8���N��[=n�Y�9�+�A�<UcK���G�k���?!�-�A=��<�#�;Hu���C=P�`��/�5�<�!�<e�=n�<�z<`x������Y<R���N�� G�<l�T=3לּ�je���8=�.E���=���;�'�<�~߼�`�<�X7����v��;G=?*̼HTS�cj�<H��<�����߻`����'�<"}����<�t=ՓR=`2u:/껊�=���9��8^s={��<�Pb�bYg��BW�k����ϼU�-<��<ly��a�;�(�������:C�+u=��;N�<d �����;�[={מ�cmJ=)*
��Ť< ^d<�%�L�,=���;�;��z8���!�s����L=�J@=����H����<��<�\����i=$�;�=����=�P���L�<�&2=��,=��;D�ϼ�׭�G�:�h==�<�����6�<�.�<~����d�����]2=6�kJ�=JQ�N� =y�P���c=6�=�<!�p��<D��;}�;�I�<W�T<ޤ<?��<��p��7��x�:�)=>Y=�ѻ���-�
=t�]�:�=��ڼWU��*��>�;k:�; �(���W=W)�<7Fi=YQi��um<�	�<��-=��;�*F�D�@���<�[b���_=|:�<��'��i>=��Y=��<#�ֻՖD����<���\�>=<�4��<�4��Ꝉ�g
�<�Z9xM<��ؼ3! =x@�^6��=��l�==��ü�������=�����<yz�v����3<�������s��E#)�C;)=�i�#������<��<��)��k<���xݒ<��)=B7�<��4���S=ڣ߼/#-=P�><b�-���7<��仌������`�◹���<&D==γ�ۇp�)�k�4�M��T�;*�?;�QP��=�<����z=`X�;���<�P(�?w�;)f�<��V=�'��A�j���<�r�߼�=jڼ��K��=��Q��W7<�9�<�T��;��	�@=;���=��<�}�<���;{ �z����]<|4g=`�P<^PJ�i9<u��<�l��R�.�=�'=�`I�1I�;��0�#�o��)�=�d�o�	���)='ꍼ�(K=	�H������/=~���	=���<T�=R�=/G�=e#�;�W�<�O/=�
�<�V2=�Zܻ���<�w����
�=��=�?`<�Iܼ�^={9d�P?�<+D�ra��ûڤ�<Z����p=��<�¼�$:K��;��>=�I�ޓ�=�6�׻IH=4��<T�5<�cq��X<�荼R$����G=>j�\O=9�a<5u�=&YZ�����s�=���;o;�<z$;��H�<�>׼&�,=n���h���)==�H=Eo1��~@=�(?='<��<#�c<�@e<�p�;��J<�Ո�<�7<�R�6('=��u��<��I=�7=Qz�<:h<�N�<�m&�?��L��a=F�&=�?�1ڸ<����Iڼ̇��Y�&�JF���=��=���T�K��<n�)��y���QC=&.=;z?�jR<�:;�_��P����<*�<�*;f-���ׅ=F\���ͼ7�x="38<��I�f.M=90�3�.=6m=v�T��"=W�q=��1��#=�=Z��;��Լ	h�<�s7<d�;e��T��;��j=�\f�}A&<�R;Z6<^��<"�<��
;��	���(��׈<�_�=-k�<��]�aFf���~�D�6;.0Y�'�ü��c=�񑼿���=�7����<��S=H�><+Y=���;�:=��L<!��<�%�<�<�v}�ϛ1�ք���m=�&�5��<�h�����ɓ���a�F�=�D-<��*$U��<&n�͋<��6=%�ؼ�"���RO=jL;�T�/�}���Q�;ϗe�ɵ����׼ �=�T�9<��+�B&9��rY�~�u=�0��_k�|a��d�:��b=�<�=��Q<5�Z=m���k@x=� �8��;�\a=Jh=�`�<ʦ��`�����y����|#<�9=�D=���<�����<ż=ӹ<�H=Yk>=wd�<�<˺�'��mռ���<6�!��W�� �D�6=��&�F��<��;��={E����S�c���f;x�r���%=��w��?�<4��<���e7=��@�H�P��<
盼�'j�Y1��:���=� �r��=�
P�<z�g<p�<�▼�C���>�2�;�;=xg��t��<�ۻjip���p��o=�-}=Q߮;$��<X�꼖�ż��l=����%/�<�1<�S=C����<�&�A<#:�j������<�c�<ш9=��=-�B�.�')5=�����^=����弭	F�Dp��^<�O�<o�E=��1=,���r<=ȕ����=ƽT�X*�<�M=��ڻ\�X��k����8=�=�hI��
��Vs�<���_J<� ��%M=�Hż�I�C�<F�w'��;4���cм����M�":U��-�Q�P�F��5���6=oC�<ދ4���o<T��<���<|�O�0�H<�Ȯ�W �!xo=�/�<T�=2`���[:=���<WRv�0�F<��;���r%�
�N��?R=��W����~HD�K�D<d=�<��͸U����@<$�:���<�wn=��A=J<ȋ�<�P�<9(/��"A=�ݼ�k���R��ٚüi֧�������;Y���w�W���Y=bV=�V�;O�����$<u�g���K��~�;Ld�bDR=�"Z=܆��H�J��4=ݥֻA<G�Ȗ/=ܐ-��O��n�F=nn�<؄"=s��<^�U�i��<��>=_��B���q���
74���yPh=��H�Zm=��%;�*����6�L�:�~<��޼��&=?�<���"�c=+�j��M<=��D�6T�;#w=v�ﻃ8�*9=_��{޼ueټ7�0=2�=�\ټ6�=E���м�e3=*1����;��<[-<< ���=�6=%�R=چ�<sog<��W�W֜<�6d=W�&���:膼a9�:��!<�z<9�|<� <��9��=p<�O=���<ﴺ<�� =�b�<'^+�E��9�b��L>�.�4�|�<���#r=�=�<�����<M�w�p���~.<��.�ՙ�<�A�+��pzy=�(�<mg��M���=&��ʖ1���1=�9=D��<T�ּx��{^�
�9�-<�;�Q?���*d�<l����7�dqW=�ټb~F�&����������>���|=�%=�`P���9�?���=�<��ƻ*��>�9�XB���$=���<�Y8<=���s�=�����w=��K=�N=�E=��g�H|C=��=�s�^�^As<�����<t
�.��z�	�.��&�=��W;a��<MA=/�L=Q#�d+J=�㩼q�Z:Q�������R5D<y�f�:�#���2� ��< �[�,C�;�s=�����,�,�1��켝ph�H+�<
Q=���<����:2��<��v<�*�<�T<��m;�)=G�ɼ��-��n�aFQ<��޼���<�)�<3�%�K�=����u�=&=���Y��鰀=<J��G��;�V���*�8=�`��=P>����@=(�=�;=�52�(��l�<��f���=�A=�h�;������;<K�p�E��r�<�sû��;�<��s��US��p =��N�/�Q=������ �0ܺ��=1�����<�(�<P���n<� <=X�A=�f=j^�<.i=�	�S�-=��߼��!��컰F�U9H=�،���r��t;���I�ܱݼ�6Z�P��́<�m���w2='J��g����r<�D���Q=�q=:�o����&0b=������=
�`�z��#簼w�X���
=y�,=2��<@�>�%��l��T=���I.�<P	=ǫ�;�=ڼg�f<�-&=�=�;@�7-���<ƈ<��Q=ު|=���	¼~{3<ylb=a��<���%U7<è.=��?��|Q�((��e��b z��;�<9�n<�ԻU#�<>+��B�a��<{X���> ����=�d�:1�@�}��w����o+=V�Լ:|-;;�<��
=� ���7��t8�	Ғ��AH��^滼4�?ER=1B=�P�����aVA��[9��/=�Io=O*R�r��:HL��0=�Fs�7z�<2�*=뿨<k��<S@=c[=ڥ>������#�񓺼?�<�4=.�)��)�[��<�k�o�
�c�%=�g��>�<����R><W�<�c�9��<�λ���uC��]VW=�R=״E��Ӽ��~��<=
L=�`$<bb���"�<l��D#<��Y�L =VX��}�<$kx=�c
=HhL��2���%�擮:}tI��GY�������<<�����;�p�L�=ދ���7�a>Z<���o=h�(=ZTP�;�F��;5nN������T���v<�v��Y}<��;L.=�a=7F=����<4�<���<�&4�~>=?�<jW1=�d��85=U&g;)!?=@=U�,=�9�;)�G��6��:	���<�=��"�;=����z����;�� <Bм�*��$�<+Ħ��?x���=<3d;g�C�Mi�-�мt�Z�s�[=}h�R�$���ʶm�)��]����](��?%�<��I�-�ҼO�<D�R=��<��˻�4�<��2=��<�*�J� �a=(:V=Al=4�<�����R=y&;=���<s�&=-K=}^<v�&=!B��70�+�d=\]=}M=:�<����<�t<҃d��w���O��CfԼ|�b����o=� ,=40H��2=�-лA�E=�&=����^=�hT=�l(=��<H�=��P=��<�>���;��<E��3[P�J+ݼzu =X��8�=��t;u�[=�� =G�Y� j��M����E�0{�.�<���<T�|�b�)=O�<$$=(>ּ�C�<ǪH;{QH�4�a�;H=_����H���<&�=�>=�gB�{��H�	�=`Z�=�@=N��;�j�;�@���2�L�I�kx=��j=V,;��<$a��9r=\�<BČ<��3��{=��=֠�s��<�O�rc<�<�<|�+�1�<�&=i�s=��=p�-��<RS9�c =<@T���@���M�K]��u�?ʽ�!��<{�m�I�'=���<q?J�X,��ܼ"W��Sg=������;1D{���_0r=�U���?P�@�[�?8�b���^b<�;=��o=�F���΁��������;/�<�X�I�"=�1�-���B=0kJ=�ü1��P<�O�-=��>�k')�&(�y�n�$�e������T��?n�c�=�F=ְȺ�/ֺ:������l=De��c��=-��x��*�<�,=��*�=�c��s(��R��p|�>�輀�p=�$�����.�<@\��4��;{��</��<2S��@�	� ��<����+�a�5=$x=�\����K=�2��e.=�j���<�$�A�n=��?���W<��`���j�.nɼ^�=��U�<�~����Y���=�I=�zT=�
=3��<�J;_j�<��;�@�<����B3=���<��<��<��i=Gѻ��H=�H��u`=;]=���V��m�=Ӑ�?ܻ��.=�)#���Z��
��w ��O=q�鼨v�;�1��{M��0��������;=3c|��,8�1��ˇ�6Ժ�S����<de�<K�ּٕ7� �=04�����<I�s�j6;��O<��$=�hQ� ��㟼w.;��-��CX�����&;<A,H���B=����#2<-ӻ@����=����ij���(�AGN<���<K��;�@c=�w=���;�0�A�=���p=�����3押��:-Z=��X=s-�4�@��?=#Ɛ<x�?���=�W=(;��Z=�_�;Y��<6����W�<��E�6��C�I=���<�K�[ =�]���ʼ�dѼ,@I��p���J���<�,/��v�����H0��晼�[������&9�*�<M4�=M��;L7»[Z�;��=��ڼ?�=�=縹���<�����ء�c�<�^��s���B�<vH�<E� ��g��Z=�N�03�<ě;�ϯ;�����=��]=,��<�2h�e�����=z�3w=T�=_�Լo91��dn�~��<�>�;�m?=��&=�z_<Ťʼ���qD��N�<u�h��=ym1=�����=(�=�E�<a b���*;>j=vpռ�ừ�<������7�.��<�p�;e�u;��`<kF=]�}�l�o������}[�o��� *�iQӻo%ټJ�<��껺�<Zd=t8���C��&��5���?�;x�#<\=7��<;����C�<羛<�Ļ��F�!�����<{u<*V�:dd��w��+�<˝s=\%1=�v6�T�r��iL��W<՘�<����h<W��P�?�g��<�	.����Z��<�V"�:@�<c�&=g]m�4����z;���=Sc<�b"=���:=u�Q&8�AZ���P8�05��S;plD<8�V���:;�x������@�]b��h����B=jI(����<?X�<�R���2��/��D}k�ߡ�4<�a1�<Z�(�(YY��R�*�K�����샼_�n��}μJ�,�rZ���~�<Se< �g���"�YF<E��x�r=o��<�����H��Ǽ9q6[=�Q"<J]b���\<IE{=6	��A@=g��;yS�?�(���9�
����g��)�.{p=��x���Q���i<�f=�t������!a���i�F�i==.׼^:M=|ɛ��D�ŋ��e>�<[2��k�޼�co<�Y.=#KM�gE)={�=��ڼ#���* =Sk<��漫�(���9�ld�X�vN�����伩j��a���YP�$BG=V��m)���泻�0�*uC=�|<F�>��xU;��<��[�:)�N��6=,m����ܼa�<g��< �d�
=[I��~n%=�>$=�&��q<��I��:��4=ٽ<$��w <{R<�� �]D=�ܓ;���둓�!;��	��Ơ;p?==p�����<�g�<��E=u`�^/�;R�o���J�r��#v.�3�Vϼ�"��<�<��Y�Bsr=�>j���Y:y2�<�@���j�����<&�<�@�I�,�@�==�<Y��pC=vYQ��uh=�F ;����p֥���L=��K��v����)=�	n<����tT�+n��~")�B��<��A=~wʻ4�<��;qF="K=|?q=�����[��ʈ;-��:��<�B��܋;��c�N�=�a=;�F�[=�Sd�SU�;��M��`��[�UPZ��;�<l`��N=��)<'�$<#���ϙ#=�4Ӽ�?<]*�<��I�26='�<��I=�[�����n9�;�Q�<���<3H=��M�ԧ�t��	�=�׆<;X�<4\q=�KX=Dy�<ǅE=��8���n<T�=jn"=�v�<-�R��=xlZ=��G=Qč�p~�<�޼��=�p=�?i=��;�1��D=w;)�!G[�<s�<[�<^��&W�<�C���l�<�˼<K�!=�O �ϞM����<M�9�,�/9��`<�ɼ��==��kL&�j,=]��<�����Լ�Pm���<~(�;�μ<��;��,���:��9��8��*@<��=�p1��rX���==ӹM��/@��{<����}<i�(<qh=Ȃ;=̩¼`ú<hZz<�,h;�==��=���%��uؼ�������<Hk�<�/=��)=з=?t7=��{�1�����-=+���G<�͙�Xѿ���&��=�ϼ��;�I���[=�@L<�r<���s�<���a>�Q&�<9�<=ڥ��/�����<�޵<�3�<G?T<����	=w���,�7��A �+q=�2�<�&���=��2�0�p�N��<����<��d=�5ݼ_b�ͤ�����<NU0= �Ǻ0��J7<@�<e%
���H=�� =N�������*;�zt�YL�'A�<�9��t7="+>�*�5��������=��;^�L��J=mF�<i��W��!$��LL� �=f@=���<�f<����<ծ<)q$��t�=�)1=�*=���<닼������A=��X��2����<�<��I�*;O�Z�"P���s�� E��}κm��='M=qr=�eV=\m����':��H����#&=9o��
$�s��/F��s��<M!�:�D<�Y=+�̼�O���y=@>�$~b=-��)f��g4������p���p=��<;`痼#���RԼR�=ۃ=|!�}ZS<۽Z=j�/�܈�=��B����3=m�_�<�<���j;/�C�.TU��0J=T��<�ȭ���)=(�*�t�0��8];���;�ѻ��*]<��2=�P �8M�<킐=XY�<˼= lh=�@T=h�%�֔=l@��"�<?�&=cW������(�D=��t�{�<��I��Y]���8�V�4=��:�΁��?=A�8=�3��氼�+[�Ћ<S,��uaR���`=�N�<\K�:���
 0=Ԕ	��x<ٟ���X���of=���eP�<$�"=��ϼaM�<�0�<���9�g=����a��O%=ǳ��),������1=�<�Z�<9|�'���0=�=*k���<�~�v�IU_�M{�<. ���<�--�I�<|9��"5�6�[��M�<�3ͻ��<ǯ��W�����q�h=p��<�<3;�8������:T���`3=�WC=cU���y<�S�<؎T�{���֩��\=(`)�@y4=��n�m]�nð��@�=M��>)��諄���~<�u��f<3S����<=-����==Ȃ��\�<Ƌ8=��<t�Z����;ź��aG3��������;yA��×�HƊ<aY��Zd|��u�<�X�z�X�0�^��A=$�A=v��-=n��;������0����<�X=%U�i��;޼ n��V�==��<���<5><���<��E<fS%��z����=����̼��_;�a=�RZ=�?9=g錼b��<7�����m�Ԇ���B=�1�;��¼wx�2���ZB�V����]=��A=�WZ=>��;0�;�d����a���R*�<UT%��g�<��=�J�<���b�<OH¼�o-<��=�W='�1=�]�<��?=� ����*�ty7�S�*�Rs�:<]<�� �t�4=�\�8������<T]�<�>�<��;����H�����=��q=�/�;�Fs��S=��9n�;U=�#:�G�\�F<��/��٠��Q=s�G�6k�B8伝�='8	��;�l����:a�3=�ߖ���U=�4S=��==W!8<-C=$���3=�)	�s��$C��N��J'p�����1�b=`����>
�p�=�@�<�� �=��7��3=G��3F��8=�.<<�<�^=�)L<��<R�׼�Z��� �b}&<�(�;qL@=��7�'d�<͑^90p���T=��w&��?�T=�\�<s-i<ݼ=�&=��M=��`;�ĥ;v�޼�Ǽ�+=���>=!�)����<�U��d��?��\=�j?=�<,<��-�J��
�P�f�����Am���_y<������9�����<z74��Ī�;���*�:��p�ɻ  p�h�2=RT=d�<P�t<��\�����J�[#.=����� h=z���q=
}D�H��<�.:�ZW=wQ1=�7J=�	"��y<��#=W	U�G�4�1�7�yB
=S�f<�"f=�:<���<���U�=� r�ڻ�=f�N����&Ļ>:�8����:�弸�f��]Y����<�����<�"<��n�-����<J\�<�zO=
����.��%^�ҩ<��I=y��qᅼB�X��'=yb�=�@e=?ƃ<�
����<i�9�k?=�U��E0����,�@;�|P�L�]=r=/����	 �DN�"��<�U=<6,=�!: %��5=�p==0�;o�K���Y<#8��ύ���)P��''=���<�0=<֕<�D=h�7�#��<�6=�v�U�S=��:��f��n�<�|�;^	^��-����;�)ɷ�P�D����x<�4U= ��mfW=e�$=TI��R�<L�8<a����;��T��8��y�<��e�]���M���"#=�n �蝾��-<�����ܼ���<�ּ�k
=��5=vDU�Tn8<�-0= [4��3=�݂�oP�=я<I��B4K=�￼<<����۾<e\E=�N���Fͼ�Ì�A�_��jI���=q��; r�Ǖ��	���=~�=����<[q"=�����X���M<4ڥ��¼$S=0P�<f ���*�=�i9��K=~O=��B���V�tLJ���U�ZK����e�&�|;�r�<
�<}�� �7=��Z=Z�����{�1ԼM�=$��;ʌ%��1=���<gY޼i�<�[5�����҇"<]#o��i�l��<W�:<�ͅ;�>=�4���$<%)0��N=�~-=DF�du*��+��$=��_��V�<t�2�=p U=8��<��_�s����M=zs�<��=�rZ�d��<}���):�����깻�D��S}<@l�=˘�<�,*���/=`7#��"R=������<�ȏ:E%=��׼N%=8_O����<oC�<�ϟ:j��;�����C<2h?�ַ��^=�𻕭�<�i�$嬼��8;�	6<C�@��5�{1�<DЏ<5��fqӼ<�
=�A �n嵼Sk\=�᫼���Sޟ��
=/U=��?�6�W�]��_ ?��Ku��������Q���`<\��A���<b<i���E8=L;=�Z8=���־�=�N	��=�)/=P�=�Z<��=ɧo�*��;6"m=���j��h�n��AI���<5޿�E�9;ѻ]:I��NP=�PV����<(���`�����Fe=��<|
,=7C<���X2#��j/=N��<�j�<$�= ��Aɬ���!�<�E=��μ;a>=�ʐ�hB>=^���"�0=�ZX�_i���;J;�<ho�< *U<�ɘ<,��;�sd���<��E���<�k<fO�ONd��(=�Bg=l_)=��l=�3<4(=�<?�l{Q<�J=L���+�_=,H�<��j<���8u��=-쭻R�%�ί-=٢<J�==cf�G�\<R"��EP=O8E=�&o:�DH� �&=q' ��G��;��J�����:�Vz<��nQ�<����]4�C=�.=���7PX;_�t=��gS��B<�P��d(=���<Xޯ<�=:�w�,�:}�<4=�w!=5AĻo�a=m�˼]��<�w��Wp�ܒ��=�Q�<��ټk�I�ǟS= y=�����	��;��@D���e=Hy�<�{�<fW޼��C�1��<��j=&⌺�^s���;���;aY�<r'㼱<�6/=�1F��߼��!�A��<FM=1S����޼�q-=BSu:9�(���\=k�)=:>`�J�@=�PX<��y<K7��8P<��	��9G�1�l=�-0�����~���� �� �;͢o=��=���<q6�<�=+9�<�m<;���<���<bq�<��c=��;b������;�!N������;Q���]��<�E=����+�=�4*=q�?=�!�:�ż0�B������ <yM�?�(���{�=b�K=�b4=g�*��h=����Ż��4���A=���[��;�M=&�E=��V�N=?��<�ւ<�����;k�;|܍�Y��l9�^~����M����s��=�"����<D���7(	<ou�$y��ͪ;}�/��P=����M�<�S<�"��\��W=�z�<�t���}>�~��8=1=L-|�.h�b�$=�5�|o ��E<�6���w�fv��EM=Ǟ�n,$=��w��Aۼ�6���P"��ۆ<�[=��i���Y=X��<�ǉ���<�3�<<.*=��k�P���k�|�� ���=�沼C?���6=2u\=�v@=��<���H=������<F{-=�;\<��+=><�7�R�=��4=F��<dh	�N�����<�����P=y�'�R��<. 2=ޥ&�ac<(�G�"B�<6H�  :��c]=�ӭ;�"=�8	<������%�(z=��<)�E��я�NH����;��;=���
���2=)�L;�JX���<�iA��H<�o��ؙ�:��=x�=a=E��J��<ǁi=9��:Aު<��"<�3�<�]���S�����퐼a�_�B�����M��J=�<v:�g�t]���Q=��W9=�y�%�ż����ת�.\�<�������W,`�������8�4Pg=ӥ=���M�׼p˼5�<6^I����<���4;=��;�=��=����g=�=c�N=0%=��d�B<Xca=	Z
=|kZ�M�?< �é�<�u�<�YM=��S=/ex=F��<��d=����Х;�%l���r`�����C2=�c��@�A=�=�]7�L�T���5= @t�A���|x=_&��ݤ�dE<&h��N�ռ@���"R�������h�<j�<�>;��(=��c=z�;�����:=�G�<�Q�<D�0���m=�����\�jvp��m?=j
�����G�X=h�8��<l=N�x���=�{�<�\��;0��=
e�0�&���;�H0=b'�;p=r=kCV=��ż�M=L��_q����q���pOL��2C=^�%=6�<1�8��R =V�pY����l�I<"v�=�cp=�S�X�T�)�d=�14�b�ax=��<3�8;��y=h=�MT��3Z��$G�O#
���<62-=�P��:�84 ���R=��=�;�W�<@��<N��< ��U����%���=�[�2�
e<q�J�+̩�۵T���i<%G�<�*�<��-*�<��/=�����AǺ��<�S= ��<�c�<'6;<]g<�B�2=s�<�ǃ�����W���漉G�<�=,=�9���ż=b�<6,a��j=,m�<�Gc��E=%�=�a�;K
�<�Z�#XL='%���İ;����+滮��=�:7��׫9��=4�a=��P=Ɇ���v���f/�0�2=b�$��.<�D��G*�^Q<���<�J�<8+�T��<!��e��;�&�ր�<���<�z�<�4�;��<�;�/��5r�%)1=�U�<�15=ݮ=74�<�J<[�����=
)
���_���S��<&�+�d�R<R��:5B�<�?�<ۣ���m��{[=��=b�J=m�������瓼��)9��;oY��󵆽�*<Hn�<�hּ��G<�'�D4�<FuV=�z*=J�H����vY4����;��o�k�6="�K��F���=H�<����<�Ӽ��Z=�b�wFG<)��V�j8y��A���ֆ��0Z=2��<C��%��<��=�9����
=�:I�?sE=5�Y=���=�7L=Gl����<$N�C�伽5;7�D=\	S=�T���L=�k}�"�+�2���)g=-,=e5+=.�ӻ:!{�U��<���<���<�I��S=5�=t��=c{~=[�:�Z�����mI{��k��kfr��?=�.���0=�5¼�ks<M��%_��8=�м��;�<�<�2��t��<
�4=c5����:��#�����U����	=��L=A���3�����1��<Z�Ӽ%�f��C�!᳻ |2<�I=˳��n���5�����흻�ݼ����9�㇜;�R=�s����;0?=��
 <���G�=�K=SJ�t�h��|!=E��<��Q��R=��7<y���0�<�	=P��؆ =[-#;�Oȼ@s0��q	��$=�{<�ܸ_�=s�#�)��=�S���l�ThG��Kk=ڌ=�+(�c��Ό���`�<c��*�<���<��2=\��%�8=�6O=�雼&�=9:Q=�[@�n�=�k.��B�u�R=�Y;MQO�^&�:�=V���
�<t4�;`s�<$�һ�Ṽ���k.��m���<>Vμ��b=�=>�;����:B�T����C�;�)C=˲�;/EL=oV��c��t�5�Y_{�!g�<�y����;�����;@����l���c?=ʤ:���=S_I��z�=�8ʼ���^����<�p��k���!U��+�<�.=�c���<i�<�����羼�lE=0�D�(<�;y��x��E[M;tgG=��8��D��I�䆱�%FM<�'���dS�*<�%j�h�<=��=��=�e�T�J<T��<�|����<��<Z�;��(��6q�K;��;Z�:~�=�Q����z�����7�=��;�)��B��+7�� ,���<��.�>��8���r~h=$!=�|T=KHT<�ׯ<�����<�@}<�&7�/��<�2��)�;�%T��1&�2���{��*��L�ۼ$�>=O�h<f��<�#ռ�弃�=8�<=f��G����^=r���T	=�W���A-=�=�pV�h�D�����Ҽ���=i�)=ėF��ֻ��M=��;!�]=��<�<�byO<��'�A�!���,=2�*=A��<�t<�w��,2=ʅ<2�C�vh@<�W�?.����<"c�<�G=�g
�ɗ�-v�c����X=݋���ԕ;
�$�vּ�|�����:����(����<l��<��[λ%l]==�)<~\�P�8���=]�q�џ��]�H=�<���<��μ����J漝eQ����=��g��q����tq�<���Pg<��v��S,=�<5ʁ����<���<�!�;��
�Lx<Me5�;Ũ<�ް�SA�����gh�w}R<5tּ�dn�*�=a�����<�''��w}=��2<@	�)��<�1=�H��Ņ���#=�p����Kn�\�;>|ۼ��+��=���_=�\=��ۼ���<�w5=�?�<�'=ֱ?=� �Ms=zK=�~1�L=�8�ы<�����l���P=gz���p��f�<¯;��"p=?X=��=wi<�/=
�"�VZA8�+:=�����һc�C��ʷ<�[6=Ktټ]�4<mc�C�d=�I�<׌���Za�ؤ���+��q<3�;;�<X3�_�{=g��<�D{=�}��D����,�>S-�|��w��T����;�?=�!=krt<WJD<�2=�|+��2�n�^�A�&���_����</Z*=��,;J�m�/�u��^5<�YV<V�R=b{*���㘊<S�,=�$���H|��U==*���!I<�#�
R��1�<������;�t�<%����S>=�q�<�;�����%�=^����ѕ<�c��pU�"q�<�OX=f���=�P�2Y�G&�5W���a��?��/=�8�<�t�<�ﵺ��*�H���1���|��C�<��V�Σ?=|�*�{�H�ID�<�>��.=�?=��? =^����	x��] �h�?�R��;�=����ڼ�<q!c<0Vb�o�n=�K!��,Y���=���<v�Q=M�v<$�I��3+=�K�<��Y�6��<��U�<�O;@c�<�^:�N�<4��<�A3=~����up��M�s��@=w/X=й��V�����=��X�i J<��@�SU�<J�x<��<%~�<�τ:�i:cf�<�=�S�w�W����<�M���x����=B�#�1N�<>p �NQ���.=�Fڼ=={;<� �;&���K<J*�:�d���<ɿ��$==6�<���pw��$^�=�m<c}4<@�;��;�J=�l�%��<��=蒇������ǼG^���9i=y�}��V�<�[a=��E��oJ=:O=��٨���<��";-�C=7�A�_���=4r�����7��<��+�f��:���<̸���w<�$� �0=Z��=�V=�FJ:���<�U=�τ���<��:=9��<l
!;��<���.�<���;��q���3=zb������<R�;�� ��5�<k��ZZM���=�M=��P�t\	�����=F�z�A(D<D�ݼR�/��5'<߶��z6�<&V��#=�V=*և��v����L< %��c<�薼]�<�z�c�A�D�9=k�=�%�K�W=I=�=�2�<L[���9D9F=�Y�;h� <-'z��"�<�I�<0?(=F��<Z#�v=�<�-=[���L��X�	��!=>�i�)@����<�O=F�<�S�'��κ=a@�<��X=���<�)=��)�qV7��D-��kD=�@7=i��<]0�%})=|�r<�w$=�=r^=� ����?��=�H=��)=�rF=洲���l��3i<�R�<������@"&=M\2=�j.<;+Z�c�<A�ٺջ\0b��;����"=�3d<��8��~*�qR=�k���=a=?�ܼg�]���T����<�%�;��л��J�a�y=<j/;�I�V(ջ�����Q=�/��M����o�K����k�1=Y�Q=!��<��=�^=��
�=:�+����L��E�<m_Q;aߡ�/K9;��W�<f#<R�]=��2=��J�P�*�΁�<��=�T�<~�4�ƪ;=K��<ޑ׼�*;�M��w<�w���с��f�J;��]�������Aa;K����bG��Ĥ�D���r�=k��<������Z=0�����5<��񼓽<a�@��!;O@N=�[�;𱁼;o=g�,;��L����P��;�Ջ=��<Rh��w���CM=U�<��$=��)���o��C��
�R�H=}pռ�4O�.Y=��<�O�������Q��Q=�m�;J1=%O�Y��Ι^=��<U7�<��p<���<	=w��;��ݻ���<4]><��
�]\��%;<H�:>�r�8=��=D�,�R�L=)�`��SE�<�>�ڍ�ROf�����<=�4�^�=ŵ�<��{��2k�# �<����4o=n��D{\<@�L�'�	�UJ=����M=R���B�<_v%:�=�y�<و=�vI�nWc�B5<��ռ[@�<]A�O!=�ӫ��H��14����$=N�;=��<u=�0=@��=��+=)�ڞ\=X���{M�������^=� ���޼i�;<�W��.��;u�f<s;:Je=���<W�(�5E�<�2=���}�d�"��JuF<l�0=�k_=�#"�&9�g+�^/T=lO	=,� ���l�9�#=��T=u�<Abk��=�,����7���c���<(GB=�A��ܰ<�d=���:o%8�*q�<�5�<wN�<u=�1=�4h=�ƍ����.� ���fQ�/�h=`��<>��<M�K�r>�<�+�a+�<�U�<�9G���L�3e =Nn�;#:ּ�<�8��Y�j��<��-?=����`�E=~K������P%=�O��2}=�Y�<���3蚼��ʻ�"(=O���~�:b���E
��!"��3=̓�Y�<�Ȁ����<M3���=���:��p=K�F�4�<�F����"<�`ѻ�4E��z|<�A�;�n<��$=\��ά�	5�<.�~��Kz=(���4�=�
�o��<�&<:��<�]�h{���˻�û���t9�<�ּ!�p=f�f=
�8=�L<�r�;���<�gJ�<��E�;Bi+<A�=�wt�/�<�����%�:��<R�Z=o�m��"=S����Z�
���{��:P?�<�uO�s��<��.=��<VdB��=-Ws��~�;��û�Ǽs���Ɠ�|���ڼd��� ������S<�e漖��| ��;/=�=�����<r������^���"�<="�B���<{��r�:|��'-��u��˼b����a �%���(���n=�K�<p����N�@=P��U���+fi�h:a��]���jϼ
��;Gk;��<wԻ��H���K<u��<,Fû�8ͼ���ټ�2;#v^=>�;�={�]=��m��4ۼ�RM����;�g.��3+=��=�KI��C=�S5�'o��7=^������<���;�$��#���C��=�RL�/�I<h�<ws=�ݺw0*��;S�*c�K+����Ƽk�ɼ@��;Ʃ<k=(VF�*�'=Ř�<�V�<v�=�:W��`=fl6==Ż�_�Vq�V�$�!�!�r=K[�)��;�5��qZj�n8^=�[=ߺ����<�a���,�<"��@d=B�|�7�<��'�۠�ɣb=1��<?@���K=�@�<n�<	2*=؏= L;���;K�C�mE�2?	�"�Q<t �<�,;q�=�5t=��I=	�=� �<�t�[��K�~%X<)�u<ڣ��:��;�:��q=j.�0:�;)��%ڶ<Pf ==��:O]$;l���^m�x�x��N=j9���=WƼ�N=5-�<A'Ѽ҉4;ܳE��Ǽ��=��=�o�=c6�:���;��'��t6=^i;ƃ�a�W��Q!���s=�:n�
=��=8�,=�a�7�׼�¹�h=;$��1%=Һ:<�?�D;��A��H�=�A�<�>=���<*⼚�(<hVp�s���k�M��"*����<Tc=����gd=�yݼ�<ؘJ;<�u���
��/u=1궼WG�����P=`tE=-�=�J�lp�<�����.h="�v=`Y�� �<�@<��R���A��@"<1w=X�_=P�#���y�l�<�m�<�lJ=�b��L{R�O�=<��<	KU<SO�MM~<�4=b2<���0v@�a>�<�wf;V�z/=Op=�F<��<��4=�͂<�Լ��ʼ�O���e��,=1���ڼ�Z�I=��=~��<�qg���z��b�V =��<��1�9K��eH���1�<T��;ww ���<��I=�D�;�H\=����\K#=�
�9==R���j�V�[����ӆ߼ch ���<NN={Q���C&<B�ܼ�G�0=<�5=�6�<�g=�Q.=s�@<NP=�:�<۞��0�T=!����/<Nķ�� =����8���<Q����0������X�U�=�n��.=��E��*;z�,=�!X��WQ<0L�J�p=�[f<>����Si<������<,=�<$|=v\�"����t���S�9�=QZ>�:l�.n�<�����K<o��<�>F�DpA=^�9=&ā;�X鼥����)�Q�ʼŭ�B�-��z�< ���V�W�&E�X�j�:CA�U�=�R�<OJӼ��;=~�����9/�:8�<�	=c��<��&��RL=�5f=��x��=h=�)�
��<�e�R̂��̼x�=¬��3=Z���w��<x#���n=o�|<�Z���S:�:1��,�;]!��<�)�����ٗF���p<�$�E�&=ڐ�<g�<��P���1=�&�<��<�$^�������a�Q�ߛ+;u�}��.���]=*.��dm=
� =.���Hw�5��=Z5��/O=
?��F< v��d��qȼ�&G��|�\G;��# =�nU=��
=G�;�.��*U�]c�Z�
�dي==%;?Q=P���b%ﻚn��u�<u�3=%��MP�ï=�DT���m=�(=Y���.�M�<�
^�>�'=�m]=��
�x{t=z`/=u���B�<��&�@ �</Q ;k��Ws&�^^,���"�0v�N��;��<�YG�Дf��/<nBO=ǋ=M}q=��[�~`��Y��/����<>�]�lO��ځ5�����w]�Έ=��<=�@=�����;u�V��幼�:��]=��=`�ļشw=^m�4r�<�eP�ὠ�;�=���<a8�����<�Z����=�}�<e�W>_<�lC��lJ���;�<�_<�Ӑ�;��=��=���lʚ<��V<��"=d�5=,t�q�=X��XR���Z�=�7=�T-=v,]�9�%ؼbs(�¶�<��'k�~N=��n��`żA{�<@$����ļD��=K��;�^�XL��U/���=5
���"�}pj�rC=~$���A=��;N��Y�J=n�[��^��76�?=����'}R�n���m�=���3��;M���㧼ئp=���<;A=F��<���<�_Y���)�\x�=�ñ���=�:'=�~V��H��|=�--=k\0��Y�:�(=CF�;����m�<�D=p�<U�<l������-W=ଈ��,�<@�6�E�a���-=B�_=��B��Ugf=��R�U����<�-� }������0�o���[���u��|�?<�"<��Ǽ/a�;{��<Ϧ�m��<�u�<~ޣ�\7�R�)�'`K<��P;��B����<�K��;�D=!��<v�.=+d<�x�<T>_�����F�C=Ā��?�J=�	��#���Ǽ�}ӻ�1=�[q����<DSo�,���?�;W����O=��7�x���!=�	���-�6��<��==��F��Q�:7XO<N�lX<��;��?;���q1<"�J=F��<�_�<�vs��-�;"�= Q��P^ռ�l}�L �;Bk&����wy<���<r���]�N<���<叹< (��w�g=�>=� X�Qt�:�=5);t��<;5L���<q��<�3�<��<}T��+J�(껼��=���ݠ=�/���i�\��<�Q=RI^�U5!����K|�5�;H����v1=^��:���<�b�=�΄��D_�P�Ƽ�)�<��O�	�<c���;����ě�y��<����U = �<c�Ļ!�'<��7= �=�Mܼ^'�,���1߼�_[=J���gyn���>������� ��F�<vQ���(����J�a�B=M��; ���i�:s\=nI={�<W���=&�5�V J�{j=T$��=�$�<�p'=�^="t=�]=��*=X��<��׼��<4��<�=�=��<��~<�� =Sf�9���<��F���<�5������U�<m�u�;�<BU�<�9�����{.=��\���\�k�;1��S)<��@=�|����ϼ��'s�D�����^<��T�53=@$F� d1�$�9=FSN=�w�:���<�<�<RW2=��l�T ��+������<DO�<�k����_���8;< ��������M=Q�O�x�I�")��w==o=Ճ;�,=�-�J*��lh=P��<�)E�X�˼A/=;��G-=����#P�r����n���k=��i����<<���0=����м�.��r= ��;Dv �1j�:��2<
_�<���H�<.p��~F��7?<��;���<�E ���&�P��<�aS9+ԇ<q����5c���>���]�����m=P���L��<#��<#k�<�j��:<�n��D9=%���:�
��< I=0[�;2�K<���;��<��<yd��?3�D�==MS=]������<�R<��D<J�?=%��;=d���pO=2mU=�9���<�3=��Ǽ�9=��4=�͵�AV��*<�S;"��;~�
��Qa=�2��w����<�6
<��&�In=;�<�p;p��߀=��2=��/=�Z����<��N=�i͹|��+�<����i��<w6�<\+�ݼ��o*F��y�׈P=�Ի�=t�]�v<�<È-����7=��<�=f�m<���;fv���P��%�<6�d=o0*=��\=�Rw<h�;��d�Y����毼ȹ���h��(=�����O8�<^��<h[c���B:���	Ｐ�;	�=V�Z=��FK�<#E=�v�<��W�
�?=��Y�ji�<1�|�)=��Y�`�s�����<�h4��>�,1�;����uͻ\���X=G6y�A��<�݇���:��=ְ&�y�;T3=�0<��Iz=�g��FOQ=�p���u�<�II=^����N<=�h< K�Z�1���!�<fn���7��:�<�;������^�� ��<�~<=
Ѡ���<������<�#!=%ü�Ň�R`�"k��$J�I`1�*7&<d#��h�c�������H7���ɼ���<�"������ނ="N�� �
6�����{����&��}+=�S���&��IH��޼G~9�I�'��~=�<�=��T=�a��y�<��#=���<����U�<����n�bIZ<V��<Ar<���)�%����d=k��<P���d<p�ż�����A�&�d<��j=E��=%�.9-(;��e��YA=��=���<�Tb�9,=W�?=FD��F6�9���ug/�)Ү<�k� G�;�#�<E�ۼ��H���z���t<��ἱu =8Ve=aT=�`1=�ۼR�K�F�.�>@̼w;���H�<8��<�<y��<�<�����=��U��SG=��<� =��L<��8���l��o`F��{o���'�㜭�Y���b,=�@��
�<&�ٺ*���X�J�rjP��6�O+o<��}�U�:�ȟ���R�<I���a�<���<E��b�;��<��Q=FQ���3�%�v;�\���6���;���<���w@��)k_�g�q16�ِ�/JA�^=��t=� =��P='X<�Y�nm�<\m����<�_���w=<���ߗ�:l=�[��:�Z<><=P
$=oڪ<rЛ�Y=��7=��&��{#=O�f���7�m���6��G����<5_ּ�	�<�k}<��=_�&��q�A�e#o�J� �Ӧ��K_��Cȼ�[=®"=�
��i-����<CW<���ڮ�<�""=�`���Uf;���<8�$=�`G=u@�<<�*<>��<q��7BM�t��<�y�������fD	=y򊼪)%=�&�3E��v́��Dg�2�t=2�̼�|2�2`=��^<�d�=����76�!r��O=϶�w=Q<�Q&�c�<�n�'���F=_qZ�˲ߺ�F�%r��+�I�[�<�}�<��k�o��<r9=�e;=33�;$G;�<��*��Ve��Hɻ;*�]<�:@���=�D.='=kV��Ui��/�]��=�u/��H=�N��n�(�ߝj<�=��=9��wg�<���6=����<��G=��'���� =w�<M�B=z�r<��q;�e�:��i��$o=ǆ������C���Ȼ����$��<}C�ZY�=��<@�5=~�,=R�N�$4�=]ߛ��?I��Z������IļPW�<�z��~5��ו���4�t�`��M
<�Nμ %ȼɓ^;��C����s㼝$���=�>;U<�w=TkR=-�<;+7=���<9���aB�;<���@w�Wf��|�28�<Ф��e���-����<P�|��:a���K=�|��弍�>��a�=��<W�����)��M����A�Z{�:J�<�*<	�5��o�����Ply<�3f�+T�������Y��_Y�ǐ��$�;Bme���<�y�X�j�ѻ���<��<0�-=j1k=�(c=i���1�#=���;��<j=��%=����
=�=У���ao��D�<U�=%�ۼHS=�M�<0=��=���;��6�me�<�1���u�AT��\;�^�=jC�<1~�<baS=��;��=�1�CQ��Sd�<��̼	��Լ`L��7<=�Ƕ<�N�;��=0�E���`�{+d<_���pq�<0����fb<��^�$��8�<x"��=2=a��)�S�覭�&��;j�u'=�v�;1f=Wl@=�0=ش�<8[���xn�6��[�F<WV��?��ܔd=Q9��M�;��<�;*DM<�'=�r�S�����I�B��X��/e�<�l0��+=v�<��T4���W��$��9�jq�<�`R=�t=�)A��ޘ�OQʼ��w={�<|5|��eļٸ=t趼�+=yt=Gj��� ��ˢ<!�
=k�Q�P�����<�+���,=p�|�ln!���Q��2[��>O��-��9ߢ�_�;��;�+�:~T=�`�ȏ�w��<�_�JE<1�F�.p<o�1��/=z���8������V���s�=�� ���5�Q=�1y=�
=�C=g�=��<���Ͽ�<���}	=70e�|�<=ŷE=�ѭ<7M=��o<��5���<�j�;�Y=.��JV����.����R=��D=��ؼ�6y���%��͌�7��=>vκ�9��/ǡ�8Ki=��<��ܻ��<� �;� (�t�
=D�T=F�#=�r��mJh��@�=�=��A�;<�Q=ݟ6<�ׂ�%��;A�"={{����>dh9=�)��$��(=L� ��^�<Ɲ8=��=�
=��<�V�o�<݂ǻ5�=��:�B��z����<G.�<=>��<�z=��޼{IG<8E&����R�<;<a��e�<�=;���ӟ<v�=�u_<8b=��<�5e;*�U-=Xn%��&=k-�<j;���V��*<H�<�y�<A�t=o�ż�j��L����*Y=I���]c��<�-�<�%=�O*�w��<���<�i�-C�<�#2=�"�<=/�9᪼���<�F;tA�d�4��6=-孼���<�uO=Ue/���7���N<ucQ�e��<[�$V�8�=ч<�:^=4o��;P����ɉ?���b���,;W��SM�Ϣ/��	=��=<�ZN���F=K���	�O�(=��B =�����<����xK=�E�vץ:t�Z���.<p��=����B�<Da���+���,�;�Fa=5i3�Sg+����<�;=�n4=>ʍ;c��p�e��:�M��8=�!�-�]���0,�=�^2<9A�<X�<rh%���<��5���=�Y�{��<�&�wm��	]L=�7`=F�5=�$;�r�T[��/:)=V[�<ǿe=<�T�tx9���<��8�����m =�E=�~#;䰑<��"��\.�˰8��j=9���鍂�!yK���¼L��<���<~<Ԯ<���<5�/���%�)=U�t�������^�T<FS;=�i�;̙�B��)�q�0^�< �~�k�{�üh'h<J7��Z ���9���0=2}�;��<̶m���9=Y���Ͷ�7�;u�¼�N��s�+��<�?�<��t=�2 ��v-=^߾<�����i�<�
�;y:�����<�t��r�@<�Q���k��!=7�/=M�L�g����>�k9����FS=��f=�����G��xμ}8�<��=�Sɼ�j�<Q�ۻ`=<p����=�Û��k�<G�d��q;�jC��g���f�<
�=s<#�׼�Y=}i/=\��<<�5�z^_�Z���DJ�b{�	v�퉼 �#=?��^Hj�Y�g�vJ=�������T==.�=�����<M9=����kO;���<�#=`�L�yT=gh=8�f�����I�4=�ܼ�@��ÿ����=H�3=?�|;��<2�C�ާ5=���<wj=.FK��;�< ּ�3
����<2:=V[`��l��"'ؼ�;'<�8 =}�E=p۵<J��;X�G��LK���j�"�\�t� ��Ǻ|-~=��<��|�s�<�L��c&=Ps�<TB<�K=��=)�����3�=���<"�c:=#[=�g	��F=گ= K=��=2��<4�4����:E=B�U<b�<T>W��s�<��&<nR}<H��;���1"H<6���&�!~�;�U,=��:<�n/�`b =�D�:uM �w4=�+l�s�!=7�`��PS�0�w����aX��'H=<A�1�&=�i=_����2N=�O�<?�*=��M=���fn�;�/��۟��}�b�,=H<��;
_=�w*��@#=8�񻍯>=��$+��u-���]<���<�g��a�;�K�<=��E�MAO�#�Ѽ%(������>;�8�=�c3<A0�<�<�Ҡ<�꼆QS=�𼜐=kԁ=i��;3ѷ;f�h�����P�9<�S-=.�H=PK��-6v��uH���0;�%� �w����:n�=�μ-?Ѽp���_O=�0j<�T��g2�o1��_u+��\-�v�	=4����R��9=���;�s^<��<C
�P��.��&3���"=�r3=z�9�C�a��H5=��)�-�f��Ǽ���;�!���O<�<i�9�ݼ��;����*�jH��g#�<'�ݼ�,h�CHB�pca��N=�u(�BKa��F=�;u�=�&�M�==�|��c*��:=�Q"����;���<���<u���w=FMB�4�<�U�LP����<=O�=	��*^=�'ּ_����k<���������B�=��=%X�ֹ<=4
e���V��N���������=.�$�?�5;_Ʈ�l��<(`)��|j��(=��;-�<��ݼ��<Z[Լ��L<��;;�R�v��<B�"�Z�:�HF=#�n��e-=!�=��E= }7�^F��"T���, <<�!*�SwC=#��a=1�=���<Z�:�5��;7�){L�S=�5=�~��M_�=�{=���D����h���R�)V�<�u0�SM@=�*�<�]-�gj=�yj�X�	���Լ��<��	�D�=��<�ꑼ`�<ߌa�"��=X�9�"���^�8=2�J�[0�u�9=���;�@�z0�A�K=pVF��g�;{���ڻ�����q\=��:�y:��M9�?�
�=)=E���:�<�`�;�xO<I&�<4����<]~��(U�Ս���<��+���H�z:=�J=6LC<Hq=si]=�G�6��I�<��,=��e=s���?��Dy=�T��%=z,���I<��'_$�V��H��<j`�4 =�t ���<�N���$��=j8��B��6x7T�=2P_=v/���v=�0��X�<'�'�x�<o,��6X=Zv�<2ހ����6b��ZV�<)�=��	=�&�<}|�<0��<�o�<x̑���X=��軇"=��̻[�n<�e,���ڼ5��<M3�<�)��*�F� h=tG=��=�Es���;�o)3<vb�<�� ��⼖�e�l�뻛\b<��=��]��Dj;��ϻ��L��D����҂=�po�>*=��n=ކ��(:�<�����9$�$%&�Wkc<��=��"<VV�`VL��/=�
���;0��<R�
�ùH�K;�h�!=Р�;��M=<̼�x�<x��<z�x��ZV=�v���;1�C��$ =�W�<ă<߾=���=�I;����l�:==���h:�;0%)=���<�ָ:�z :��=?�A�N<�v=�}-=v��<�#�<�O?=�Z<�t<���<܏�}4=Ӟ"=.�����<�</��g,<?i=��ּ-��<ra���v<�p;��;AW���׼�@ּB=�<̼���;�0���V=�Z���;��~�=��)=ٿмY���g�a�f�!v��ns�$��LwW<]���h�5�<i/�<���;����ZJ�*�;�R=�>��[�<����v�;��d;��A��=�<��CEO�!!޺���=G"=7����6=�6=�<�a8=��A�<�"�O�j�Dx`<��l=T�2�Z�+=dY�;�e=��)='�:��ּ��<�r�=��w<��n���M<?�7�i�</�!�1Ud�1�/��`9�T����I.�v	��^�n�T�.=5j�d<�S��<��T�o�r���C�`��m�!=`]<�qh=t�����b�N� �=�	=�٘�2P��o}<^��;)3P�~�׻���u=TZ�R�T=٣�<]��!�@=�=���<a�K�Q��Ѻ =�� <$�;���L�=��#=��S���a<��<h��<�i��#a\=�a=͔Ӽ���|R��<�<�w�<��Q����;����X o�S�\= 	�ňo��=:h<g���;=J�=��<k�:��1��/T<`;��<�3�<L�����<�<5�ڼ�P�i�=?j <ţ	��.�<Xּ��=fqG=�%���2�t��2*�#�=�F���r=b�E���3=Tˋ<�}����Z=	r�<9f-������fm�%�f=�8M���T��6=��<'�Q=?H@���6�\2���˸�<&= �o:���?�==m=�<�(B������T=�]p= 8=������<q��<Cμx�;0��S�A��Hμ[:�<yF�Hr��d��<����$�6�F��kM`�!�d�(.H=�J�<Dꝼ�;Y�h=��"�����$~�<N�u3j�vTo=���<K�S=��6=��
=�)��R�<<�b<dF�=�J��5}ؼ�4��o=$$2=+`=j{�<�d�<�-X=�Wa��ˀ<���;S�����y6� �l��n <8$��B��<_C�j��<�2W�w��<�=���7��}�<�]�<ę(�Nm�H��<l�=�8=�}{<("A�AX����x�=���ʕ�M�*=�M4=���5S>�#�`�g��3�B<P������L��<\~�;��=���8��6��=���;t�̼?$�<�sټ�3���=H3�<�pC�T�O=�D=�X�8G�M��=/Ff=+Tȼ�>�<g�������=@�<b�7<:�U��I(u=��0��@�<�l�<��)=q����;ri优.s�ﺑ;=�<M�����v�=��'�9�<𼷼��-;LJ��s��A���.=���;���;,�;�Rm�<�=��ż�ý�f�!�[q<ux=z�n�ف<���<���7!=I�<�����c�� �<v�<�}b��y=� �<��<�IQ����|�C=w�i�R�ӻ}ʼR��<;Z=�Aͼ�.<��<g�t���<N'����R����Q�(:��=8��;���;���<���<;�S=L��=&I=���<ְ�;L&=��@=������4<�a��o�<E������<���������L���;���4UM�k�=>������؀���<L�6�}W+=y+��=���ϼە��q��;�Cb�[~,=/�;4��Zf�� =V6�<��1�\��<���<`�=o&%��a-��叼	�8�E�"<�=���yʔ���O��p��d�=�x�r=sk��Q<�f=-������<��A=a�m��� =�B�<�S=!4==�C���;N�� �����D� �,���<=��2<�=�BA;���^#<q%�<D��<Y����#�`�(�Y~=.�ԼP=�I�x$ �x�]<�TM9FXͻEކ�������s<$49:�^F�� ����)B�;�-=�hļ�Щ�ɒ�;�v=K�o=O2
�S�=h��<?X�s�=��?<���<��=��;2�����<?��YN�P@=ɰߺ��I�O���V����=�I�]�=$���F��<��;=4�==+H�;$,�ҪO=;ͼ�F=�H<�-q$�?mX���#���v&˼ۇ���׼tA�0s�	��<��D=ERp;S���-����,B=��;=�+��V��V���i���;�:�΍��LX�=���<<��<B�:�����v)�i,ٻK =�$B�)n=$*9=��[<��==�=��=�s5��@=R�<�aԼ�s=�, �!M`=�/���n-=�&=��ݹ�e=��-=�T��a��ی�<� )=���o�ּm� ��;��>�)��<����� �<�$=�p�<9n,� �k<�&�"�<�<<=L�=�r=wX�+�ʼ�0<Fּ�uj=ږ8=�`���<����&�(�e<����F8=�t�݊=���P�c�<N�==�=�ĵ<�	�<��#�A�<��|j=d/a��>�f���k]������6�=�=5RǼTRb=���M=L�1�8��Σ:��Ѫ>����:]�<W�= !�<_ V���6���=�{��=R��m�7��<��I=2��;�4���l=�~Z���!��{o= �;=�b��~��t<䨭;�X��o_�,��[��`�;�S�d�<�;������/=qz����l�YUG=�f�<.�N��=�c=��<<�J=η)<��,��:=f�)=��<�C�����b�k��<Pl�<��������K��:�9��#�;��0=�R;��I=��'<�=�����^<��%;߲���<�wt=�==m�<PM���0=Տh�_ꁼ6����-<��<Th=�� ;�H�G�j=�[;=�O��Q0���<{�q=�2�wK#�ڧ1��s-;\=���<O�&=��=<�PW<�2�;ʿ1�eX|=P�%=b�r�.��<7D����2�۫ؼ,>�<u(^��D��� �;'��<�Ϣ<G�=T�+��<�z�<���<�ۡ���4=��{�m�3�8(��=0h����k�����<3b����V=-p�<�x�<�g=�{U��g�n�=��:�0�9<��<�%����<��=�<m��ڶ=	���k�S�<掼$�h�=�3�g㺼M��;1��`=��J=�P�<�s%=�Vo;�,#=���<��<^o7<�6'=|;'�*Ol�#��;j�l�ZR*='��`��;P�&���A=�T��Kn��[�<B2���p=���<B텼'�L=1#<����_�{=B꼯E��䓿<�dC�L=YsR=-�1;��-=R�=�+��L6=`^���3�x�;�y=�<�"���=�\��I_�<U~=�-<=�^L<��=׃=��!=`��<\@���Q?�l{	<�0)=&h�{t���� N�;�w=��5���3-H�qA9<���.]��"�<?�=<�wt=]�;k�o<��U���S�����={f3<K]�<��%�)F8���2��%�;>b����;�a��T"��Z�t�5<��z��L�ĸ���-�<Z��;��<�'9��`�;i�;�I���&=��>���V=�	Y=�%�vT�<��=��	=��=/@�Z �<	�H���z<����@=	�q�_���$�9=��w<�P<cH�:���It�<3t�[L��u�]��y���<�h�;�Nm<ợ�����%��<���;N�7=Q=�O��6}=n������3��.�9��O<�l�<$�0=;��<쟼��;��1�< �q���\;*��<io��@8=����$y�Bc+=�=fޯ���
=D�/�\�����-<�-q=� A���<X�<yu�<y���ԹD�N�=tɼ��ͼ�,�4�輮��K���_�<�z=�K�+�$=hA�Y�~=aW�<�f\=����g}���=j7��S/1���N=���<q�
�o^3��$<�&I�	��<�4S="м;N�:�L=!�!�bW=S��sM=��<=�9�h��<Y�h���];�Z-=&�-���Ն�L�P<��4=�*"�!�=*�;������A=c��<�2=4��<]�;h�_:�i�@�V�R�F=��>�u�~=��@=��	�z].�W�<�Z.=�;��`�䆌<Dv�G�Y=�_�<?���}�<#�p��{�<"A�B=�T�<5�:��<���<�e<��(�ʷ�<�	�����v:R�Y=RRs�������´�<v���)F����=��׼\C߼r�<��W�Vy��dHż��O�1!�:�\��{5�<��^=j�p=�����=��<�<��h=��:���<)
=�:��� a��A)�.�'�o�ѼZG=��:�{�s�g$_����<�p�;���H�̻��	�����i=~�>�'U=@6<�<]4���<���<`L�vY�<��;�h�9O�� f��x�4��G�<u���k����/�b�;�̘��˅�y�j���1��W�;�M=�K��8|!=w�;���=�U�<qZP�+�缍�<�C��<�ƴ��\�sH�<@h=M7=�2��='<!�@<E���,��q�<4�C=�N;�B�d�<�ߌ����<���<�P��%K=*1�<�1���=d�]M=��d��l���7���v=,��:C!���<��=�,�<@�<��[��1+=y����B;�=��L���NH=Ӥ����<2��e�=��6=j=E��%K< H�<z���_��SX�<�o=Y�[=!j,��*=6dj�8
���4=q�]=��0=�W��<���=��f�Ao�:1f9=n�=[8���<q�F����`";!B�p4�<)���9��o�-=���;{9��4x��D>j<�I��+������xH�<T�}�Ѽ�Ʀ�Ft=�ۮ�H@�<��<�=Һ4����!=a��<�[��ƛ=��:,�g�U�o���B�q=54P�(��*�~=��a<��]�T�D=��:� 
=�+�� ��<��<�8�]�j��n=���y1���ἴ�[��lѻ79=Ղ<��ܹ���(����]��g,���]e�ǁ=���;㤦�|x�������;n��:��>���=�G��4?�<ZM����򻀒Լ�����8<<;�<���^>=�3�<A�H�K����_=Q�
�[���;~�m�B�;c��<VX�$+�pt<�e;����D�u�(�<��=_|�<P�=�=�<+�X���'���;���>�ɰ��#=���<���9�D��E=��Y�{��p�<P��<��==6{q��儼�^K��(=��_��^=k5�M��<��<XȆ����;�=�xr�<�;0H�c}���B<}�`��]4�d�[<�?<+إ<8X��>��M��R���$ܻأ༫K3���n=m�3������c<X�����F={!�<?�B�򫖼�
b=��;�ZQ�CL=�F�<�����I�}b=��<E�=(�X�r��)c�	l�<��<�"<�IN�|�=Z�Q=��4��{'=��L�%��K��<t =pI�<�=`�q=TD4�M�A=�U�H�1�_��ǻ{	���Z=���;�-E=�@P=��=��s=1޻����u��Q���}QR;?�.=�f�(=(R�<�م��F��@�\��oɻ��-=�U��T���6=�dnW=:7�<6��sF=_G��n�q�g�v���ё�=�=���N=c�+=Z��֋(=���!�x=�ч�\K=����¿D<S�l=Θ��w�<'b!=�vܼ,�@<�cz�4�=:B���6���$��C�<EVa=���<^S<�I;��-=uq�<ϐX=�C�s����</�?+�������)ƺ��:U�3�/��H�<ɛ%�:/\=~*ۼ�9=<�_����2� �6� ���bI<�pϼh�==z�Z=WT=0��M=�Y=s�=�e+�m,����
�~Ot<k\=��+���6�������N�%���:֓�<�X
� Xi��f�<��@<�X�;n�f=9�h�k�k=����Q<���<��8=n߄��T������]�<�:�����ټ!��=`nc=�;9t�=1�<1�,�U	N���[<�6C=h�=p���'=��f<|��<#j�<��<�?�S�=��u�̺};61B�&�i<�!�<gc������ 9���<^S=D��X1���+�P�=`T@=z�Ƽ�d�Z�Z���}��#�ڛ_=�-<��\����ܼ�)ҼtS�=	�<"7�:�b�<3c<��)<�Kn�u	"��� =UB%=^� =退��'<�\o=�,�@S�<�L#��J缕��<��f=��~�b<��;�'=w�]��5,���<=V��&{��H�w��������D=�=��=q� =6�r<Ad���Q�<���Ｄ�)=C�M=�,P<��-=#���a?=go7�&��:,�J���=�Sm=�3!��ar��Y�L
�<n�D<=�'�p;6=�㈼K���*΋�2�;�����DӺs�;� ^�<[�[=4)�<��,�r{�;KSe��(B� ��sܽ<$�;����]�;�1�^\<�wX��G{�B�C=�X�<��7`�W#_<��������Ӧ����<n��&R=���<���1���FR+<T��<X�2�Jl߼g�;��׼>æ����އQ��μf_4<����"�;=��=-ϩ��dH=����i�%Q<�Z��J�|=?��<##��
[�>����7�q�4�$Q=4�g=S}=�|+;ĝl�]�`:���<�X	=��;=�L=,�U=K��<�"S��f=}p�s�U��+�=��d�hO&��'[=`�׼c?V��!=u>=�=������<��Y1ټN<O�j����;<�.= �^=�RX=�{�d/�<ŝ1�\F�&Lu=��<�Ra=�~�;��2=�E�<��i�e�׼�\�<�*=�yF<�5��m�<hG���1�<��p=߮V����5�<�W�\�*=>&'�F�
�$#��B��H�]<��T���üf��<�+0=�c�<�hw=m�R=�˫��4�c� �E�g;%=�Yl<��¼Yv����筞;w�0�z\ͼZż�h�<��<�[�<_�S�>}=����h[;U�����=������`=ha���<�_<�~6���m=J��<�G=�6=®�<�AN���]=
�=.���į���f=Jy��K�?�@�E�o�G<?w�<��ļ/_��h���"=
�2�|N=��\��-='�y�W*���K=�Y�ơ��q��;���n�"=@�|��N�	L����̼ӳB=D�L=&�,��p1<�ݛ<�?�R�L=�CK9��>=���υB�GX=f�_��VL���<���=�tH���<X����v�;��"�-=P��+�F=Vx>=�U�< ������l�<�<�<������[���;,��4=4�j<�m�<�μ;w���!:��P=u��D�����4<�û����k>���#�+!5�[S�<1X�<~I=�l�Y��<�(;7m�l������J=��6���8�W�0m.�tU2��xx;!GC�t�ǵ�#	=�yA��мN��Ɲ0�Kf=��<N=5B�<v�a�f�\�;<�:4�r=,�����=T9_��r��[<��<��=ۏ�����=<�LB��CL�sr*=���<���<��C���(|>=A�����=��[<h
�;CԌ=�u����<K� ���aH��0N=xfѼ|V��=��"�i�;R��<;�ҼI�k;m���!�G�4��1=�i漩=Bo=�3=�|�K_=��<��f=�R���cQ������<2cx�GT>��KF<�_=��p�K���������;w�Ǽ۟<଼��<��<����HB�}=�k����h�N�E�h�B:zU����;o���*٠<��1=�u&��zO�f\��4����t��)p=�b�<Ɇ���n��w�a;��'�-��zn�<?�7=~���j�|�dϯ�caȼa7�<]�<���<_@'=�<�(����<�~?=������u<�c��°�e�e=�	D�R0<��[=BL��Ɯ�;�ø�Rr����<�:.��i	�W��+
=D�;�G���<�R�m-=��1=~|#�����/�$Oe����<]x�?N|=�@�GEo=fIE=R}��@�l=ƣ	=ס:��{*;�y��G�D����QI���k��%��G���;h;� �<�=̯��MK-=���<	�Q��P�=LS�N�g��V�M��G1V��Cl<�S1�f��v%�<Ds��=^�<4Ty<��鼠+L�p��:�N���q�<^fx�(
���;�3K=��%=��;B�#=�BO�M�=9	z=��J<�a��n@<���<��=l?仢��<��U<t���3�5�%=5��f�;.�=�F���j=, Ǽ�3N=�pQ�x@=�4<Y��;q)< g6�+�;�h�<1�S�F��1�<�x�<4 d<<F��0��](�D׼�$#<���<:��;�����G=����*/=�:9�FP�<��<9�a�;�¼{���"d�&�=*Y�<OA�U~9=��ߺ��6�@�2��9<�E�<ۂi<H�-=�����/=�h1�j�=������<��<�~ =�Tļ�$�<�VH<�����:ڽ�<�.���X=gD�<�S��ܴ�<�~<1m�:�F��Kg�<r+��M[=��D���)/=�.�6;м���<��<���<z&����<�;\�伒��;\g=��o��c�����<�h���=ZQ�;�첼��=oP�<
�K�x)L=I$�c�������[�^�ڻ����<��,�J�</���D=���<�!��޼sE~=\��<"d�<��!8����=ދ{��%y<�\�<ړ�<�`Ҽ�ȸ�6�S=�����o�<�܎�:�C��HK=��ļ �<���<�o<�h��<O���F����<�!=A���qT=���<'K=�\�<����?t=���<VZ�6#<�"c=1f/�Z�*=ϔ�<�^V=���<�< O[��Џ<�{�<*^!<�>u=^C>={T�<������=��<v̼�����T9<�.�bk�6���-t�=k�=��<�5=ݾ0=DvE=!�<n%=�s<����(�Ҽ��{=���/�3X9y�O��j�:�k���R=ߍ`=�V�2�M=��3=��*=��C��4;\tt=��<;I��Oȼ�f=��I=xc4�FJ�S�r�R�B�7=��%��ϼ�e�����<�<�=	$��Ɍ���<���:l=ߋ��`=5\E<9D��1μ��ϼ�0���,Ҽ;�<d;���>F=?;7<�=�e&=p�R=cJ:=�84������)��q�;N�ۦ<�覺�R=��&�V���P7=W!ȼ�J<����=Ԫ��#�$���ݼ���EA���I=�A��rP�9-=�| ;G���/��<�ڥ<���9�Y�l=)�.��N��@�|pX����<T7<\*�;P�Ѽ��=Y�H�~��6s<�ۥ</�2���|<�����9�<���U�b=K���τ���3�jQ�"���A*=	a�<$�<T�C=���1-=4(�]�<�<Y=��<8J<��KP�YwH=��m<8�;5�<@!=|
<�A=.[�I�ѻK��<�}��g޼X��;E�<��z������C������;=.p<_kY���U�:��<�]�swϼ��y�W�G:V�]=Yљ�6�	=�b��!�^<V=��2<�6�K:5<�dM=����$S�>��<*MM�����.��^=];�V�<���;%0f��c��>5�(�:=�ˎ9[>�<�=��(=��<
p켬���V�����9����<;��;��$�z�M�r�`=l�p=�J0�ґv<�<wmG�LD��
�=��<��|<�M�|�L�wN�( =dS��	���<�f
=��`�����>f=t�;7��<d�<Qq0��3<=��o����^�O�~����ټ���+n��� ��5@=�n�<�6(���<yȼ"���=y�@��Z˼􌌽�r|<�i�#ƶ���f<�hO��?�=<l�����<���?�<'9=Y�f��=B�I�%tu=�q�;?K=�B���2=�+��$$<r�(;����]�*���A�g�#=#����=�l!�������SJ=��W��;����}r=ʏ��f:����e�F�T̏<L�<a�I�pٛ<��+=�_=`Gn��QC�l$�<t�=O�L<DzO=����[<$�~��>D=TS����2<��:�Ӽ<�+y���=��c����=bU#���"=[+�Op=E�7��<�ؘ<uj� ����=�'��rb��#�����<��<Iϭ<Z��A=9=#�3�2z<<iT��|7=�Ɔ:%��
�<�5��2˼|��G6�L��<^���+='�=ʋ=T��<�^�<w_켽��:q��<vӅ�t�'=&�����<�GU�1LA���<vg=[_J=:;����<Z�<=�߻�`�Z=
�h��++�(Uu����<7��
��;��*=�78=jS~�?�=PZ껬v+=^��;�$���@$<��p<AC<8�4=�m.=0h+=ݣ���ɻHtF�&>���c=��<���;�=�+����:���ude<��h<�d=诱��:6<� h=b�j��M3<S ���Y�Ց#=<�L=ڊ^=c*�%�鼨c�;,�\���:W�0=$'!=���;	�����4���'<��Z�Qԅ<A���� $��{�4�ڻ��e=��3<ucɻt#R= 
�K�<��P<n�=��;���kF:<�����<ب-=���*K<�c�(=���R�`�������<�)�<G�5�D�<�t=�� <�<�/1=�03<��!=��q��(5�R�
=��l���=]�<�9Ի� <Q�%�M6�<Yu|=X==�Ȇ<_=f�=	�;Mx5=V>v<�.=B��<P��ņ���=X:����o���J�џ<��g�;�	��~q<nK=&7D=���;\�<l4�<�,Ǽ��=��ļ`ix�BLt�to�:Q�<�I=�8=7�̻�cмV M<���E�j<�Jġ����=ҾH<�;�<
�Ȩ���)�9���z�������ס��4�<N��=�DB��3�/�J�������9=E�j=g���Wh;��<ǉu<T���1�.���	�M�=V��<Fp��9&X:ob���=Q��4e<BL���=+T,��=,=~H[=yF�^,��|��=�=&�I���n�L𵼂I�;X-ӻTaI�[P<�ŗ=^���PQI=ף��Gü��7=7I=��� #�=2 _���2=Q�5=G����N�rIe��~Ƽ�@μ���8wj��6B��Ep=6%L=o�<�&G�� ��*�<_�y='�]=Z�c:���<+�����&�~�5=�Ix����<O�(=�F��k@=�p��
R=<Bf�+�F=Ҙ`=��=^A_�x�=79U��S�	cмX#P�{-�;�����l����<Q���<�Z<cCW=+�=/����e}���Q�2�8�?=����oN=��O=-sI��2�<��K�Y<M�;�<��E=%y��+��<�x!=D/K�����<�X��
��Ӣ|=9��<хm=����8}���9=�K�<'��������=Q�M������<���"���o�;��A��j�<Rͼ�p�<�=%�=�'�<�A�򨖺8"�<��<��м�W*��%6;�ē<�o�=Sj=��Y�>nT�[=��<ߣ:�zo �cY!=����q7=h��<�{
�X
=4���=ѶJ���<U���kZ=��R�T1���������X=�)�8V=)dl=@�><��z���Q=�� ��(1��}�;/YL��r���0=Q:�;��_��ܕ�P�^���@=��B��&M��u2�=$|��=����	�5�}������v�<���<�(3�:���6=ÛU�p��J=� �<���<x�1=SI<�N�<1�=��J=����C��q�<�:��-_K�Zl�<G�a=�'=7w�/A�Hś�WV=J#�<>T(��є����B͈<�+=.|�<@On=ƈ=s&
==!��MӼ4�6=�%�C�0�o��;�/���9���na=���<��K=zJ�<�9��Ἱ��<:DҼ��N�˝
��	$=��b�]@�<�&�ٗռD�L���Y���V��7\t����μ�H��C=D,����ii�<�u=E�4����[W=!�F��}�<pꉽy�=���ȻX�<����v��"���J���iD<�I�<��9���<K�f#� =ay�<9�g=�w\=�+�<h���ߚ���7?���<i+=��;RU�Ȟ̻B~<�=;���n�;�<=�Q����^���p=�"�=ڻU�R��<�=>�);^D)�v����<�
Ǽ�6�4u=X�"<�o]=P��$cU��C[<�Q���j�}-��2J�<P�=x����]�"2[�y����#=P�O�|��<�p=�L�d'g=�U.=�"=N~8=y��<M�=�F[��i(=:Z��;�<�'�<�'i�}��=LB_<�Z�;i|�~�� %���tػ�(n<�!���<��Y�B�<�LI=a�c��/E�� ��?��U��{���|&=�=y�;��8�@��/�<���;2E@��_��n���Ӽ_̚<�c=�Z���r2�튁<f_��l�ͼ�QO=��1=�-�u��<M���5��
��=�<
+p<<���W<�t/=�r�<� �;ט"��U=���~�|�16��<!E�'��=(F\=�Z=
=Y�缭�ݹDռ�����5���
=���<�|�;S�=u�<�
<x���i=Ck�k�+=ʬ+=�KH=�̼:�>���v^=����P�h��3v���:5�m<�0 =�)ɼ����I@��G_<!�"�0��<,bj�Sߴ<y�\�SP.=��B���T�)��<��X��A�<�v�<N��<IdB;5��<�ԣ�|X=
=�q=<RR'=%������a=�i+�-C��V^'=�kq�05�(v9���U����y����v3�D��<,QN=[�u��.�<T�=+_%=LɄ;Ϧ��C=m|���=m|<+?x�k/�<�q�9>�>:��z�W�3�׼��k<o�ּS�3��"=�/ �P�=?��X���� =D���E2�{��<�\ü�L��~7Q�o�f=n���/IC=���JC�����^2<#��<ps%=�� �Q�'=Vc
�:�r̼i&�:��������(=
L�<ԑR=�
=��\����6p,<��A=��y=O��na��ڷ<�j�<!<�<�x�����<U��f�8f�V�6;��a�+�b=6�e��_�;؜Z=	tK=zC����X�Q�K=�=��<M�:U��<�FS= ֻ^VO�Ƒl�ź
;g�<$�8�Z��<mڪ�&='	�l�<؃0=7�4=4mN=�h =ps�<ɲ={y�< l\=<���m��颼8D��qn�{M��B��<�p�bO<�=+\`=l��<�e��ᣣ��UJ�5�y���+=��=��=�/v<�D�:i�h=�m3��=3���MIk={�c�6����.�A;U��;J��;�$�M����W�<�Z\��'�:�;�H!�e���1=�����['�<rʻ�c�f��<��^�<�8�<5-��p�<���<��<uu*��=,�E=��=�j=P`�z�t�v�"���J�^=��<u��<�7�<��<�M��H��<��2��M�;tvu=�>=��E=�K=��Y��|�<p�#��5V=Vo9��<\�P���{���q;�8J=�D=��R��hܼ�t=�Ǯ;nD=��;���</-��˗<�\��-Mq<��p�=�`����<m-
�%�=���J6=�Ѽꢾ<�{�<�\Z�s|=Ɂ;��
 ;��9=SS}�"�n<��%��;�^O=i��`�:=���������gFl<���|sf=*i�<!�@=�A��Qj=�K�JD$=��2�
�ü�A��ۛ<^@�<A��=e�W��<������<��l�d^`��q=[�V=��;~���ze�I'=k�B=��}�:\=V�.=�إ�ۺ��`?�QɄ;@:�=�5�y?'�AXO=�^K=o�<��2=���<詨����<F[��n59=�g�;{�L=j'B�>�U=."<��J=��&=���<πM��jԻU��<�ۏ<���<_B%���q�ۼ�����k���E<�0�AE�<��&��"�ľ=��=�y�D(<a9�<)�L�t1���*�ׄ�<}ú�
���=^�4=�|5=H�<T�]=X�[=�+�+��d8�:	��%c�<��-<�|=��v;�N���=�8=р��<+=B)�<z�(=��C=�P<��<��<^�`����e<ּ5P��w=t�N�<�|���<�Z'_<�X��qn��a�<�M�<с�</��G�2��A��Y=+=,�<��ռ�Պ�T?V=��F=��5=6l8�fjB�R�=�=X�=18	��X+; �=��(�2TT�~
�<ڈ	�G��<�EX=@��Bj�<��m=N�=�B=�;ƻ���=�)Q��k'<��u=uON���<�]=�N����.��H��^�������<�OQ��u򼰓9=������%��p�<lR���=$�=�̼;�"=�~=$�A='k���=��Y4=����y^D<!�?=�A�<�m�<�j�:��I�������i=�D,=)y��γۼJ�qg1<�j�<>��;)�W�D�!�2�=��<�!�2���ꟙ9a/_=Q��<�_�;%�=q�� �	<�9(���)=]̲�y<H�L=���<u�<Zp:���=��x�������0��S�<\�&�0���5=�F=����.�=���V��<����s����J��B��%�۪�Q� �|=9�Q���R=�@�<�'"=v�<��i=��%=��<��C���I=y�);��D����<+��<5μ�>�<�Rb�����5�0�ח_=§(=�e�V�"��9��[<��q<x��<�|���)��C�<t�Y=�^=�	���<=�q*=�a=�T<�=��E��<I		<]&;`�=�3����;�<���e�;���;��[<
y==�D��"=�T��".<�ƶ���T���$�95=Z3=L�X�0l��S=����ϼ�ǐ<�!<�9��;a~��5���/;;�"������!=t )=�����0h<+p<!�=�$v;���=9b�<�썼�ℼF�<Ûo���<0�׺��W<V{-�Oֻ�^���<����T�ܐ�;��%�e_��c��<��.�P�̼6�G�=E-�0���&=��~=v��YL���Sq=�1F�x8���1=��b=ˏ�<K�#���<[q��_GO���*=��D���D�gm�<�s=��=7Q=Q�<�l���9�-�I;9����:�"a�)�L=>���^S=��=���<�?-��Y�=](<}h�<�M=�+�<J5ɼX�	����<�k<n�= O���;�Nr<+�R:�<f�T=��E�K�<p�7<w�0���W����<�OP�}�&=�2I�S<14��ds�� l�����^�ӻ塺<�'!����:��<C+=ܫ=��U=P �[�T�J������h!=�u�g�Լ�	+����<�+�<�q=I(���ND=��鎻(f�<���<,��<}�`=a�u=V��Aμcw�|�l���C<��<��T�5���y��}#�k��<�����up=�U�;m�@���<�b��G��2�=���<�R����< ΂=t�=؟0�Q�׼�G�����<Ť�<0j�;���cL=$�)<Q!�X����d  =���`�\�d0L;�Ý����c�!=��<M��<�j=);�<�����;M�m��i=K�"=d==#�N�ۚ;�hѼ{�<Sw	�r{�<��<J`=�י<��[�߼3VC=�S�}G����<�"k��e;&�e=�lպ��s;H1ջ`,=����</<�w_��g@<�ӝ��)N=��%;�H��ML��`�<��,���c���f��	��,M=�k�<se�<^� <�S=^=b����^�^�K;���T-=�s=X�;�һGV�P;���76=#n�<`X�� �:O$I��W$=3#��\�\:���=1 =���	1$�e9���pN����:����3�i���>}�82�J��K���;�0G�g9��,f�<�q���zZ;�)B=�=ꗼ+�k�`O`<OI�V�ۼ��J=>��<�ż`�;�S���=F^=�j�<2$@=;�=��X�4�F=J�a��Y1�Yh���F9=������:fl=�#��k@<��<���<c����z`��!��ģ輷���)>�#C���|�S])���7�[���]e=��=m(!�^C=�����T<����3à�-=k�̻�-f=����e����
�Ѽ�=/V[�ˌ�<λj�<�`<��Z���ϼ� /���g�Ö{�`=��{�+G�<��=���:�
$�⪳<Q3=]9Q=�!�<Z����X_=+hl�R�V=���<������<T�L=�޲<��CE�*��WZ�,��}D=�v<���^�W�=�w;=�C0=���:�*=Ql=��ؼ~��ۻ�U1=fx���Ϲ<~�1=VHd=��ؼ#���a	��B�;���<�w:<��;z	�<�ۛ:��<�Ͱ;v�<��(���a�!������<�҇���X���=<M_�F��<���:�0��`�< d�<��U��^>�8�<�+< Ka=��Q=	�P�ƻB=4ѝ<�<����]=�;?<8��<u;�<)�&=�_X��r�x�>d�<��E��\뺵�<��a;�1�<̬<�������-���R7=��=�d�<b�=�0�<�ͼVS�a�=f��<o���:c�'t=�P�<�U�z_:<���<j���f��,�Xf<䋽�=�$�R�W<
b"<��S�K���u�=q�(= �c<LS=o+4��M=�U�<O�;�/:��-��{,=ԏB<�J���6=�K�+�1��h'=�[2=�ȋ�s9�;���;o�o���<�(�2�h��(���|���=���;'(��+��%<�	=�ˏ���<$�=]=��K;��ܼ8��i�4=Nܫ<�vݻCr+�Shv�[4@�����x��6�:=�Hz��.h<K�D<�j<�En<�_���);���:]H�<��R�Ƣ$=�mB=�*#=�OD�B�>��j8��L��L�:�h��Go9=�h"����m�(��H�<���;s�6���<���<#�C����"%�<�Ǽ������:���S��;&���+�1Gλ��);i��\�=�Bj��u<Tt�%���d��u�&<D�\=ܲ�<	Q(;A췻�;N�	�;��ͬ<Y�1<3�M=�<=����{;w=�����I ��T�#�W����:�cƻ�|��+<x&>�I.:�f=-[=$�<y�ڼ?ݼ�B=��h=�e��ؕ<P ���6�o~�c<>=�ZJ��t���/�T�<堼<z�:�r<�d5��3�m�F�MY���<=kE�ˇ�7`���ͼZ���>�<�G	< o��)�l\.��O�=~h�<�j�W<5^�<��a�k8�	4����]��=����'Y9<�}N=�w�@K0=�׫;&ޤ�9���}lV���;�I��Qݘ�Fx�<;Œ������=��>D<S ���ǔ<�&���Y��R�v1`=�\_=_�Z�}jɼ`�(���Ѽ"�.��:��Ԃ�og���p<�]M���M=,q=b�-=�tY<6��<�������h�n<|sy:0���z��<��;�m(���μS'=�k�����;B��Tf�z�<�ؠ<�.P� B.��2W�q��<��[�/��<�=�?�<7��7�5��Ž:/|�u�;�U�=}Q���.�Kr�8�����o=F5� %��h甼N:����#=FfN�mGD=��T;��<�7�<`j!=�x��z#!� ���IѼ��O=/��6L��12������T�����1��λ��7=w�ڻ�;�8�=���<�Gg��a�<��3�W�x;[�<�	H=$yJ�9߼�8=; h=R'=VF��=7 =9&�<WX�\�\A@�9�+�x>��1%=�Q��wL�n?�<{�ռ�"#��pO�7�Y�	�p�	><�J��eL���=���<aD!�!U>�	F�������=Z<�<)�-=h{9�ܨ�:�򁼢��<WS=H9�K��𙵼mEQ�W��<��9<@!<�NB=����Yۼ*�J��ҼÛ<L���^k�������.=��<�H�=�T=�Ϊ<n<�Y�*�=*Z4����*Ȼ�L�#+-�g���ּg!��#���s;�lrD��\�Ւs=��]<���b�<���<�X=j�;=�.d=��;/n?�1�=�tE�T�4��i�<{�c�^!
�1�=r,=m����l=#ļ�6Ǽ�=aS�<~��<i�R�P��Ƭ��c�5$=8�<�'!����:�<��K��@U�A?��C�<o�W=x�#=��K=/H�<w���y�=�AFb�ᶅ=7�;��@ͻp�(���M=;ZӼFA�;�FO=��C:1J��'���X=�֪��bh���z<F|t=6V6�����~D1=�%�;ʧ��&�=�ü�����C��1<ǜ�<Sּ�b<�x�<lm�=��<�w=={�=�0/��
�4N7�ģ;ko< u������1=��=֕�<2���n�<:�B�އ��-Ƽֆ�<�'+=�X=T Ѽ!u]�a	z<<J��07<CX�:J6=<� =�8����w����\�",
��ռa�<��E�p�<p̎<>~M=ͯ�<|���+<Oߤ;+��z����:���;����<��6="�:��t�<��F�bƤ<�=�f�;j 
���h��C<��,�Z=�띊�d7<]m���=SX�<�K;=Q���MԺ����;�:b��߼h:]T\<�=*�i���Y��v0��&�;�<	�;6��o|;=�B���);_�=�u�<6�<j�ڼ��'�*/�<�k�7�0�|��ڝF�*�K=�O�<*��o"<����=�u�;fj=��^<Qs&��=��Ȼ�z�:�<>��GJ�#Z/=�v�^��<��M�iP �3}�:�1��ZT�<@��8'=��><��I�6��N �?���
P����<�h%���<=�;����G�=%�:=�
��F_H��.=V�л=�V�pM4�8ZҼ:-��7#�����j+<ƾ8<��b=jLF�_0=]�:�1 =4���{�
��S>��@==�?�<L;H�B=��g���<4Z9==�<�#v=�~<o�<��C�ӂ�������<H�߼V�m��V=�r�Qlb�I[=�EP�����Ti<���<f�q�~Q�<��<��[��3�<g��M_i��{T�Q��<�Ŏ<V%Z<�=H=ߚ<DȨ�3/��Q�I��z�+�d<z�(����<�ak;ԽU=�c<��<u�= �����<:���d��ڠ:<��;��+���==�C�3 P=�5=�.=u#)��w�;���<N�Q�+�z��-��=�QD=�_���}=�
=0aG�/`�<e&��.�=qF�X�==$�;��������<ɳ�֓=Lӆ��d�<�`<��4���(=��&�8=n�R�X�=z�<K1�;�\j�I�=QP��G�<�E��zV���\=� s=VJ＀�N=�-?=>D�"2&<�����-��"i<fB|�+:���;�9���+<ѬB���K/p�_Ǽ��<�kp�x�c�+N񻀁�!�(=A��X̼%��G6�<�_"�&u�<���9�N<,�:N�<qw��	���J&�<.�;F�<���he=�M��r��<��d��:]=�! �=�=1�<�����z��=YDj���\=��;;r=�
L=�ϙ<��=PN�9�&=���<d���Z����}=U�<?��=�:��3=!Z;=��u�� K=U��<a���N���8=g�{�#]<�h��9�p��e�_�8�]��G��I�<��컟�=-J=/��<M?�<�?���o<�Ҽ>9���*=z��xaN��7=vpY=�l¼0��g�;<>.<�dI=��<fn+�~�)��0��_\<"Zl��j<��=�%��i����<b�p�U'��3,�<6*㼄�$���=�<ն�;@ݑ<�8r�н�<;�ٻ��X���
;p�E;�$=��;����BG=��ѹV6c=4��i|=�c=��<�8=Q{�-Ci�@�f����h�;m����<�%�Ϗ�<n�<N>X��/-=��#r2���9=���<|�%=���<`G<�S�^�����<WԹ<���<mYN=�p/�3`R��oF<�L
���?=">=0�x���<�#�<�4U<w�z��W��?�<Z�j=�u6���L9Z=*=9=�ϝ<��ܼȮ_��<����iԮ�\M�+^a���:��=[����)=�	='0@��d�W�������.s�{J �o����@���<N�::<�y��>�<E�<Bo';�-=?�/=���<}�;�<B<���E�uX��C��y�Y����S��+�-�y�<�.��j=�W|ٺ��=qq�<Z�J��<-�(=��Q����������<���&x�����,�#�'�,<����N�'�=�m=F��vQ����Ƽ�5=��3=�;�_�6�ޗ4�`�K�;���</��.؄<�]�<�jn=��K�#��<1�6��~��o޼:2:=K�F�9:��M�v��$�<կk����< >�<<]�4�mie=��μ�<r��N�=�K=7l<��=��;D����=�_Q<�^�H����	=[4�9�
�< �=Lo�<�i-�&-���19�1��<�l=9��d-\=
4o=x&����;2�Y���5�ե�:���<�;�(@=��Ǽ��<�'�,�<�I����":=?�"<���B�~=,��<��]=N+�}�|=�b����|<�w=n�E�uY<=���<{�Q<�����)����Tr={(��w�<S�2<9�;i��Ⱦ<��O=���/�0=� �<�C�4N�<��<)����<j�Y=�������t\8�3P����V������/=�kc=�%#���;����4�����0S˻��*zO�V䈻���=H%���y�����B�B���W=�Ȼ����)�{ ���B���d��3=	�8=�=�}�<��;��T��C6�
��J���S��%&=�(��ּ� e=���;62�<%��f5�:�j���	=۠G=�ab=�v���v���E�<�P9�v��=���<��?=h��<�7ּ)�e=�&�;���;=�v�}?I=�)=�-6<���� ���<+�;���^�S<�㘼j�<�I=�u�������&A<��;j�=�7��T�Y��<��d=y�޼e17=2&�d� ���+���	�"P�Jl�v�<r��<�*=aU=y��<r�<(ke��1Ҽl�Z=M�D=�!#�k�;�_��xN��T;=���<��<<�w ��LS��~'=	IL=[TM<��=�x�<K�p;�&=�Oʼb=ahq�2�1<�虼X�j������
��=O<0�|<+u��0���=���<K�)�Ǫ��(�=�M���FlV<O�?�'���O=?�1�=l� ���O�mX�� :=j�2��<)��43=䈬<h�9='�8=�m�w$1��}�<���:���AN�-�J=�����t6F��뀼S<�Y�)��<l���=�����>�74�<يR=]bټ��$=�B!���Ҽc�0=����_�̷b������<=�+=��<)=���<S���ss&��H�<sԼUM=hm��
�+���%�[=�>�;!����<���}�@����=|�M{R�2%=L�L��=@�g<NAK�k�;��5=��=x((=���3�k<����:JY�<�Y���q�V+=AP=�0�^�м��O����8=�D<PlF<��=%*��PB�ĺ�Oy��|:d�A�<y�*������<��,=�Xp�t�L=9#=T���E<�j=�'$��]=��H<b�<9�+=��HH	�cI��S��Ԑ<�+߼�����ϼzf���?�<i��<�0<=��I:�i���D=jl$=rI�j=��S=��9���n=7=����� ����=����is<x]���@=��<��\;���< �$=J:�<	>�<{�n�ſ�$�9�.�k�I8����@=��<�N=˱�\d�����</��RK=_�)����o5��@K��px=���<Ln�:�I� N<��h=g�1<xOo�T�:��w=[]W���:�G��<g���2������=�cJ<a�ʼ$��<sg =%d=l
���{=-��<P�=��=T�<\���b1�:��������{�X=|�;=�]=j}�<��"<o}�<�r=⻣��e�<3=x��;/4������L��;<=�����ё<�}M:��Z�7=N��$�Cݘ�V�k���<��<�zE�kgֻ3�#�-E��7
=��ɼL"����<=a�pLD:��V=�^B=Y�T=�9޻ȨW=g���&��I������:м����W�:��Q��F*�y�'�pf=!������'Au:�})�)�{=��
���?=6_)�TFۼ�T8�ۿT�h=��_<[q:Ms*��Ά<�a�91@=��h��C =��N=�f����<�	�<S	T=(��<�q,=���;ϰμ�����<6����)<���<������I=�&7�s�h;U"�M�7=)(I�%Gn<x*�@�]�5�8=`bü/�����-ʋ����;�E���D�O�S��;	�<�P<�H=I@�;x%��V����� ���)<���	��<��ּ��l�h<�D8=�r;�r�<Hi��Ud��Q[@=��?�?+=�*A���;�d#=b �<��H��*Y�H�"��o�߱�;x��; ���+��;]p�<@��� �1<�0���6g=[8h=J�'�AT!�a�}<�4=��v��<#=�a|=Ղ�����l�һ8X=�v=N�G=֖μ	-�����h1c=�z���g��R�:em��@=�hͼ���8Y�<�=��u;é��ꁼw@�<��Լ՝̼mm;���Oq�/Vb�e�g:I�5�>�;a�ɼ�מ�u�-ÿ���=�,5���m<Q�<�21=#y9��^��n�H�UiѼ @q=�5��aV=���<�=��s	s�s9�<=��$=�NF:2�B���#=l.=��H=�䟼m�;�H�3n�=��=�.;<�@�H\=��T����ۨ;=1F =���<�I�7;ݼ[�K=<�'�^�<_3ü�`.:|^��Rr;����cP�<�Z��������{=���7=����ڼ;��<D�Y�v_=��h㮼>�=��<Av��E<�<M9��-8^=��Q�g=U>=�s=�P�M�3=�	U��}V<*u�t�û�a��fM<��=Ȟ���3�QP=�#�y�'�B�޸�Lἂ:U;�m<�D=�H�k�M<v5�<0��<$�?�a	�;�N�6	����⼾Ǭ��].�õ.=4�P������i�(�'<��&���=�HԼ׬ؼ3sn������ol=��ռ�F=Qna�-8P=)�'�cr\��c�� �<(ju�j"I��ԭ�8�=<cCL�7�-�"�X�B�_=Q{V���`�N�?=L�ϼ�3��3�3��*=wK=7��<wb�x� =&\��*	<��j��A<W7������W��Kb;��"@�A/�=�兼hh���EG=U�<�
=[��<Q��<��=�+=���<JD=ނ����=��3����:���Df=oY���b��q=D� ���Y�-����M��v�Q?���������n���R��X��ݜ<bp=��,=
�=;�Z������H��#<��)���<J�\=��u<��2���%=���<t�� ـ�=ӣ�X]$=�H��{
=�1�?M�juM=���:�$=7yܼ�\=�+���f=�2���$�!OټQ'�<6`�<6�a=��<;E<)�<��_=ѭ �����^�<IZ`�J ۼE�p��8���?|���Z<cߊ<����}�C<F����]7=�:�<�<= $�<���;�:=$d�����y=+�j<�]���j=v�����5���6�E����k;�&�=�%�<�Ւ���l=�!�;��9lM=�Y?��w�<�;�>��\x��RH����.==y���lV���)�&i?=
g����e�?=��=�6!�͛=W6�|�=�+	<��1=�(<M	�/] =#�O��_@=�P�<:�<}<�d�<�R����<W��<��\=b$E����������<�M�<����A\�� =��P��z�<��I����;����4=;�'�]-<�v�= ��<7;9o0��7g�5�9=�� 뼼�}��ܼ��-=	}9=��<$Ԕ�	�Q��$�;`��<�a=:��<�6�^���N=��<�5S����;?�s=t�=���AǻU-5�O�*<>A=�Q��\��=�Y#L�/։��=<M�G�t�g=D;�<�f��{-���=���L9���`=U=�=�h��+N��m=�cV;���<d��er:<�=�(=�Ļ7ѻ��
����<�h3��j�Dx�3@,=i"Լ+�+=`��
�,=+�:=� =��<�8;t�R�n
$��8����<Z�`��W=���ns�-6>=�>���/�h���7���	�X����k��0�=!�P=�2=��ܼ�K=J�<�"f���I=��;
�+=+�E�Z�L<�M�;%k��G����T�4L<�y@�P���D<�j��r\e��E������w��R�]=��<�
�:K�=;#9��f�=沼?���-Ǽ�+���=��;4�����c5
����<���6��\=\�<r7�<ޤP=�5<�QἩ3����9m'=���F������;�;�����&�;J�мl[K��]Q���0��%���m�neW�������<�k��L�>=�ż;Y��뽼'��e{�<6!<=Df�~_n��ɻk�=lA��Es��麼D�&=Y��p5�$m=�|���	;���_�S�Z[B�_�9M۹�m�=E)�	5�$=j�<��%�P?��ZM� ��ρ�<v)�z�4�
֣<S��<��<5)/=!=�
��	��
_��1�b�\���l�ց�<B�9�X��������'=Pb;��8ۼ���;�pV�My=��<=��-=�=&�3=ܿ������V��]++�쬖�c3�<��W<�'=�l:<š= w=h�Y�R�='�;��+[X��TN=RT��Ku=T��<sK=u0������jO���<x�\=�X�����Ǯ<ΟN=D~����<�aD���e=��[=�}�3��b�x�޽ =Pi3=�to<�"=��B=�6V=*!=(˼m�W<|%<���,�<φo=�j�<�@Z���b=g�2�Ww�<����r���ip;${4=��ɼ�u��I���8=�*��p�=FT"=!!1�_�>=�(�5��<�:=8Ba<�nx�e:�:p�y\�_��=3��/���h�<�"4��:;�@P=ϡ<h�y=�u2�ձ{<�`5=."�<���qQ���<a__=�:��٥7�?���b�!O�<�8T�Z)μ��5�	�Y<f讻��b=;��=���6����+��#�y<��<M�����w��8�<��:xx@�
m�<��h,�*�=��3��w`=�����c=׿D��K�:?YQ=C"�o��%E�<w��
��<7��<(�N=�=x�ܸE\!=�E/�y�<���<2h�<�r=��	������+k�:�T�otn��G�<rC�<��<�1�;(S� �&<*��<66e=�H�;��B=(?=`�
���k�w<�_���
���$�v�9 ΅<�T='��_=e���o�=�s��\�_=��9(�03�#��33:U�9=��載[k����<�=�x/�"#=}�<V��<:`j=W�-�l�<o=��v��a�N�ϼ�w�sm:���+=�h�ziS��Eؼ�+�3�=�-=��H=�����-R���\=^`�<D@=�r|��Q޼&��<�a~�5R����}=)h��s{=�D=�"I=g�-������m1h�{c<Q/<�Q_;g��5�D�K:}��T0���y�:�>�<^7=#9�<����yr��J=.	:��h<B��;�����2����;�dF>=̼��G��<|�<�E�;� +="2'=ԇ���	=�y`=8��{Y�<;���J��a���\�J�����;*=�jR=�@=�ջ��4���a�� V<eͲ<�K�,0=����NR��`=Fa9��*K=��9=M<V�j���+���i���"=d<Q=�'�<��=���<E��<rE�[mC=�Uy��:��<�	'�{���+�<<�f<e�<���<)�<)X<^Y�����;��T��^2<�g�;2@�Vh���=e��<������<��<��g�>��<k�+���غ����:�M��<=���Y�.��f������=�
�ɍ�<.���<!��U�@=��C=�a=��t=+�K��<���<��,a</v<G)�}����<v�/���(=���lL@����M����c��qc=���N,����|=�$�<�pƼ��7�%!&��S2<m��eiL���y<�'�������D<��޼�Œ<d"=����yu[��N=,� ��Ĝ��"���<�q=���� X�텦;�iD=�^�Ik��r5ἨZ>=�]�;�&z<�퇻��<?�\=�6�]�V=̢���<�D���#&=^�!�A�,=��q=��<H�<�Z'�[��ӂ�<�5�<���<�� <�G��y-�5�ѻ�	<D!N��/=?, =x喻]��<Q�,�c�
=�I���=U��`Z=��<5w/=������ü+j=�  ��a�:)ﹼ�,�=촼lxC=���<������)����<��=_�R<L"����j��;
�4�"�3=�Z��Ξ���=�;�kK����<]�J���˼|PA�?9�=��e>��:4g=�5z<5��<�Η<v�4�%�;�/&=\O{=3*<�"��4�)���Q=��H=�9.=%_�^�<)����>#�O=�N`=�&��==�u=��=C�U�&=J7f=Q�/=Mc��
=Z�x�<G��i!�<6�$=q��"�g�;kY�<Jaq=�����-�ЊR=�LA<��6�yў�gi�<�z=�ɻ~�@="B��F�<,��A��<B�==
����;,�;K���ɝ;�I���Gh�rw='\I��u�<�v�[S=�bǼo�<�����p��2=�洼0� ��c�tR�=�-�Q��l��<��(=�l�;}tj<�]�;�?� �Y��
Y��y���Ϲ
�=	�;����bF=�U�<���<qN$��.z�0�<�os=K<M<ѹ>�p=ߑ<�I,�Y9ؼ��'�	�/=�/
�>=5 a������!=5��;z���W�e�a��;��|=J�i<��c��	��p�����<P�;IUl���<��ݼ�3��6��Xϻ��6=EhF�ut[=DP�+~�5���Q=/�<)��C�F��9���:|�����U�r�=)��	�<��1=�aμ_�ռz��W��<	�<�ֻ��.��o����_<�¼�7����P<��<��;�$<�~�_�<7�������p<ă2�m��<O��c�i<��
��\)��M��`��+dC<���fL�;���;$C�R�<o�<<���<�-;@�\=���/F ���!=^����;��H���<��M<��<7z<H��<U�s���:�1���ny�1�=�j�W]p<2�<@�8;K�_���2=�=3����r���[�P��<[x`��_	=KҊ��I��{�=rw�<��;BU�<^��?��	=<wf=��}|��=�$=?Xd��=���<�=�n�!NK��0��j�9��)�� `�y
|��bZ="�=�����ʱ=�6�;c�=+֖<a��;x,N�G")�߹�=-y'��I��3������=={��4z�8<�5:�u�<�92=Mg꼽 =��:��/���L<y�Y=Z��;��]=���L��oȼ�1'�;�!�΄�D�F��Ϫ;Q���C='�<L'T=(l�<oQ�s��<�?k=X�����<W�y�)�E=b�+�I���k5<ÏI=�@���� �;��<4O���T�S��~Wt=�l���r(<�+><]1��P7=��U^+�!�����I���r�<�z=��=_-��_[�q�!��0=n	뻣{A�=j�8��.�'��z�<e�[=ts:�N㼺�4=k-&<\�7�E=��C<�A�I<�<Q;p=��BJ �zU&=(	�4?O:N2D���(=���<��(=I��g�	=S������G�����	=���;�.=^]�!�߼�)��c8=�/���
=���<`ߴ;���<�&e=%;��P���<-�1��9׼ =*�<Y˨����7�H=(�a=X��Y�o��	���˷b<�	�:�>���"�;�����S���~�di=.==?�=�?�<�=1�x=ƘZ��Ro�Ѽ�<�0==]:t�_�4�V=�w*=�W�+��"e��'�o��UHF�p� =H����N=TvH=�$=�5=�������Jd�=���#̥<�I��M�P���{q��y#<����y�Ű����=#�<�5ʼZ�Y����2�E��_Y;���<�h	=���<�L�<4�]=$/���j=�"e�G?=��q��p=��=�xS��<��Ly�ޅ<M��<='�<G�<�;=Ocӻ7(L=�fE=��=<��9���;8#b�ؚ1��k7�"?W��E�<Ķ�I�=^�$�����5�����<��R=��s���c���	��<W�W=+.���Ҽ�:�+�&=�#���P=i�<�3=�"
���=�_O=��4���-�Ȫ!=�$Z���������vf�T`[��)��5�<N=�u�׼��X��v�����0����h=�ԋ<٤G��b����=�Ｋ�=�<"�{++=��o�Yl��}�ϼ�m���ż徊<�=���;|c�<аN�Z|�;y�C��-<D;�>�<�h0=�j�����
=�ѻ���fz	�V$ӻLr!�.n�<�?��e����6=7=�q����<�Z<�_�<H���[6=��^��	ݺ�T=h=�9���C=)���tfN=}F��Ϩx��M����h=>�l=�7}��l ��3Ժh>k<,��<D ��t��l=e]'=�`G��n=�#H=0	��B ��U�K)/=b��@�Ӯ�<w$=��M=��);��=��=���r�,<���6=�P�; lʻԵS:hň��\�<�μ�*W���=��<��G��tP���<�n=@�P��&����0�=��!���;)�^���0�D	�0�:��;L=<?K�E%	=׳��z/=�r�U.=�׼TE��4U�Y=�a̼)�R���=)�8��P�zl:-'�<]|'��==�R�<f�U�@�s��jܼ�'=TM%��_;]&�d5�<�U=�#j=�k��� �:Q����	���=�����v=Vm;=�V
�����*��E���g��4.��|���
�:��5���<��$�PZQ=K-M=��3���&=q�T/r�h�<�O@=�v=.���&3=�>��J.=^���Q�����<n <�[�#���$�^=��"=BPC<�.��x�<�^<n5�<5����Ά��ؑh�
�^�Msh=����f�g!��nU�{��0c&;���<zǼ�	�<*�¼�t<Ɍ2��=���:n\D���z��������6=W�B��y]<�F��E0<^���B=N�����T���R�WA%�<m�<*��<�;J<G}ӻ! !�f�T��,=;�><���o�<k��D��8
={�q=�ռ$'K=N�J=��Ǽ��p���s����<��=~Pj=8��<�w��f<��=���z���O�;4�+<6[�o<�y˻�w�Lפ���<E͕�>��<P���Nм�=/�O�����.==�P��;@C29b{��=��==w8e��V������ܨ���b�ǆB=.n=��,����Co)��X�*\�-���ީ<�k(�:��;��R�A$༳����a��<���<�[����(=�"��}��<�V�:�L=5G!��⋼��<��v�+�7<���r*�<��a��KԼ���<��!��d�<~�t�qu�:�ߥ<�5�<I2�<�l-���X=.e=� _=�M=��X��#�Ĕ�<���<ݸ�<�;6���_�1�z=�r��Z<��b,W=k:l=7�~�cD���
�\��<K��^��E�<��+=`o=L��:
k=�=nXP=�3h��D=Qk�;lE�<#](����ꓢ���&=m�b��-˼�\ڻ%�ɼ�< <������&�ļ|YR�nv=�S0!=�$ü��$<�pz=	��]"X��@j<��ڼ�&�<�Ñ<]�=:�5�$+��-ʼ�6�v��m�V=,�漻=���<��f���d��ɼу:��o��zR���&���E�"��;�*�.6����M=n=���;�I<0�<e�;�[=��;����yI��zQ=����Z����E�X������ũ��*<f�P:�c�<���I�=��
�^�
��-<O6�<�v=�^l=�\��X[=��3=
u�r<��-;	k���a=J�==�O�<%�j9æ�<��g�u�1=�A=�l8=�(�<:8=g=��v���i��������:=5{༟�O=���K�D=V���i��-�=�g�����&�;*�B��=e����O����;�U<]a�7��l,�<i�YC�H=��@��V@��3Ǽp�%���u�D_,�O
��&�<��l�7&��
/�<a��=�Q�<�U�<�}¼���<�7[��_�<�N=Z�[���+����7���q�<��^=�@=>��<T��3rQ�����$?=�mq��M�<�P-=�R=FI��X"=俼���@���=���;v�c=F�<`�=�;<��[���"��ێ<Om���<$O,=�{R=c=&�?<�:>��46=N�u=*�i:H9q����<�m�;R[��X=�<�Og�����'+X��D���:� �<��:�!��5{<��=����۩<A�
�$+*<j�<L;L�/=��q�$�&����<�3Q�P2�<�L�<e�Z���{�Ͽ�<�®<��p=���<�K�<�C�<S�#=�����-=.�=@�ӻ��<q&�t(�)Ҽ*E}��޼V<c� =�uC=?@4�e�U<�����'���H� $U�ʳ�+�X�(� ;�ͨ��{G=�;=f=��=�����l<)�<�d&��?�c�<��;�#[=��?=B�:�<d�EaP���|=D=o%2;�A=�����U�׺�A:�a�I�h�;}������g�u<���ͱ<�&=1�0�m�?= 1b<^Ȼ$=�6<��;��.��q�kx�6bN���v<�+<c�=o�z��@=�a��	xໃ�b��=���P�!�E�u�C�j��<h;}���@[�'d��[���V2����!=Ĭ=;@�<����e�<�i=�V�<5S��흹�@�R=֐<�;�p9�W<�=B=3c뼘,<�$#��:����k=��"��F=���;�c=��<�n�9��`=TiD=��$<��Q�4��<?�.�&�:�ր�~� =�2��V8G<"}-�we�9N����SL�mQ<�y=� ��o$=/�Լ�����<��=�Ǵ<2u��&=mJ�����z����<�9�;M��$ɼ-=u�u�9b(��Ya<*};=�/�< @3�v� ��١<��/��/5:X�5=�k=����1P��ů<ޓ^<�`�H8=�W��PK��,�<��[��:�Z�g<��d���T�k�P����;�yT�Z��<O[*�q. <�����cH=3e�[����T<�=Nb�ƾ<���k=6��;����,����9K��a�;����0��v>6=��<Y��<t���9�<<&gм�B\=��=Q<=��;��)�g=�{=��k<u��r�9=���<�$����%=�к;_?λ�l���L�7���*��;X=�[=�^���ud=�kY=1���#�+�K���;�~�<���<��P=�w����r�h��<���xgb�WGc����<�I�6P��ڂԼH�O���<5����bY��L�<׶�:��n�� �������<$�=�� �9�S�^����=ӫ�;`d�� V�<�O=�k��L�B_<�*�7� �Eg���Ć=��%�Q<���<ץȼuyͻ�<Ƿ=+zҼ��m=�=߽�<J}�<�f��ռ-�u=R� =��9���"�zo��t��:B�Ǽ?X5=��pIc<��h��*Z=Kh���e�0���.�$�/<��/=�w<*
V��'�<��&=�g�<�ڀ<;5]<�9+�i׀��5�=X����1�6��<Me=@Ы;���<�R<�;�y��F"	<�V�<�==���I�AD������,,�8JD=.&=诃;�9w:� ������s9��$�|���ǉɻ�=D=	[�
�=:H�dݐ�;�Q�=O=qr�<�u8�3;Z��)<�ta��8���e�;�9μ`�I�|H*=$�?=�J˼�-�3�T={�<oDI�|��;�%��M<�ܳ�= !<��=X=�ۧ� &=)4W�Iz=�HӼ��<�.�����[�kE�1xf<g�<z��;�y�j����#;�aW=�e����j=M���9\<�W�<c�<kw=�",=ޭ�<T��,�O��vj����ȝ?�
.��=��L�ڧ3=
���NxK�xD�{��ހ�U:�1�X�=`���=�@=xy
<�ߨ�k�`=ɟ�<k3<O$=b1��v�|��B�<�k=$�<�X'��@�Ty��4�:��C��C=bc=)�9=i�!���@<��~<�(�<o�<e���I=G=�<���:�d缪�<`��<��;K�r=b	=�+5=�����Q=�Cj=ZR�_h=��=f
P=�&���D�)�|7�XX<P#O��Ȣ<�:�;��,<��h���`���i;Ц��:�<�n~�z���%��G��2=9p4��G:=��{֏�=I<�?=�l�<U��+V=��}�X���Y,<��2=�bf<a�H��*<Ǌ:�D弶ذ<X�̶p];���<g��4�<��R��>|Z=�
��=�=J�1<���<>��<��<�x=�޻I4�m�*��q���{��H̻"#=�S��k&=i�D=f����C��D!=�P<�����%�<�<C_c=eP�y�h=�0���<��K=�N�<�������?�;!�C�xI�;Ex=�K��#��_�������
���_�<����,S=��l��	(�>�r����<B]E�o��=�D���5=+'��t=.sK�#׻���<����R������p���g�<�Ŭ�zU
�hK����< �G<��g=�UȺX_�=�kS=5��i�gS����<ڊ&=OQ=Ȇ���pS=��L�Q=KmA�d���7�����s=%2�<L=?q��ܹ<���<;	�;?f^=���<�(N=߻7����9�Y�<���<�F�'<Z�(���	��<J�'�A��l�=�)�Ư�bZ<��﻽�=��V�º�<���9>`=.�:*HM=�q�=��;�+�;_�$�!=y���L��("_<�7��"�+���N=4G.�b.�<A�c���,��;�~P����<�*�m���i��(߼�-y�ѓ,<\%<(��I�m�c�5`���	�S�-�W�y�P;׻a�������ܼ��i�ɓ����<���<��
=8ך�l9==��ؼ��`��A����N9f=�[��%m*�f =L�=X{�<��<oZ<e���N}:=޵�X	�<qԮ�Q��!�#=�uh=_g�����<$*�<�P=j�@=�c�<'z���d�<^7T����tD<���<
��r��<�҉�"-�/i��Nq<9F<9(=}�2�s�S=�Y3=wZS���=��+�)�E;a*9<'���	=y@����t=NI���<���5]P=��<���;5����FP=9�˼�=�c<p=I�0�qlc;��<��&=<9a��_H�ۑ�<;�'�Z�9=�9<��I�r�[=�䀼�>��+)�ceV���t�����u;.�W=�j�8�<��|���;�;�����6;N���76�
�#��k�;�{=f�м��������hX�P��<g@���#<<G=B��<���<(fѼM<=/�ݻd���+O;��B=|o���1���v<\�T��$���0��@��5&���Wj�O�����<󷭺n_����E=]�Լ"y<�I���v�<��Z ���p�ׄ]�/�;a+$�	`:��8=Us����0���3=��̻*KQ�;3=/�<�6=����t=▀�%!Q��(���g�=�>=]*R�j����<�p<��\������=��<�	=o�'= G<���<i����e=�p��	��<a��P�<L2��N�u�w���i���~=�4��+���ED��#�=��=��<T.q<������<�ߜ8���WR�@eǺ��t��f��#=҃7�ɇ1�%����'=�f��z�=���h�A�F�4�U>�;q&��A;=��j<�x�q*4={�ڼqPv�sf+��}��aw��s!�w|���<��\�e{K�YH�<����㼻K�<�D��rAY�������@
=�'<�@��8L��I����U���=���<ǃ=��;u�h=b����IA��n�����<-�g�����h#<�r+����;�vr��Rt�BK�<�`-�oKM����<�ļ�x���j����F=#	�TҬ��n'=|����$,��G=��=Q=��nUr;��¼�z��"�5<�4�f�
��;��3e�;�=��:m�</hY;OSN�Ϭ�,�̼��ż�fn=��[��l�;}N<���)Ab<�[�<;�#&=�}z=��N=�L7==B���;8`=�I$;2jl���E��4!�'�g�$��B��>��m�==�7C=ټFe���Bz;�  =�L=�rW�kE��~��Ş���g<C��U1�0 �<����?:lw(=y<UY��<�}��~�hG�J��b��<�Լ�M�<�4��`�<����گ�<FQ$=�G�_+$�>!�<r�`�ġS�J� =X��	l.=VEH��P�����e]�<�+=6'<�˷��h
�!@���*ּVu��ꌿ<����Dʈ<U��n;���<*(����;{�;f=���9�&C��`�<���E=���W�<�O =�8%��[�;B����x�I^�<��M��U�;���u�/�*�=iN�;�^�5P�<���<uB����=cnC���
���<%_���5ż%At=�O�:�(�<Sl�<	�=�zL��W�;eQ���le<�����>Y�D�?SY�w�&��;A�������\�ڹ�<�?B;�=x�n=G����,V�D2k�f�=��4��G��5I=Q� <��7�U#�����+&�2��<��j=,��:����\B<7�#=��Q=qa�<�%�9��$�#Fͼг4��#�<=�ϻ	�=�hJ���ʼ�,� q�;�5�<89m����
�= �U��<��=_0�;�U:�`�<#R6����=-�=��=��b�GU�
봼���<�&�<<ʏ��P=hx�<',��l��2������aN=��@�a��xݼ���<�<)���#ad�7�^=��4=3�\<ɞ�:���<�R��vT���<��V�P|=�
=*A#��<���v=ݴ5��B����;�)=��d=XK<#Z�<���<a~<�����;w\���_�hR==�q=�K<��<�[(��n�lK=��t���5�I��=#�y<����.Y�nf� ��;�m�=�����Ҽ�˾��E�< �޼ÝC=\�H==k#w<)�U���&��%�6i��X�L=0��`Q=�==����A<6�<ʅ�<7�n=���;__=���ؕ�<��Y�p��<��Y�t�<>�������&=R��;��n�����5��W��<�/V=B]�-�%�KR�=:��;�5���j��V=h�����C��n=�j��r.<� 3=�����ӥ��ߜ=�@�<Y���---<t=*�ݺ\�wY�h��}=��b<s�0�(ݻ7M�<��<�vt=�C=E,�<KC8��D�<�<y��jҵ<�<�'<��F������V�d%=k�M���Z<��;_k�Y
�<lj��h���;:&�<5��<�=#UK���?=�"�S�<S�b暻*�(��yv=�/�Px=�ࣼ��i=c�<���ƺ����c=�������$)��N=Lˍ��<�3�=W�=���c)=ݒ$�c�����;<�g=)K��C��K�<w+�)�R�P�a�7�(=s��<�r=��2=������0��;��i<��S:]q�;���<r��;Xv
�wJ�<��<�M�<���;AK�<�"���qC=⸃��@@=g�5<�����N�7��<�)��
*ּ2�E��1�FG�m���mB\�H ��r<�k<�1���K�<�u�=�8�6*��M8��g�����r!�;�T�<y=�#�<|�<(�l="�6���Ļ���=X<2���5���Z��"c9<�3=�/P;�?�!0��T+�C�$�JH}�n�=�
<���<���;���<�C$=��k=��;!�?=L�<�&A=���:߾3�xt����*=�+�[�e<pt=�Q޼�.<W�s= ż=a������+Z =o�e��cj��6���v<7�﹓�_��<��T=�ǻK��<��M=ċ�<Ge��(��<�O?�
�<��}�l��=��5�e&\�0.<������"=���<�(k��VD=���:�i#��܇<y�*=u\�BF���-=��k�	~��F1=�K{=��i�?5��-�8�S��<���m�<"\�k�"��Pe= >�M)O�PuD=��μ(㫼�Q0�> <��,�l��� =�6���O�9�&��7��_:�)=�໑+�;<=�F��}4�-[����
�*�����[�1���q��<Q򵼃�=��Q=�9���	�=��<��Ѽ��x������ü�#=�� � � qg<�uB��P+=\�>��RD=?b��'�=2��-�<�0��G�4=�&�<��<�JT�Ld��ǽ�s^C�}k"���0�&���=��==�>8=?�@=�O[=6W������6�,��ܹ<(v��]<��|=��>< ��AL=�\�<< =E;W�H-m��?r�u�	����<����Jż�|=��7<<���ߌ伍a�<36�9�:�<]��6��<a�>��.g:�����+��B���N�<s!�:�z;�B�W�=��=��1�M�u=��|<t��;VoM�6�:�ahU<aI,=*�$�{C�<�ȇ���`�SY������^g=�K�<�1����Y=<����5�S:hq;��=��1<B�=��<Ѻ��W<��-�^�X=�S���^Q<'�#�}<ڂ��U�[�]�Z=?��T6D=i3?=k�L<�{:=�.=��X�����BS估v���<ؾ<�}=c�3��I�<��<���<�^_=�N�;1F�y7�;A=`��}=�7=eI�<r��<*������g�&�����B�*<�m��q��;�X=P	a���<h3=��)-
�A�7=N�R=�z="e�Z�E=�a<���<,F=x˼/=���� �>=%��8i��<#�O=v�N<qz���eC��a<Pl=Ω滶��`<ْ��O#=;2O=�'%=��.=l$s��h�܏��5Q��c�Z��<&�ļ��Ż�Y==������<��R���1<���<<�<	27��EC=Q��<@>$=��P�̯H=u�o=2�E=q
�;�Bػ���:;��<iA�<�F<�i'�xqg�*�;��$�;��<<��tyɼ��3�7;�!�:߄�g$�џ=�W<%쐼9��<��!:���<T�*�P4��ՔҼF�m<�	����$�ƥ�[��<����UJ|���;�!Z=c���n�C�~���&�<��q��2�<��7=t9F=O�V=�cF=e��<g�Z��+�<r����=@ L�lv}<*�^�0�h��e�<f�L=��<1&=Qf=��=�~���dR�u�:�s���=Y��J���o1ͻdw>=��=j��<�@&��s=Y |��:5�uu=�=9���R;��>h);�'<�.C�b=�<�Gz<&a=O(�<I�`=� �9Ń��ԜD�m���{�D;��)=�$���r=�)�<,k�<�,�J���>=��<ϸ+�1��`��;�l*�X���_L�<I= �t�_+=�� ��[e�"s��t���;�R���I=]�ȼ�S=oc͹эf:�g=<_�
�(<�2�;7�"=-+�<R��y����;��ȡ;0���{Ǒ< ��;��q��TJ��s=8�<�=H=�tQ�{^=�T5�8瀽�Ȼ�!�|�<u�;�13=|�<l�)��$�;���<��h�r�d=����� �G��<N���<ݠg�c���8�3=���=<�%��%��<3�<� =�'ļU�'={�,��mT<d�U�h�;�w=k�O�^����g�`�F��w
<�V;-�=m.I=J�<�;UlL����A<J.�yG�"ě<�\���式	(=�8a<V��;n�T=��Y�2O�C=Xs�;��<��#�B�I=�f��m���G,��c�;&�:�:}<������<ã�<>
f�A�޺��A=�q=4G��R"�o��`ٻE�e�".�u=�}�;%�S=���<��0<�d%�<�v_��ӌ<�C7�m,-�7	n:��]���&�����0h�5�	�/��9W$i�`��<qD<�A����f��BpI���=�@�p��:��;7��;t?�<�2=�B�<���<�=�Y��`
�g��<�$=Zt�<ǩ�:�|�����8h=<�=�u���<	�=m��<��)=�|�|=h�=��Ӽ���V왼���b����=�t��/A-�
򍼼 �����`�pc<<�K����J��=���	<���W�< �f��F�}k����7�_�g��_=t�K=��b�XV<Ћ6�\����<�41<�Y=vм,	�و<��V=Ԟ.�)�=F����="�R��m޼a�Ȼ��^<X!Q���|�o?X=�A�[�)=JiG=d�'��~���*=���<�#=jlM<x�J=��T�0߽����<��?=�q�{�9=S��rޞ<a�8=�>$=��,<ОD�J�8��c�<�u:��wU�*�n��m��j�f���.����� �<�s=[�1�0YS���1=,,`���=4MW��7ֻ���֍�:%H�<U�o������R�=�k=7�(����۫<a��};���}C�1��=�b=yp1���'�`��Լ�=����c�=u�<;���]����2�/Id:<�\=��D=�-��9���=�������üW�<:���rX=�d��'*�f�J�- ޼�L��E9�z��=�B=������<�<�!�����<����h����<xc=_���4[<]�P=�)�<:��<�w�:s�6=-�H=|�<��==ֆ���=��=��X��)<=T�<�b�<?/.=�v(�+Q6�,�<|o����<����<�����;�<����<�P^����^=�7o=�
�<�od�=H�5¼"�
=�H-��"=x���@�6��<,~I��>�x���K=&�|풼r�:�
����<M� ��~Ҽ�T��]�5=�٦<�#��ws=���;��[�9=z�����͹��{���ͧ=�KaF��Q���=%}G=0�1<�7%���;j�~=�m=k2=�q8��K=z�V=8z�f�V:�q�<����b8�:x��<��<�<���<�)J��/=�;i?��e�-���1����G=T=2OA=�j��Z=g��<�=i<�<[�a�T㨼���:o6�;�F=�NC��x�<Y�=�%��E�L<���<��-<�o�;�dF=�'��q���Dp���=�z�<c��<ܙ�����è��C=�s�Q�Ǽ��<=ē��d;P�<�{�;/=�ą��@v�60?��2�$�<�ϼ3f�0��;)�=F.#�Am��h�b�F�;}�<��=��<s��:V =�~�����^Ļ4$��
���J��4S���1��	4=!Nk=�==\��<!
/<���-l�*Ā��W��=-���ݼ���<�39��O=��<3R��j�<4?=���@�<.����z�Q�)<�q
�()^<��=����7=�w(=��/�T�:��S=�Ƶ<D��<+�;8<R��竻Ѣ&<`�=_�ۺ�(=���<Í,�B��� �߷���;�3�ud�<�������6P$�Qf���]�'�;��<�v�$��6FC<pj���t;�I�	O���e=�\R<e�<s����;��Q�q���ة=�[����<x��:���a�#�|Ax�#M��[�����<E{�	�3=�%�<��*;��X=q�����<ㅽ d=z��<�$����<@��J�޸b<�����O=rr�������q�"�S=�D�P�L��7=�]�<e=W�O==��;�>G��ۼ��.=�]e=�%�;�Y=G1[���<K6)��[<�zl��32�z�j�' *=kʃ��zc=w* �f���9=�Xs��#<��7=-���jἃ�;�����=������j�4���>�"�k��u%<W¶<��M��V�������^=Hc���=��~�45?=�KP��Ǽ�t-;T��\���:�<��<�I=.��y=���<���<�����$�j=l�=(%���J=	ba����?�K�+=�UN�o�¼�^=�V=�=�}����d3K=�{��v�<�.<��K<%�=Bm6<=�=�!T=��^��M�<Y�y�w�$=�nH�ͱ0�%Mq=��=Q_���ܺ�<�=�f=C�=y9��,��<=�J<졼Mj=.x=/�9�[�y/,=�{�<��<��W;��<�S��.1�fHz�e:��lQ"=�;<�D=~�񻤇��U��n�<σ�<��6���<��<O������BH=�p
=O�i=bX�<�����_�Q<S-X���==�+� מ<H�=�Ç�9�u�;�м�v�y;=�)I��*<J=34���m���+��9I�`���3��Q�����=�G��A�:#8r���K=�w'=�e���"=�����;t0m=�F�4,f��i(��U=�4Ƽ��<R�Q=Ǔn<�E���"-<��;�ҧ�D�<�p	=.�8�8qW< �����:=Κ@�ʐ"���b�����&�Y�=��<�C�:�����#=r�7<��Ȅ.��Q3=����;�.6��1:=��2�p�6����<:�3r�9Q�<t7ټ:3׺j#Ƽ0�Z����<�}�zv�n����E����<�ȵ<⟄��u��=+mv�4�?�S�K��\��&0!���=���� [��[=|�~�w�;x�u��+����\=��p�|�=ѨG<��<s#��+�<q�!�k��<U՟��Y<��;�4�<!q5��`=�'=��ܻ���<��=�l��B/<�D`�8�<�W�V��^+�.(Q�<}]<�L��6�<B b�={b=��2�5dD=��=�\-=t��<���<Db2=NF%�������I��p<�l��a�RX=��2��b�=t�u��M�߀�h#��:�<�����U���-=OH=ɠW=8^��B=Y��EE�'��<�T�;	&��A��<�,<w�<x�S�&&�,W�<�'O� i$=J�;�{?=o �;�'�s��<�*�^1�����l�<`V�<솼��*{o�~�3��� ;'�u��N�<sH�<t��=��9�c�=96���炻0,S<����s�oȖ<~�L<4�G�`=�3���XټA)��O=��9kv��ʝ<^�=V?�<>�=x�<z��<�Ga;�PR=8d���=Q^=�:=z�)<��i��/<]��<�	2�m�<��;�6�0��'�Y����B=�\\=�B(<�>�i�w�g,�<(�5��������<i�c�p�@=U촼�HA���<�W#�)�|=�6�%�!<���9I=�mZ<Uo��`�;H�o�6�*�?��)<[=�����"=�M�|�=
='=
tQ=�JX=Ŝ=�dJ����d0=��6�M~y9��<��Y<��y=�k�wuS����~b=s,����	=�T���<u�A�h���nO���h��Y=]��<�n�:"U=�x�G=�<<J-���:� ,=���<R��K<=:�sx�Y�b=�$$<�~�<t�G=g?U�~T'�U��m�;�1�\b��vռP�9<�=w�Z=`/���=>�<6 @=����%:��z�
�ݼ9]*=;�<�@?;+�Z;xM����A�N_A=)~]�}�=:�;.ē=>6�45��=`)��c=|]�<Ǆ%��V^���<�4�;�lI=F�������v�<6�=7P���\t�e�/<g�s=O��<MD=����3$ʼf�)=�mY=WN=@���W=0���/�=���<���G}��e=�Z�<[i=�nN��ȕ<�<�fȼ�!�h��;*w<"��+��;_��<I�<��;��<^5>=��^=�$=�4H��L=��;!�t)��ܡ8�����j�߻�s:��%��K<Н=/�ԻCp��Q��rt:=�G�<s�D�P���<���{<kf=�bl=��	=N;�E���y`�<��E==57����<�v��n�+���a���Z�J�=>����P�Ļ�Kɼ�X�<�؄�?�<�2�P����������<m�}�}�z=� ��v����d;%���U�<s���;�/=uC:=rX�;�ȼ��c�3�
=�Ǽ2j�U�=����<zYn�@7���!��FE�:�Y���O��:�L ����*�<���H�h=�-�<�M%=��<���<�H߼��a:x��ʡN��Ƽ�b<��H��IC=Q������;kV�<�C�<QK��&�<�W1<RО<O��Y�x��+=J�����ѳ=�i�<�zM���=� ��ڟ��GH�����<��N�P�:[cV��=W�$=��M=n�<�腼���ף�V���=K9#=��#<ʋ�뾠;���k�ؼG��<
��N=Za�6�^=��2=�; .�<�(�<��;�s<H��N�;H�:<�<*��<�B�h =�e~�馆�F��;�a�;���4�=9�<^h?���<��#=��2=k�^<�5=ނ���=���f7:�Q:=[Ka=s�Z��j�;��
�JY:�~�?=$,Ȼ�E�]=�'�=���"�Q=\�����/�D����o<��=8�<s�h�g^�=��<����I�<��u�w��<>�?=��Z��%�����\��@X�&]�k|P={h�;\b=ڢ���0=^^�cN��=3�=���r|S=�N�;dp)��ň�:w�"����.�99d=KO==�?��㚻/�;�Nȼ��<��m=fX�<_6�;�Յ��a>��K��y�=-mO��A=������uq���'A���9�J�k�ד%=2�;��ӻ��=:��:K�;��<@)����ƒ�;��=��'�d7,������6=�Ɖ=�&7���==�0<.�����u;�C���=v)=��(<Y@�֨#�A�O��f<b��<�R��m=Će���`��Z.��'S<��M<���<�"��AG�/��<K�<�cE�U!J�aI��϶<Җ��%D=Ӿ;js�� <=w��;�1��"�<���=�����2.\��������=��:P�5�$�i^)�Em�<�W}��)�<��0��e��"�<����-�=�����F�{n=��y=-k�<�_�<�һ<�a}����nԼ�Y��Պ<���<&d�����Š�<���<�7�<q�<�=�Y�Y==X����:��������=��E��n<bE;�9gN=�=����O^=F���;��=l'=�_�<�*W=�t���+=�?<_��;T��<��W=
�i�F��;��=x��;��;���=;F#��{%��@%��\@=1�O=	24<b3=�о<a�9=��z/����'��@�	�B�`"꺿�;���_�ümv�=6�F=�GN=��<#/=	��.�=6Vx��%�;�d�<A��lDM�V�R�	ז�t�'=R`h=N��������<���h!=�+J=:7��4R=���:ď��
�=]����/=�i���^=g\�< ��/F]�<@ӼX'���g���G=d����:�<x�Y=���<'��,��Ҡ��&�9<$n=��<Z4��z����0�Gɬ��T�<5S�i�D<TH�r*���K��z���H=��s���<�yR=ڲ�<TS߻�? ��:�<{����F�
G9��)�K�I����<���<�󨻰� �!=�N��~�<����U�<��!<�y`<.�y=��S�D�;�z���a�0�d=�+7=��<��_<(��<�;��}Z=�5��%Ѽ9�<�A ��U˼Nm�;�$[=\��;����7W=�G=F��2�;,ST����<7�$=�	�;�}�<r�;��;�bV������H�X��q^<)���:��h�<�*=���<CUQ�K�*�u�;�A^�FvF<�D�<$c�<��x������<�ݾ���;�R�<�q<�(�w�}����<p�;��	o�C݆=�_=e�<�I0=�k2=���<?1��K<�<03\:<$����P�oI��w=��h=_�,����p���c��:�=�<�!'�[�<9���*4:f$�;I���vj,=��˻z8��S�ya�<�2#�u�N=燪�����"�;^$=2�)=�C=b�R�0�>=,�<O��<��7��j=�c��]$�< s����Q��lj=��=�=^k	����Ӷ���ؼ�},���_�|�W�Gx���(L��.=m8E����<���<f�緷~��_��A�<�؁<]]S=p�����t����M=�!K�[�A=���<��=.C��.#=B�Q���Y=y6��2鮼t�,<��<�[�<0�-x��OB�<���<�&�<��,����;�j�<6+=�����<4N�<�m<����%�9=�?����<�U=��sh���<^s<L�4<ˍ��|=g�q;/+��ݼll[=ߟ�<f�=KM=����z��<�4�;}���X���w���<�K=�?�\�=.����/=�M<�iG�s�M�WC��x�<]�<��3��@�<��=*��uX0;�#V��n^=�=������+t*<q7�{R��S�����<��'��"=@����44<�?<y��F5=%~.��I$<�l��^=�L���o<%Ǟ�аf=�	"��}= $<�r)����;ƚ�<0�;��<�>=I5C�2<��=
_<�Uv=U���~�=G�l<�A��s�-��zU�3+�8x���G��/=='j� <<B�������� �A� ���������������ƿ���[���|���;�w4<��=@w�R�=��=�����E���żB��D$=/�L<��<�rڼ_!<) �o)���<�� ���;1d<�,`�=�@=j�>=�A�T��˺]=�'�;������=M鈽@�����:`��<��`=UԻ�v�ȹ6<�g	=���)���i��n�3=��7=:J��<��;�=c=xf=��D�q���<H�< 1���lV��8@<(-'� �"�(Y��T�aI�<����U=�7R=<��9g��<��=���8�E<��v����<gS=d;�|�K=��=E�W������(��¼�Qh<RH-���!�'����KB=O�O�J�S=t�v��o��&E=4�޼�-=>=�g���=�a漞F�	<�F=����'J=t�<}�;�����:�:5��<[J�?5=��;*������6ح<u����D=���T!»��)=	h�<�&\=;ڼ��<Ț��3�Z=��]=�!�<ƀ�<q�F�qX4=�ȼ���<�E	�b�8�������#��G��B<�gM<�Y�<^����;�&[=���&��=-��Q�	=@L�<>�o�
<�v^;ܰN=C�)�(~R� ��� ���之z_<��A=�<�䡼��Ｋ4=D}����<ž~;�w���#�d��<��=}E\�\垼k]�<
�Q���F=�gټ��ҼX�;=���1�.=���<R��r�Ⱥ3��mXF=V)=.3�<��V�D9<��;\�9=[
H=IC/=7�x<tӣ�+�};d�	��:�֯;hU�;�)��AC��9���8�<B���[=ì�<$��������mG�:b3�;
�Ӽܲ��«<9�<H��<䌣<��<"�E=�$��#���=9��$�
�%�>=�B=�eK=?��<�n��vy=J�	=�� <�K=�񩼣��~�w��XO=���<&���Xx=�Dn=�$��^s|���Y;��<4��<�ZM=�j6<��2=�(�:��$=w <�lE�"=��<-3^�T�7���1=�Q�<,��<,c�0��<�0;IP��5�<^�5<��ؼ��a=�=sN�	K����J/Y=8�=I ٻ�6$9���<6H9=���=op=
,/<��=������<�h'=u�O�t�7=^��;U�=��9�=�[��0�{�y=�)2<�����=E�<=n͸�,4���>�6=pއ� �H��]v;����}�;��P.�;<�d���s;���;9o��XP=G;^<!V�Hƥ�Ar�?=dT�<#x޼2�.=���ʹu���7I�< O�<b�=�ػ<?�弉�=sy�R><�1J��n�<�J�<*wR���?=�L�<-b��o�6l=�LG�?��<�}��n�:�V�<�N=��-=9��;� �&!7<�%�<M�;��2���:=e���=S!��kU=��D;~��<�5U=Z�[<��Y�����b.=�a����<C�����<�b:=<�&=OjU��� �Z!��k��<š�;�2�;�S<C 8���j��Kw��N�<<֚��>=8�D�/�<9��<�Y/=�$j;��!��!$<o�3�S�g;nM5=
(2=)�j�!>h</��<��H<h�a<0g=�!=YrF<�z<�O^�T+O=7;���<y�
=X^�<��9=�ܼƘ`=:==#J����<,�<���WrQ�OH<�JB��H=�8q=G��;���4W!�t`z����wT�<]2��m|��DX�"r=Q���j=����O=]
= o ���	;ٽJ��<�޼K��<�Z<���Mi���<��ƼI��<��U��m)�I���4�<a>� �2=8�u�(����s<�O�<R{�9���<>f%�4o;��G�� <a��<�s�:嘫<�=(=O���i�.���=�Y��/z=�	<�\�=��)�J?C���=��K�=�T�<݄7<�$���;��<J�N�������}�i����<mߛ�d�<���<IIA�qi�`R=�弜@�;%`�h=(�o��+��K=�_T:k�=�$�4�#��<w.S=�爻g+�<�������=6���׌;�����cE<��ܼ�R&�YV�=��+<����$߼���"x���-=ټF��<��P�<5��ڔ��<5�==�v0�@�{����<.37�Jw���C�<󗯼�9=���:��
�o=Ȁ1=��<��"�+��<�����<�ߓ<X��<���T�=R�[�Bh=|@��M����K=�P=u��ۿF�߅�;4����_�<L|\=�����<�u ����,�[�=M/`�,}98���Z=6H�;-�<�����+��i��<��r�&�M��p�=�셼I�W;��ܻ����x<|��<��
�)P ��O:��_=�i�<��/<F�N=�����A��G�<�{G���r���I�ż�ʗ��<�c4=�p!=U �����S&6=�����%=E�@=�l�m���ɼ��8�I=�e
<��"<�c�ȁX��;�<�ϔ8�O-�&,4��������N��~o<��<`�K=b�U�����k������~H�J�?��� �b�P=�%�<��H=�.9�2�	����-�M�d�
�-���I�.9�<�ۘ���Ҽ	ɪ<w��<�;Y��#=S[=,��e������0�J=+O%��%@=hsU�U��鴼��<H�u��(��m=�����<]r�:Kh�S�r���i���=h�J=�O>��Y˼i������<���,�x�;C�)=�4=�;=��#=e=j���$��ա��&8�k]�����]=����<X_(��Q8�
eK<�һ�eċ����<'�P��؊��D=?��<�=\��J�����9��<�}B��D=��Q�#�H�2�k<S4=6�=p��<���;�9�}-��J�/��m��[�*������o<>��m�޼��;���W4���������?�=4��<��j�T\���'=]�(����<9�0=/^&�)rE<���<{_&=��f�=t���w�p3�<c��7e?=��
�9͖<n��:�s=���<�������_==����{�<v�"=�>>=�7�<F+�<�E���<��s=h�>�|l�<���N^�$�I�	 ;&�-�V9f������f�<��$<�ѥ<�t���?=|�<U_?�Jx-�O�$���L=�!>����9@��W�2��a��	f<�!=��y;f�k;6���Չ <<�ڼh�����<�M���X;<�<�<�1��0=v4ڼ�|-=݆Ӽ)C���c<~�B=�躛�<

���]=k���F���m�Ą8=�h0���@=p�I=��������<�e�L-	�{�=s�E�*7�T�һ|�R<y��u�%��<��^���/;f�C=f=a#���%�m�`��LZ���&=
�=m��K�м)�2�M�,�)
�.��<�1a<�;�*������gƼ��k�2�Q=�,�<�=��r����=�i���=�Ԁ=�B"=�$G=�_ü��Լ/�L�]�2=m-W��'�T!y=v�����R=�:5��*1=�����������d=9."=B�N<�r�;�Ws9-Č��.�L�9<��;�K�<�=�5;�/<úk �bR=��b��dl��v��^�{�țK���~9VEټ��Q<�Y��֠�<�+R=X=YA�<�G"<?a���G��:5�?zN�X�v�	~��M/��Y8=� Y��P
�1sۼ�c=+A=C�<k�<�'�<1�9���:k����0=��<Ⱥ=���<���<��F=�4<�L��*=�eK=jS�<���;^ =�F���l�=)+=>5��ļU/�(0G9.-ۼ�='��#=���@����%!=��v=��Q=@ =Ѝ;=g)t�		=*�K��AG=��n���<��ѻ/����p=!�<Yj�����z=*&��P�<=5<s+=�Q=��;q&�LA5<ڥ;{O��O61=t:��?&=�ˀ��L�i�<K&=e�!�jA޼��<�(��	l=d��I3=�yϻ��m;�����,�s�M<ׄ�;Zi=��u=9�<X�U;�P�<�7��_6=�2Y���7���U=n�_=��o�� �Ӊ��!y�;+��v�F=��q��Z�<���<���f/ =O@¼֔�<\逽�-���\=���9h�=E�伟��������;��=��	=�鮼=h�l(o�!��Xh�L=�<�j+9
�ܼ�_������%���;=�?w=��8=�]=�q<���_;:L�=�_"�����F����4=��=f�	=��A=Y��sqS<-W&<뼵���H��ё<���C�ը�<�[�:2A���R%=�+�0μ�	=A�<���czu<bd*=�d����=��;�H+���;ȃ���%'=�*���=��B�;)�\����g:Ql���6m��y��c`��c���Fp���<`�a��\.=���I#�:���:J�=^Ȝ<��<"�<�w=*B�:	�a��,��"�=t�=�RQ=�ŏ=��:Z��;H��<�0�{�h<���<�^Ӽj�����Bw��w�OVQ�L�d<`�1=Ø$�\ �<��=U*�;v��<(-&��_��e@8=�5�)�s�k{W=Zo�}@[��|8��w<�\==��ȼ*�>�񹉽r主��<�ݼC�ӻƔG��()���μ�V�<+8�=4�o��VE���<�=��j�,�ؼ N;``=<'�4=-��.@�<��]=&�?<�@���
=�ۅ<���'�)�2=/J!�0A��o5=�Jp=�����=����#7��;L==�_=�Ts:@��;]����-��s(��K+���:�#�<H���=�, �5y̼
'����<�]d�̘�<�Z<��<W��;��<����0=�腻y��<=�C��ǆ;��T��<H:^=K��[�t<�R���Ǫ��w�;�c�,�8���4<p�_=;���5�_�U�W�@e�<9]!��Q輞��϶��;�;0��+ɼ�)�	��<aѰ;(/m�G�=uj=�����a<� �����P<鼡�=��b=B�����<���;3�dР;�<�;i =:= ��4�=c=��<˼�"��ؼ��<i����矻i�n=�W��<�<��%�4K�<�T�<�&<� =�z}�u�ּtt,��P�<|:��Z� K(�6�<!��<Y%=���<��D�;��py���yN�4we��j=��2�\k��U�Q��]]���y=��R=<:���F�=#=pck�p�<h���<����<5S=L�/�TR]��0+;^A�<�!����������L��G=*M_�!Y��.U=efE�D�0��� ;�@=I�[=�#b=��&=�vl���=�=F�w��9�&=4�<[C�<���=�$Լ��i�;��G=[=ُ3�'Y7<��;y��;��<J�;�T�]=����)���2导��M=��`�+�U9�Xn��!�¸�<�	��Q����C��Ă=���;;�}��D�<�j<��p=]鼀84=idV��`9��h��͈"���;!!D���C�2=7!��3!�9�7�'#&=vud<�T�\�d�I���������=j��[�Z��ZR��&�<�8=s]�<���;��N<�4]=��3=8K�"��<7�V���ݼ�>�<kZ�<|=��b�#�_�pRv=?��3?�����q�<b��<M�F=���Q�<=$W�����{g<�����(��v=��4�K�V�E=Ą=�^��jg���J=�J�:<:�c��:��<��˼_0���E@=� =6�a��&=�}I����+R�F�<�̼��<I<A�]=����v=wr缺�5�r�"=�׼�f���+�3J��h+�N ?<�r�&�=�K�3������;�Im��~_�K�t<�hi=e�N��l�<��:��,!=wڼ[����k=d+c����;d��;l�l=��<Q��1)C��<�6=�/��x����R�gY�<�ֱ�Ze<��[��),=9<żM�;���[ei= "=���0wA<������q�	-�I��S_��1��Cb�JmU=#u�!H =<�����=�����~j�VK�<�f�@ =?��:A7��k���-|=6�<lt<��޼��;����(�]��)�_=��˼�X'�t�C=�F�<ˮ;F���)
9���Q��� �X3�� 6�;`L<Ϥ�<�J#=1;�<�?+=j���=p�=l"�;uAc��t;�^;��E�����=�)�&j�<�F�;��U�:F�8�j=�=��0�j�=vl'�-�w��?T=��<�A"=��<�� ��j'=b�!=�S7=�7=��B�d7�=�	c�,s`��-�<$��bźs�)���;<�oF=����%��K�<^���r1�88-<�iüCF=��;<�CI���B=N���=<ʣ%�_󅼘���{=�� ��W�.�}�]U��;Q�o6�w�Ļ��=�a
�\>�U���s%<�'���<�Q����/h�:�lV<�);�xq���^��g�;2`N=c�b=@�<L�1��J�X�a���Q�V�7�8=m <f�.�H�"� �H=����h��i���ɛ<�&���%=���!�=.�:��<�(�;�w$�����E ,�N�߼A<�M�<�M@�Y�<�M=b�� �<�kB�{��<��%�!^�ؾ+=�<}��;�=�}=��!�͞9������X?=�|�� ^�g�l�3��:^����<L�@=B��;9����ԉ<Զ���R�<\�=��=�4�`�s#D<����e<�n�=�~��+=^�?<b�S<���<ixj<��x=-g��"z7=_�"��e�<�F=_n_�?����;	��<��-���ݼ�@Q<�"i=�%������<�OM����<�o=--ҼC+S=>�<b�<��S<o�:��H��u�"=����l<�m»��=4
r�v[���+�P�o��ۈ<�����!���
��*�9ʰG��c�;.0�Ev�N��Գ�< c޼��=;K��.��oܼe�<���Cx�;�y-=���.�`�ض���Xd=�=�@ ��2��	�e<�o���i��H'��[ ��Y1�*e�(]<=���<�xD=�-��\��_s�;b%ϻ���LM�;��=�;=�x.�5UK<bˤ;e��u���o?N�}xڼ��ɻ��3<p��9�?=��<(7a=�^�������[�#-J� �^< K��p�<a?8���<_�#=ґ;��U=Q�g���%��l��
��LZ'�pQ�X��=���J�b�򘉼�F�_w�<�V�:�yg<ջj�3�V<�C�<�6=�%���:��X�T<��=�H%=����`�~=;,#=��*<����;������
�hQ��?@�7���˭<��%����x���_W=L=<�!�<�h����n��;:=�"=S�<��H�w�
=�F=$�<��{;�.���G=�$<ʜ��3jD=��<��C�+��t0O��[��U��TV�7���-��#.�i8=�"=�м`�޺��'=|�ݼD�?<"o�5E%=�RS=�d������N�����<Z=�L <� =�$"=��4�fD=�~��Y�z,�<�<�����+F=�{�;��X=u�>���:=��]��9��S�;�T� Z��HB<������=�����f�T[?�����;x��JE=��9:�b�&���z;<UEO=�QT=GZ���;��0=�	~=����oI�'��<]<.=�����g=��<��n�#2B���|d4���;��¼S�K=�*F����<3�8���l�<j�2=A��%q�;��W���S���9<hp<� ���*=���<֏�<�I�"�=���<��<�)=�:�r�G<�Թ���W<C����=�߈<=J�1�_=�i�<Y}�<(�=˨=n>���I<�^=7����=����=ᎇ�Gb�ݳ漮�y�]��<�%�;:U!��6:��A=�	g<����¼J�N=���<��L="Y�:��h��b=��<���;Cļ����g<S��<C���Rb�X�r�I���/=��]��i=�u�~%3���ּ�K3=��κ���<1[I=4��< �!����8��%[�<�+�D�.�o��p�8��}W=;8�;Tb=��<)�!=��
���<�<��B=zO�sjӼ�#?=�������Ҽ�qi=W~ֻ��=����:d�b�<����_��_��<n`z��O������:�'�<��:=~S5=�\�<��"=�!�pg��<��$��Z�����&���w�4/=.��cK��J=�U�,2�T�=���==<\�<��w₺�fм��N� (���U�<0���ͧ�=�g�|I��Z�<e���= ��������<��"<3��<��鼨�w�̟��D=� =�R)�Q�=��Q��\��=�uI�7�E��0;��Y�^�<��H�r��;��<fS¼*����q����8۵&�� �<���$��H��<����Av:��s=��Ӽ�C"��[V=!N<�=�[=S|7=jM�:�c�����?a<��}<����W=�_<,��<����q�-�q����;g����R<�'������=�B<�,���u��=����C:6��"N�F�3=fׁ<^�=�ZP;DaF;[`�<���'�T����<\2��ZUy��G��Q=M�R=��:Z�
<����in=�� =}�8=��<!j�#Kf��3м��0���=���}�0�=Ҍ����:�D�`��<l^;���=&���Of�+i�T�<��j����o.;_���5���1�k==���b�<P���M��qk<�)&=;�<����i=w�c��,�<Ӏ�<*�*=�}-=؆�<X�/��c=K�м�;\�1�,����>����<�z=�/L=G���3<d0�mu�����:C=X-�<��<Q˯;8��:xxܼa�u�	�i�R�<�== Y'�WS��-�<��]�2�����8<=(�$j=�F&=�li�=-=u���a;��*=��f<h�=�C<��/=��J�[0���<D�<�8�_�O��3=?>��d;�aT�C�y<h�:�!H��X[=N����<��9:��U���]�4�P_w�ME#=��r�L�6����<��S<\��k�=�]��P=�Q�pF�<0Fd=SR[=�*g�I�����;d
�<�4��=���=q���lx<�����=�u<�Z���=7� =+>�<eI-=)Þ�8E���J�<�_<��=��k���O�*�X�M�O�Q�,�-͉����<�T2�5�<�0�_r缛M*�`n����h�77L�3<�4ƴ<2D��s>[<f�=��d=yt�<w�&<`��<t=�:�)T���||=���<�h=�=�8=�����Ļ\��=Zjü�~��V�*;�<�iaa�+�"��sJ=t>=��=���>� ����<X�ּ�^��w�9=rUp�9=z w����S>���<�M5�
4=�[�N^O<��
<VuI=d��<�t���.=h:�c�H���/<(ƻ���=�'��L�<t�J 0��s�<���<����<�9W=�T��Q=��;��?=�E=�\]=��Y��y1�r�׺��x���F;ڐ%<��-�Ux���S����L�� ̼�'�hю<��~=Iz"������)=���<p�<=�\�=P'E��!�u�<�ّ<�q�գ���r�=E��X�+=(Pr<��&=�H�<�k�<�o^���ϼ�0�;���:�)�.�ƻZ�$��	��7��~=��=G����|κ� 9���m�c���
=�G�����$ǧ;���<���<ф�;ʄn=�`.�{�,=;λ-�7=�����<�/���y<��;hg�;������;��� =����>�<��I��^h=.�$�^Q�$�f�G�p����a�5��.O=�W�:�|v�Z\���m�<��<o;��D=κ2=e>�
,��;!�!�^��}��`g��9�s{<�ph{���;� $��B =�8���P=M��;�e��MEP<�����弙T=�3<]�<�����0�67<�� �'z=�:���jI��t$=��ӼY=���]Uu�ΰ�<!��K+=C=�	1<�|����<D<!;C]*=A1=^a<=��f��/�JZ�<�Ia�#i�;��:��@=;�.��=4�I={O=L7��W=��=S�����>�ƪ�;�#4;�q��i�<��Y<�u\�ړ�<j�g='!�/�;�nTj=�J@�Z�6���\���=%=��h��=���E =ǁ^=�[�Z�E�
�<8g<+�d=e��<͸l���<jF;��?=P^���F��м��缋H�:S��<H��@�$=fo��Ƽ;v�<O�=�F0��8=�{u��P���=��<�
'=F����4C=���<�a�|�3=�K�<�I���;�N���j����;86�wR�<����z�<������<��HS��.���Z:�x���<b��<����ʣ;��ؼ�_^:1�޻$=D�<;��M��;`��m���O���f����<�˴�'�h�� �T?�5D&=]��+�_�IU�`x�<���<I�O=1@=9�I=2� =�m�<_�	�WD��T4@=t����Z=Ϛ=�#���'<��b�f�<���<h��j[���v<h��<L�<&���-ּjn�<���:��;j�ֻ��V=Tn=풼9����A� �~�D=Sd�;7(��p�4�x��;W�7=L9�Q�D���
���<z(�<�~�0��<�Ƕ<�5�< ���X�<2�˺��<ڮ�=+'�<Y�<�	=��Լ�����C<��j<P�D=�k����L�ЄN=�=��<~˃<{ɻ����P<-�"=�ƨ�OX�<�==I���R�v̪<u�?=qb�;P1=��,|=��=p�l<Z�a��A=ɵc��S���n�w+P�_/��7T=}��<�Rмʤ̼U�A���x=(�!��e2�2�i=p����'=��<=H�%;��<KQ=��e=Nb��Ż)=<�g= �|=�D�<:��<��=���<�F�<�j�x�%�w�;�1�;�t=���<��;�d=ZjＮ�%�]��%��UF<88����;O,y��}�jۼW<��-C�;�;S�����b��Γ�;N��\j��o뼉�<��q�QiI=��r�#t|�+��W�8<G���MJ<٥���
Y=��E;��!��!�<4s=��D=H&��k<���pl'�:�ɻT�<���<�0=����N�:Ȓ<KT��U5w�= �ӆ����=Bp=;��� �<�>?<�$�.K;<枬���<;i��N4�wx�<I@#=Ѫ��+��<�2�:��<�7�f��<�������x�=�
�<�]�&tڼ�J�=$(�2e+=^��<���6.={�u=�y���5���#�����R�<�h�<�������Z=X�=��p<�/<lx��=�p#���<��<r��o�*=A$*=�:�i�W=�!E=������N��
=N���|Z�..��e#�㾼b{.�H�<&=7q���;E���=�E=|=-k���3=^��ypO=i�;	�s�E�Iqa��H�;�Z�A��<��8=d���6=�e���.���S���>=�\$=07;�ν�;�Hu�U�}=���;&B�<�*L=#r3=��O��M��e4=�s;"�����:����z�<A}=��l�<'2=:�>����濼Cj�=���t���=�ǻ��=�Ӈ6�k���࠼	@�;�ԻY��<�{=O�<Wd;<OS
��\�U�� ��;�2�<�-o�:�m�a����t<:�
�F���Ba$�s혻C�==�)���.����<ɇ�<�<8I�vƼ:7=��<o�I��3v<
��<r� =�R༭' =Hz�����<�ɼߦ<��-=��Z=�Er�Qb�<��9=�}7;q�"=R�=�".����I��=ںB=A��<��<T�2��4�Z_U����<����#;��-=e	�O��<�]m��.�<S�F��'l���<
�`�;Ƥ��(�<�f�R�����=�{=�=���<o	���?��Zx���_=�<���+��U��<��?��O)=�����o���[ <�*���=�I7��?=���<<�<w5Y��+=:G;)��A�U�_��<y1m�sK�<�+�<�И<@��;Tǀ���&����<]����h=�X׼�����߼�$�;�e��=��C+�< ����c(=F���`@�<6f��!����4�B<�<*;l=o��5k*�4EU=m�<��<�*H�j� =�0 =��W=r��e-=��S����<͵< �k���<�����<T�?=�^=�b�ǀ��C�,HY:��<�\�<J���#<�^=-U�����d�ߖ��ao=��Y={�6=�g�<O:6;xᨹ���<��W;�rR=n!��)���rؼ�V��'����<v��.�=����v<�[T��?_=A�<��y;Ӱ�<����pP��a'�+[�<���Ώ,�/�����<&:�lK�;b��(^���y<~��<�!w��S�<;�c�<U�d=Q�a���%���a�b=g؍��=���Ҽ%�w�UN�<�&����\=�^���.�����2�L<�
:�k���@p�g�T=�=��6����񜁼�=�<�?��dh�g�P=�)���q�LA=%�<���;��6��7���`��1�<w
ۻ���<��C=�P(�\�&�"��=��O<͝r=�~�,����:z�7��5;A�'=�F��݈ =��W;'��G�N=@ �<�R���ZD���,=�b=��QL>=Z/�`w�k�}<@k˼�ú��<+V���+�[F]<O<
�:?�<�,�<;���8u�仁<����\=��3���<��-=�Cq�+Z=D��$��v�2�<y}"=��*=��<U�l�i�T=������G� t��,���<=�0`��[3�x�<� ������8��<�b����=����Z�:m=��ݼ.Y���ߥ<�|(����;Z�$=7lt�4�<���;�Z=�
�l���r�S=�X=�-=\/�i]=%S�K�s��A��}Ѻ`t���<z�F�V=Q���l=BN%=D=эk���;-��M{<�f��Ѵ���c<��Y=G������F�@��2����>�؂�<0pl�<���<KfQ=�ʋ<Jd=U��]�n��1�m:o=2�� �]�4�!=5��5��0Տ;E:L�Ii	<��<��4=�6��_�<p�K�\(J��r��`�=?7�=Jo��·��	H���T�]�<9���=�D=�=�#B���<�n;����<،`��(�i_I=�J=O��9��7�p)�g,x���}�Ҝ�:�,=�}ļ�D=�W'�L�-;N�j<�N�<z	����ʬ*=O)/=v-x���T=��4�nD!���<6�e�c�,=F�E=�9=xf�Yn�U^[<���^�<&�?���;��"��L��;�Q<�J���l;+z��s2=#z�8�<��,<��o�e�7=aVe<�:	����#=��޼IW�<a��;ɗE=�'9��q=����&��[#<�S��<W=��n�b���HӼ��Z�`�=�`=K�;�ؼm;�tZ�[��>����k�o��<�Q<��=<i;�<(�=�������H���_���P=�s��sN =�>��m	;�fF=�֭�by;c��)7\��л�EѼ	l����j��6S�cRD=}u��� {;{�U=�<���o>*<)�+������s=�k�;!d�����'/=���c	��|�D<��G���<��<4}=��^=.��D�k;�;����t����%:��<RS=	Z��[ <�E='
< =>#C= P��5��A=@!���G����*Ӽ^�$�*���q=U�<�g�<$\�I!�<>Y���=N|�ܼ鼑q�<�<F���$�/=��<��=��;y��<�4��*=^1A<C1�i������-�<e�Q<��X=BW,<���<�ho=NO2=��<;=�ň�I� =?�0<(�;��<�S���Z�)g��+��״l;��c=Ω�<�FQ��������<�k��6t���L=�T�<��<��<#`�L�ļ�A�<i*���`<��O��d#�܈D</��+�8�0����I�;Y��fc �HC=�G1<����q��Ĵ���=v����TP���h<M�˼���x�U��<砘<��0��L9=iY��{v�;��ܼ �����w���{<[�Z<o��v'=	C9=�I!=�</<:��<B�o=�����~�Nbo�h�^��#�+Yu�]��O㹼 J=���v:<��,<�&q=�Ƨ����<b�!���(=���<�9�<M>�<�uR�H��;�""���=���<fڼ�р=�y=�s���s���,�<�gS��p�Xq-��EL�	�����	Ve� C�E9��-�-=�w��&�8=@p�<�.�<R��<�l=��p<�F�;����70i=��'���<���;K���L�,<��r=tU=8
==�����<5�H=Ȕ<��;�y҈<���O����+�����Y>�t�<-S[�;wH=�M)�MI<���C�=.;:�X耽�1���H�=���Ze��� ��:=ɀ�:�e;��<�n��#C�����'Y-<���<��=����<�^a=�d< �<����`<�O-�<"�\���H=�vZ;�aҼMB�;p��XEU=e��;���`�2�Ӽ�2���<i/*=�*�;J:;;�z���-��\K7=[u=�"N�Pl���-���2=���<�H���b=�]X=�X�<&A�����T��T��O\�4m<f����x<-l<����g8A�N�<�_�<������:=DOp=x��<I����.��6=�h��-����ͻ��N=�0��C�;�;��]=f(Ѽ��<!����o=w����M��Ċ <=b�U�=��=�l=�V�=�Z��[������X�@%��j|��6�<<YB;�A=���:������"=�+j<��'=�^�N�T�i�����;bD�<��S�<]�μ�м��Ϥ��j<�x��zN<�u���M=I[ֺgYj=U�=p ��ޑ;�z�<7�R��-=&i���=��O;��R<&��;
j���1<PF�^�1��j�-�N=��o=�z�<�޼�K��r=�N��>�h��	�?=�7�`��<b砺��
��B�r�H��>=Y�g�2��U=X	�<ǲK�4�=Sļ�r*�,�<TE=��Y=Y9���5�;�W��\�U�=_��=Lļ2̴<�WA=/�<=.�=h���|}/��PG�cc�;&PT���9��,���:}vż�<��5�� �<�'9=�L��M�= �=
x�<'��w}����=.�A=J6�/3;��<�|O=e`Z=B=�C=�R<:���ܼ��K=��O�ǣA;�v9=�n=Q=�['=�W�<s^=t���pC�<d��<e�O=�S�<= �� =;��<a?��%	:���&x�;�
=6�����<���=� M;��'�vn��[�����<�n;��So=���=&��8�ż�a�<Ư_<�B(�^<��E��W=�Sg=,� = gf�F����=s~T�_�<��n��1L=��
=�J7=pc�<29�;@�D=��i=;��<U��<=x�<Rg=��
�r�A=��<~\���[��(�x�;='VO<�	��I�4��
=�Z�V{v=�
��o���ޏؼi��<i#����s�=��+=�%g��(�<_��+�~=la��j�s=�S=T�<~��<�8��j���!��eK�WW9��\�<�ִ���������%"=��<�^)�؃�<+��l��<�/=<z�;��o�Mw̼-�.=�fI�~aq����<�{X����;�d׻I��<�L-= nM��ٌ̼:�y�-=A�O�G�d���;9�=�=9��<��v�<D8=��N���y���<�:��i*����<]=�y�<Y���;R��m�� �ʻa��ݷ=�ǳ�P�v�����'=��k;�6=��^�j?��$��,��'�;Yo3��ρ<�$D����<�",�� �⇼��e<�J��ca=�RD��~�<��= 4d;?4<�uG���/;�z�<l�&�x��<�hH���\=�!_��\��X=�]=�P@���5=qJ�<L� ������K�T�Q�P�O	�;a��<{ڮ�V���K��@tY��ŵ<Ha�O��<Vo%���<8T��ÕY=�"\=�'��u�~��4@<�;����)=�_�=�$~= d��w�u=�H=�;����/�̓�@< =���ı<5��:צ_=���;���_�0=f��ջ}���7،��bl<���{E�:+<������c��<B���=v:<�g=_�vr�<Z]I����<F7��I5=�kf��eػq<YX@�:���p����<m��ش����	=�"d�Ղ�8�L���+d=Dh%���<={ =md�<�<�f=)�;v/N��^�]bh=��=Y��'�<1m3���<Ǆ�<s���I���ͼ�s���Bw�<�=mVa��N=��F<�h��9=��ͼ�����=S3(��c�佹�F<��F"����<�p1�toY<�5�5]:� �T=�=gK-=�C�, 3���	=�^r<���K����<���;r2�@�q�~.�.�i�/ ='�(=�a�<K�<�={g�=�ԍ;�SȺ9=x�X=i��<�<7汻J���{$=��$=�I�u�����<y^�=� ;*��<	��;B�5��ڝ<<�=���<T��Y�����ż��?���+�:�!���<�|<��'��=��hF;��μU�׼�1<6����<�~�;�=�}ٻWHV�u1�<'�<�Q�<��4����j��ث<�=3v�*����7�؄�<�9&<Z�~�U!��u�=:��<� �=T~��Lm����Ub�te =#˻*�c��i����;���$�Z��=�s%=E�;��l��
G��eǻ��1=�:��F�g<
�C=�&=\� ��G��<2=:[��g=�	�;��EZ<3%N="=$���=�8Q=K�̼s�=k9̻�x8=0��ei=xhV<�5����v��H<鹇<�aU��ʋ���@���=	��<�$F�ks#��K<�u�<�7�<����9�<Bg==<ܫ���_=4�<�2�<�
=��,<��]=�]�Z�z��h�J= ©���=�����H�=�F���(�<�x=�<r=(1ż�x�;� <أ�;/I��v͟�4��<��<]��<�N�<v�%��<k7�<a�C��C��n��!=I=|�QK�'��<U&=r�
=D�M��U�<�)�:5G�<�m;�Q=��;e+=�d��R"������^�<��%�F+�<r�뼏�?�js��:�[=o�=�9(<�d�����<���V=D�<q�<�ҽ����<z��[�=/�i=�f,�a�d:�ok<�W.=����|�
;��<��K�� e6��;*�Dh=l�<R�<����@�ͻ�2h����Hp9<ɕ+<$�)=�&u=+�4���c=��-�(Q�<��X��+�?&���-G=�?�9��<�_�_F��K
��żL����=.7c�0t���<��2�<��3��mn=LP==�M<x��kܭ��EI<k}A���f��	=�<Q=�=�02��ٜ����<k��b.c�L��¯<u�.�!Z���|S�(�y�<"�<XN��|����nl�ʓ�<��m�D'l=q^���=(�=�O��f�:��6���+���<��Yea���B=s�;> }�>]��ˢ[���T=�Mi�w?j�+�=0�h�o������w#�k���6t ��,#=,�;�S7��b=�		�^�W=;�:y[�Q6���<��桼s3�l�<�"3�m1,�kf+��6�<�<������b=6�<K&=�7=������˼&Ó<{�<��,�E��@�+�M���i<��<�_<� �ڃǼ!�=����=	�<�Ä��c<�������N��<h�<|�0�l'-=�:?�H��e<�.<�]C=댷<D%�<W=�Ǽ��=C<ټV�Y=;�&=��F=��c=�x���[��qR��S�<�F�&<c%b��'�<���<���=�3D���:��9=ɼ�W@�z�`= VQ=.]B��?�si<GA�������׼�b�;�m=a[(=$��<p�}�/z=��Fg�<@Zv=�٨;<?���ŏ<�ɼ,=_�=�����G��z6�<�6�<���]+�<�==<�����Z�u�=�|\���==k�v��1������|�6i<����e�<�o;ו=A>}��S�L!<�m��ټ�Er�s5l=��_��V��������;��.=��]=�=�r�-����L�:L�_�'0�	�<�w��b��:�;�b@�E�<�ә���C=�j;�I(=��<�J<Ax=S�b�k[C�s�r����;�R	����t��`K�y���פ<�q��p��GQ�J?#��f;T�ּn�%��0R<L���%���b=�X�gP�<��O<�W
=Vyټ�#<sT��6�;Y�=�?�<7��<�nC=���p򼸊I=l��^�AO*=��<��
=��<Ë�<�����~��<tG��\��P`=��j��j��8a�׸D=衼_&i=�W~����<כ�<���<;�N�eb+=��<>z�<ѩ�������+�F�LR=?�=`mR;�<A�6=�%�>�I=Er5<;@�<��;��mԯ<i h���<��N=0ؼ�a=��W�cHQ���*����;��A=1�z���G��7��Kd<I��:Lo.=�
!=S�A���=M�e?����<�:A�+��;^�M=w�E�������s<�4��%�<?�ټ�V_�;���O�
=,=�5����;n��<��=v��Bz�l윻u�"���<-���~;ߎ1���N=���<��?<D� ��;=�.���< d����8��=�Aؼ���<d{����=8���*l��>=��;��=�V�;��M�4V[<��X��QS��<-Y=�6��rS;��M=��W�-���#�;`���7�)���r=��I=�Z<�闼��V�n�<ʞ==#�A��"� �=���;ё!�:�+<Cq�<\E=^�Ƽ��ټu��1��<n?;�L�<�0�<���<�R��V�a�$��Q�<5����a=)'����<l��<�{=��0�WU=Ty�� Ja=�
��Y,�z��~��B��S�u��7���������-=�"�c�Y�p�z!$=hI����Ǽ��=�*=B�}=�i��x5�<��=9�N���<��L<���L�3+�;�2��x��<ߟ���8�?K!=ʀE<:��ܼ	r�f[�+�=��4=��m��P�k�k8�k�I�,�=����$Q=�=U=Y���8�c<J�����KfV�d�<Ni_=m�`<&��!Җ<�x�</Gм�e��鵼��C�\�S<�����A�;�<=�JM<���;��9�����9a=!��t*��OB=$��;�-A��%=4(���b�;�Z;�E��<�ܼQ-��q��Z��C���1�#�<��I=fH�<F�<��T��o�<��^=�����= =.=0�^=����/Q���2��D�jo4������=K]q<[����K��g=[�;��5= ����d����g��"!��ⶼ�|�<�M�W:o���ۼv�,���t������̼��=�W=Yt*<��"�R�<�M$:a=i�2=3�;1�&=���<�G��nL���<R=c�B<:�1<u]0�%�1;ۼ8�@0<�������m�
�$=��)�h=T��8���_==f�i=!�>�������<��*=\p�[#f=\�z;��=��= �1;��E=-9������z��m�JHI=!��<�X�r`o���	�\A7��gn=�-=�3=��6b�<Y�м�y�=f=��<����%�=�
A<*�&�lp��˼�
=w�;9I���� =�V�b�&=�:v�7e������f=\`�<oS﹧��:-�I�қ$=,�i�1�u[v=��%�`X<=I|�e7=�]=1<�)V=8�0=!�A�.�;�9i=b4=OF��&`�3w9=�<�,3=�h=�G���<�F`=�N���;O=�R�<0���M�-��Z��;.=��-=�?A=���>9=󉽼!	�9�oH���"�����Aj=8�A=�H�<�<	�9������t@�B�#�&��yV<�8{�o[��a�<�Ғ�<��'=�o,���ܼ6}d��%��)\���'�9��2O/=����P=5�<�a���d=d�==�C�<���<���A���^�Lг<Z]&�cj=�y�=2�8��;!Ѝ=�z�<d<#��6�k=�;���*��
= (C��W,<9������<�<�hy=$�==�V=�� ;�N�<��J=�DG��cX�Kci=��<F�k<�9`=T�;0/+=�x<�s�7؛;���:XɊ<�//=�ī<B��}<�=� ��,Ѧ�O=論�\����+�������
��=<��a��$<9�@��%@=8��;g~>��
�<�N=X�W���(���%|==
ɼO�2<�W�;H���:��tJ=j�;��< R׻]B!=���1f���<�0ڈ���vx�
��� �<��B��f=:Q�=l��EM<�_.�Ȯe��dR=7�A=_�<�$�<jjv<D�;��a0='л�/=��<�F�<��*;����`�;�#����=�R=��W�.~�<�PU��-}�3�	�Ԍ<�R�;�<�o7=U4��Z��h���t�< H=���S���=v��E3U�?�<v=(�Ҽlu=6�9���%�H-=����Q���l��,�7x�<�HD������;�8Q�<P�}��Jo �I�;��;�$=W�j=����R=/������u�=qH��ߌ�<u�n�3=H�!�ϕ=��m;���y��<+K(;��gʖ��S�N�:��<��%=>�<۩'�<�;�޼ӻ�K=h��<���O�*��-�<3���4ӻ
k#=P/I=�9�;�3<�ݙ<=�=a:�<�Yr�z���'��/v���:�M�=��=�h�<�]G:�K��#/=��7=2�H=���fh�4���9=��2=�> =_xڼ[ʼM��<q�<QS�:�B`�"*�ݞ���f��g9;��^�
=K㼒�!�R^5=*wQ=�X�Ua=��<c_=W�P=;v�=�҂�%�y�ӻ��ܑ<G	�S��3�</!b=��<��q=A��<�R�l�鼦U=��9���=&Ӻ<���9u��<�܍��k<=|'=�;)�!9=7w��L���G.<�g!=�� ���=������;�$J<��<���]l?��W��ռ$K�����e=�����A�J�׻\�<ԭ1=q���_\'��_c���ԼZr�x�;?���=�=J=���=��":TEB=��B<���<�l= �]���&��NX�#Q�7f���3�F�h�8�)�=@Ã���=����<J���=�� m=,��%Ob�.�$=�	=�*���{=ꑼW�F=��&=�Q
�4x=�ne=�̓��E�2M���ּ7:��C��<3�<�=P��;��?=E#�<�ϼ:{(=�T�W6<� ��<���<n+_= =dBQ<g+R�V%$=��P�47��=���m��M<?2U=�>��Z���<��K=��@=�b��縼�tB=�'�<X#��k�	<�gɻ���;�Y�<�9�;�3=9)`=.q>�4y<س:J�2�~�"���<ViB=P��;���cNK=9�k=�j=S{��<t2�vr�<�c�,��\;�}% �G���W�A2=��!=�hݼs�`=�0�Zc��Y�(=*6
=�`��_��J=�S���|����<��N=yk�;3e=�T����Y;ck<������+=���<�D�<�݆<��0=Zs�S7^;vmʼW�<@�ü���<yZ�;�(�<����4�6;��&�*���[<�����F�<(^K=Ƒ@=�7k=q��9֌�;��#s<�Ӈ�d�7�ȅ=��%<G������� =u���8�@���़~�t�n������u
=��S=7&��Y�2�D��;����F'�	A<7º<�N���z�<�=|��6J��,8=�Ni=U�aM$=���r6�<^&<�.Y��C��i5=U�<�_h�zT�<;��ZE1=-�=�<y�(=�H ���D=N;C=��=�Dl=c����s��E1<�e�ּ�m���o�h	�<�F�ן<�<=�
�<;��h�^�F[�󾇽	tK<4�<�
�c���y<����K�;==��<�tE<>t=�w8�f~���iG=�=v1Y���N<@9R<i�ۻ����t<��g��9���T��<��-�=�/��+�N;�<��4���>�KlV<�7y��q�<� �'<�V*=o~=�޼غ�<�^`��oV���V<P���-�<� �Fv�<�<�6<=� =�ơ�<$�,�G<��B=^���r��b[=�=ҡ�< �q�❎���<�{&���
��HW����<t�d��H�n':�o1
� 2��d=v:=<x�<J��P�d<Z�S��������'=lJ:=��=��!<V��<:W7�ұ�;����>��jR<��==���<��= )=*f@�3'�7��=��"	'����C/=�L&<�Z_=T��=1�߼{|Z=in9=�K��]�Ӽ�p���t��͒<��e<u�Ҽ��C;Rm�=o�ʼ�Y;���d�eq��{�<�\c<!n�;�e
�A�a<y��2S*=��������j<ޞ�<޺e�RX�Z�［Gb=	�\=|�F=EI��H��1=�9<��;/�e:X�:=���wM=�\Ǽg?�<�]r:F|@=j�b;@=Cݦ<5����<�I=v�<��`�Lp��]�z���3=�-�O-��f�M���t"=X���S,�P�=�C;m2=פ;�	����	=���;1L���g�<�⠻��(��=��@��5=�7r<�H��8%�<�h���#f����z5=c�;Z�@=����� ͻ͒���T��}�:�1�<w��E%=xme=Gv�� �~�j���1=͸b<	��<a^ǻ��"<I�+{<�ZB=&�μӓ�e8^���N���<H:<@���x=c9��ǧ: |<Y�<M��<��=�<n�8��sO�ؘq��O��=goW����d�l��8 �ƿ��_/��=N=��u����<� ���$=e�:=Y�4�Ev��F2�<'&y=�=0�|<��x��Z�<�.=�H�H=@/����5g���X
��k��M���L»cKW�&$�m��<X�<=[N*���Y<��(��H:d�=vf�<�мS�|;_w(���P��}C=5�ʼ��V=�˨<��@;|!-��A=��M_�������5e���=�F=0R�;/^�=��<�gaa<I���*��<��#=p�l=�DP�9��-�;՚=n��T+����;�j�;�=��;�-)��K��:�<4����}��*�C*v�xk<�c=�c<q�=�Q�e+U���<P����~=y�<_Y޼�����g=��L<W<�W<�2B=-Z�%BF�Ơ߼��=,��9�P�����R~ǻ�J޼�J<>��~�<��n���<%YU��_=@�%���<>zM=&��<4]<ЂF=���<RH=��2= 6�:3�����FE��;�=ű^=��=�^�;K���?n;�1F<�u={�h��=�W@=a<V�1<��H��]=:��:r��=�F���~<*l�<�@0��=�W��_��!�<���*0�l�H�q	=���<+�,�I�4=�wv=@�2=�g,�se��};�8	ۼ��&�&��NE��=�;_h<eG=��X=���:�wb���<�R��<�������<ٝ[<5T~<V<D|&�"'�<�rC���E=T�A<+�=�Z�<J1��~��<���=<�Q�7���D
=(û��,:f����=�ڑ����B�r�v��Xc�M�<,3=�d�=E�<�^<]���<l7=q�<s�"��J׻�qм69��; �Cl0��;�8�<�V4�S����IC=��#���l;�o缂�H�E��<\�_=��#=�8���d�=����û��O=�4=E�=Q�m=l��<T=�'��k=�o=��;;�=� =p�2='�7|�<��ѻ�ɻ0Q&�UX��^�)=�5�<�M���,�;�|�<�g�Flɼ�!�<P �t�K:�$�#�g�TW=q��<�`�{A�;0�¼p��e�3=_\<�'�7�Ѽ;}��1����[�bBj����r�}�8H=5����<a߃��>��/L�|�
=TW�;�����c�O�:=Pz�<�c��#\�)m�<O�ż�s�U�Ϛu=gǻK�i<���<_r�<o'�;�G_=���Y6=Rq-=}3A=��3�\�~=�8c�xr������㖎;��#�T���yɼ�=�� �dŊ�
ky���;r�w=KF��FN��ʬ�SL~�&r>�¶�h�<2�"<޵��:	�Dk(=,�R=�K=F =�=�ۍ��}�;�����Fj=����ץ<E
�8B��$�<K��<VA6��lv=L.�<���p�3��1������ś)=/;�{u��H�<�d=��+��u��ǉ�<�#G<V�ּ���<0�꼫`���p�t�>�w,��=�<�<=��<1�� H=��\<��9=f��<�U
=�S3=�M{�����I<�2���6�&=4�y��/8��f�#�)<S�=-�&��<=�Nw���(�/�u;�)@���<=�Y=���<<�:sź�5=t��*F���a���=��O=f��<$���&-<��=�;=�7��l������v2�x��<i[=0��<m�F��o=O"�K�8��hK=뱋=�R����,�<;�=�N#�:Ԙ;��]<�+�� ��2漑���2r�A1r=@�s=v�':C�O�C��5?=��v<)�ż:�=�Ǉ=�`�ߡ�3�<���Q��;"�=!I��t���h�u����<3�O��>�<xc)=�UY�Xp�<]^��ŀ< �=�r������ -== �q,�����<�M<��b���s<p-�;6�@=��8<��#=�K<� �qz<���[
�<,oz<��;��):a]�<�,K=S0�<�Zi���ɼ��f<@��<��;�J�<��;�R0�֑5��_<=ߺ=�۹�P���=��O=d� =7��;��=M	�;�.=v =8�.<{`����=h:�&ڞ<.�=*���o�P%���P=�G�;zۼ�/��UQP=�X�����<���$/��;=_�=5��<M��;h��l���9�<������<+bp=r�S=���<�gm<�}O����<��	�u�����r>(�l��;I��<񒆼_��;v��4�h�0�<�v+=g�i<V\�<��=eQ����z�>���v��%=�ˬ�џ1=։ؼ�4м#g*=�9�:�Ma�H�n���ܼ�M5�����w"�<
��0�,��é�13	=���<�Թ��{�;l|��e���H�}YD�B���r�
� �����C=�$=�x���=:ǧ<R���i������:z =t�
=�\�0\< g*=��U^U=�0����<��<��!�h��<6��+�G�����a��k4=P�E�y�%=e)��=��<��澼 ��=�R�ct�I�C��GS<��r�M�I�ם<k�<U_=��=w{Ƽ�p=�\�<b!��O�u��z��)=�*=ĸ���O�(�C�|�<]W0�4���� ���3=ѓO� =�h=�Sd�s1��ࠝ����o����-���n�/�"=��m<k�=5�a:�y�<�[ƻ�����@/<ؽ5<�pN=�<sӺ>Y=�pm�v�2��|Q=0�X=a���J�k�}�1= �<�u��<�?=K�<:6�<��%��m�</ ��<;��(�z�p�}"�<jC;aٓ�#�=��#����<�m��x���z�A���͵=�I=������L�͌*<�Q��VzҼ�<�9�2��<+�<,~�<�d;o"b=Z����E=��X��$�XTr�͐b<�Y��ȶ�`\,���G=a�.������Z�=@]� ��<VV=��<�C����<��U=$�=����C
<"/=�Qc���,�?f����=���c-I=6�==c�O�/6�<r�=��|N=���x�&=	o��S������=)�=�{\=���<�lw=�AS=��"=���@��<��M��G;N���*/��d=k7�:��3�9��(u;xVT���r�(�\<���<�kY��3��l=@�J�n��<�w�Ze�b= �<�W{8=����>��*=e��'9�<V4w��)��E���<�Q=�w�ot(;%e=늽�+�[7����<=�?�<[p:�J`��/N�=W��ꨌ<э;�Dd<%� �GFZ�t��<�Ҕ�wY!=��6���<�c�;	�=�;yW�;�#u�����j=S�7<֌P=�J`�d��<뢇�q]��+ܼ�Re��"�<\��
�e.�<x���{Z�] �<i��-	8�Ng�<;�P�4p&=ւ��**=���;�N<*�&�1�`���.=��M��7c<��>=��=<M�h%�<95F=<�Y=1�\=�� ������)V=�1=_��<4�+�4��J��+=����5X�Ud=�u.<��Ӽ։/�'�<8k<��H=q�'�I`A��QS=�X =�|<�w��N:h��=�%=�LG=������x<AX�I\=P�<iy�<�20��	�;��̻ϚX����e�F��ʿ<��=׃E=�U���Ŕ�$�X=w�?=��<�Wg=u8
�f�=�E<��м(R,=@�V=�i��'n�c4��G���5��JI��'�Mb;sز<�v��;��:��O=2I�Z�*���`�+���H�<�xM<�s,��]�<~�==���ʓ'���W=�g=�K�1,�h�6<,�B�c���uX=y�5��S=�D�<�1�<�:=k?Լe�[;FҼͱ=��������N�<���� v=�uf�n����A�Z��<F!"<�<0��k&�����}��;7"4=��e=��˼W����l�$P='�N=��R=���;֞>��>�+ T<�y:߯9�.��<Ck)=��\=��=� ���q<R$=?�=�\%�= ��aC=�,�<U8��T���[���U=8�k=7[;�8=��<}�<�*޻�����	=��B��E�	�*�JTһ��=x��R�=3�6=.l*;��I��r<���<��<JQ�O��Z_�7���P ��2�
��;���<u�*=U/��"���ˬ;6˙��7ܻ��꼥�0=�of=����~�z=��ʼ2[	���^%���=���N���<��:�ڌ����Pp�2"#�7�<�23�!�a���K=�~H�:�9����;༖fm=S������<�T<�A!=`��=Qc�hp���J�%�+�K&B=�"��h�<7�D�j=	U<e�8=`#7=�i=�e*]<�+=ȅ/<�u�<hP�FN���G�=�
���04=⤴<�>�<֑R=��'Yc<���l�弹��h)��Y�e��D�a=<[��<^#�<��k��"���s
:�=�������:=v�/=' ��7=91�tL�[���,�;kCټC�%=^�:9��<�[w�֎8<�7<q��� ���6-=E�w��=	I=��5��p=��w�� �;ϛ�;U�h�y���_��c=2��<��T�b���3=p!��ļy�;��Q=X��ue=s�����z�:u��ct��+<�����<׶T=iH=o.�^�<�-̻��!=�+7�ݒ<"�<S�Żs�N==�W��� <l =����V;D(�<���-�	<����ߧ���<�(���b=��<<iB5�QH��oW�;�\"=f���5�<τ�;(o�'`/<�G�Wj�<r3ּ���tWA�B ��V�Լ��V�yH=�<_�����p&�o( ������	��u�#����<ݨ=�.�B�=��=O�I��s>=��=���~n�u1=\P��P=��U=�R�<��a���7;Q��?Q)=�p��=E��<�H=\
=�%0<m�;;���.�;���|Yu���M���W=���N?����;Nw=�<�_S��2���D�<&?��@k=�ƃ;<#�;�-��{n<ƍW=E碌?������x��<������<Q �;(� �=�+=Ujg�i� =?F�:dI:��?=��p=�`_=-}�<ߴ �u�z���d=JF ��)�����~3�V��Ro<O�=j'�<Ù��39�
<w=Ѡ���Q�fVX�������=�c<���<X��;n;<i2����w<kj��;��<g�<� =��[Ѭ��c��g=�c.=�tX�A�;�Vȼ��V����=Z�UM
�YpD=޺�~S=S=>�&=�3�:�==�c3���=P%=�J�<�8/���K�4��<i^⼨�<4��_=<��ʺ"�$��p�;�Z�<�꽻��;��]�U<�G���:�<�rK��
�=A���~n�����n�ܻ�݆<~J=�^�<���1%��۴ü��׻Nq~�#�7=uj<n����M�<�ָ�BC�<����]=�t�<_O�:U�S��]L��X;���\��1$�; .���Y=W�㼇.^<I�Ƽ�G�<��Q= �H�أZ���w�� ���g��,�:���<E}E�����s��9K�ɼ�{���?D=�G[=�\�<���*�9=Rs��I*�<��o=-�N����iҬ<�n���T+<�SK<P!=�
<�4�pq<���)�=�<=�⺏0j�?�7���<r���4=Ƥ4��i<��7�����3W��]9;��2�S�S�6<˼�q��)��<�!��̘<�nJ=�T<H�
�{a1=�F"=�H�;� =��:�i<j�c=�=b3���K5<���O�<��%=�-=�㼓�T=گA��f���7��=?r%<O@G:/R��ݫ:4�Y=ΐ�<֊���Y+=�Aj��e��@�~ƛ=)���=5��3h�	x�<w�=�s���W����:2�<QPռTL=��<�Ҋ=��>�b�<Fi�JX�f �<�S=p<��J���"N���K=�F���@/��ƕ=��,�'��<`�(=�pE=j���&:����9^S��0�<�i=9�4=X��<P�l=�y*=�b�1�U= �e�!�.�`�!���6��%)=�v<���E==�AZ=��<��J=V��<�φ�z/*�yR;�i�;�6�
��<nX��r��B"Q��ĭ<BY5=!��<���;f�=��<i�<�*w<���;;��:t�<=�M<��l�  �ʡ�;�8%����< �s<�0�1E=�w}<(�l=0����h=��Ӽ���;��9���=۠:��D=�&.=3(N�`=n�T<YR��mB+=�I5<��h<��K=�E�<���X��[��-;Q=�Ɋ<��=���<�]O=�U=W���PZi�}}�<9�=9�F=�ͻ�/E=Ǣ9��J��=4��.V�<D?Y�R��S�=3�R��P�<ݓ���mQ<`��;"&��,[������'�}�w=Q�� �:�%=�hd�2�t=+Թ�V=���a�<V,��j����e���<͎�;�L���ϼ�bs=� 6=��j�0�%���E��	5<�\�����=ɻ�a="�*=����1��e�'P_����<?#l���ż4��<�"����<1]�=q[>�?<�<�C<@�?<��̼�G<!+k��b���Ӊ�;��<�4�-���,< �-=�UL=;��<��Q<�t=�a��O�70-��]��&���S9RV7�s�\�cл���]bJ��>�[�μ5�=:�) <�����;b 6=;R=�r�=R����?=�z6��+���/�j�=��;�X���Y<y`B��^;��9�,Hϻ/�}=��9<�����C=8�O�	�Ґ���0�������'�Y�b=��:���<�k=4ܺ;���<e¼�F���e;��%=8:ṻ���!�=���<yMH<��X�
uB<�� �A��C�%�+^)��V����<�o;+s��OG���M=�y=�d� �H��z�<.�X=��<�<?ٌ���^=�X<c@���jh���$��O�j����ܺ�K��5(=�o0=�5-=0叽�g<�74<��<����=�S��X�;�4Q�,�=��*=Sl�fS�w�����d=qe���Q��6=�3��6���V����<��L8�<<#L=0�<%�[;h�����0=�wd<�B=����_��6-<�@���Ƽ�.��c�{��F�-=�WJ=� =T�<�J��N^=��X=��<�z�9�pK��|�<��<<����A�<�e<���<�ڐ;/�=�z�QI<{b���@wv�Yb�<j�ջU�t=�#;�ҽ�<B6c=�B�<4i=�hL���"e2<0M����4<�fT���=�W��B�<�G������^���_�#�O=�C�����;��5=�=� =�F:�F#:�ׂ���b�=�V��g�<��ˑ�<%:�<�	=����`׼�C;1����j���张�..5�<Y+=��`��#��R=�<�R4=��=�*-=��a�t��6p~�c\=!����=��r������A=����<s�8��6�;�)����ձ��<����<�֨<�t�<�I�;��<
$�)����w�;��E�,�%C0;ςp=�9=��;���&h =h�.=��*�;�=�B/;hY̼�!�{(=)�=�I,� 2<�=�O=��0=j��<��
�C�FI�1�����)c ��!8=�3K�P0�;4�=]v�� ��BN�Ȧ�=��=I�6~:t�	��`�TI���b1�h2��T�׼��[<� x=�����:=F�t=�.�;De�<�;uS<[�,�
�$=2��;]�V= =���R�=�\%�����}L�<s�<�S@��Zo=�R�����<&/u�fi'�� ���ϼ}qJ=x���,夼1$i<f\7��e�<��C����0;=]H>�d*=i�<�!=)�� F7���=n�<wP�<���<�p=�?�<��[��m񼞅^<��<�B"�7��=��=H6��W;W�Rp�<��9=P(�m<���A0����y��<JM�s��<7�g�G�	=h�C�l�<߁Q=ދ9�ߍE=0by�UL��hλ�p�;Bq=�]�<���	�=N�<m*=Ƙ*=�!�<^R<z�;<�0&���|=ST�<���2`7��]=?�'���s=IsC<�A�<����EZ��$����i=���<Y���m;�W����<�	�<��'��9F��i�T�<�b��%�M=>G ��o4��s�'/.�k�x=�<�}9��<�k=�=k��BgC�8X=�3-�I���#�A�Fx�<8FK��'�;�Bt;��H�u$<�(=]=_<n�E�d�s���E�X�3<Z�=`��;äg�<�M�|���<ēN=to2:n	�E6j�m�<��5��=�<�E]��8d<�c{�:��<��<�9�f��+��a�k�TB�=ӑ����?�1=��^<2�;Q���.�Ǻ���^,��/`��v�x��;Eo!=CRs��
g=/�v���P\=���<e�<�=3����DǼL�'���ƼPͶ<]1ܼ[XX�\U3��R+�br���Ѽ0e�<L��@g;<���O���s'�s�V�N�*�)w#=�����&Q�k��8�6=����J�<�Si���k=�mC���g��ѻ\I�a6_���	�U�:<Iee�Β=��%=5\��C���:�we�<WHt��넻j�#=X���j��"��;�t=Ay��2��<W�=53�o:Y=!-=��W=ϻ"�(������M�<et�<R�B=�O���㻑�&��'=�#û��U�<��;@��<Zm�O��<�%	�C+<]�	=J!Ѽ�¼BZ�@8R<�A;�U�mx��W:\=�S�;��9p}��Rx��Q@=��.;=�1���y=T��<���;���;EhS=���_��<�m���Jf;�)�<T����&b����d�*=��躡Fu��S7=ø<N����<��6:y�:�˼L�<�6��
���Z[g=I�#���Ż�_���#�ER1=AbB=������B�SS<<�Dd=ݼ6��G6���=�'�«ϼO�>=O��(Il���9�x���a*=���<I �&m��ݰ�G�=0뼺��<�F8=g�=��_�po��&����<�9޼ތ���:I�L証����VJ��UN<���"q�����<�>�:��)=!��:�{W=@ =�QV<�t=��Q�.4=Y�<PcN���F=�l��Pj<8�|<���VQ�<~|U=��7�"��<�Eʺ�9���J;g+ƻ5l�<5u��p�@�Y=P&b����;�l�<�0='��<sG~<�f*=#�=���<�[ȼߒ=�H���=%lU�T%=�m�=w�=�	T=uyY�we�<>!���v�<�k]=�!����< �5=P0a��L=yݼ���<�Tc=Jѳ;��%=0T'<�������N�&�%�w+J���.��#�+�F�������$� �.�<i>�<T�T��U[��ј;U�</�0=v�=��B������9�ぬ<;�_=�=l�3�:�'=H�<?ع�	Gd=�� =q� =��L�t푻8D�{�t�� �:�q����a=��=��+���λ�� =5kK=%B='-���)=������;��`=K��<@y$��⼒�a�s�Ӽa�4=��V��q��]�/b;�Q$&=��@=�ca�Ɇ='F7<�|y;�?�;膼����03���`�<������5�P�<j~4=~0��5[��@�yO�;O�;���<�oo<�]N=e�<�Q�;3ϻ;�t(=Z/x�����>=��=�m���=HO=�6��ܳP=``2��&�<W�8=&�û�=�b=ˍ��f<A�!=�=ż�%O��Q��0D<����c�๏��tA��^S�ج�w�ü�ɧ<�m�1�]��yZ�\=�-�;����ڼ��2=�8T�[�R��	P<%�>=ފr=����ؼ�<�H=�q���伿m�<E.==����B�T�iJ	=գ�sb=�! ��Is�EC#=���<P~=M��������ZI߹��
=?�!�8+�?ƞ<w�!�W�N=�t=]=��<���C�<]D���;$s5��@���
t=f�;=����u�<QH�D��N<���=]��:�X��!"<� �<�IY��^r=6�@=��=�=�
=� ;Ȃ�<^�D��b8=��2<ء}��!�<��6��</�aN]=Q���&��Q/��S]�}�����'<�M�c~�ܩS<�W=VOu�]j=nﺵ�?��>��Bۼ+���z�I���x=%S=�9^=dK�<�f=]^���漎�y�a���W�=�d=�=0M���ZF=�C�<��<OkC���$�F/��j�<�v>��U!��<�r�@�n� �)��&k<ΨR��v����<��ͼtc?=I�-<`1^<��=cJ/={~�ٰ=��=�|=�8�|	 =��l��TP=�7-���=�ȼ.��< BT������z=�@�<��P<:+<5}�}7�@���d��cA}��z�-�x����b	=�	���z�8��$�O=��B���w;�X���*���:��<L'_�w+�<ͧp=S�=j�<"9G8�٩;�i�&�<�(�����#<+�S=�!8��K��f+�:�h���I��+�<�2L���m��P=_�H�ܧ�<'�(=��=6���h@=Y����R=b��<����^������Y=ڏY�\KѼ͚߼�^u���<6j5<��U=ç#;��p����<xӄ<���=�?#=���5"�����</��Z�@�T��x������*m����2g�<�~�t;�R�n<U�<�ݼ��x�z�2=~~o��(=���-@=��=(g�;4th�Vz���߈���W�<�Ə=��<��4=*}[;�v�:�eк&H�<~�B�����6=���<^�&<凓���_��hk�(2�:W+���9=YJM=�����;REJ����<?<$<>���Z�x�){$=�R�<wMb=_6�K����qK=P<16=-��<��=��c���׼�_$=h��N
W=�f�<j�+���N�a�J�m�6��9=s��<c-����U����.���;�8Q;4�<l 5=�Y:�O[=Թ���X9�-{�j�8=[;U�;?C%:����F�<.{���N�6^9��8=e@&<��=M�[��_�<�%���=��;S��<�z =F9�<5�H<��5=E|=�R=�~f;����c=�K<�:�WD<�%O=fT�:�D�=֊;68X=�� ��%	<<G�:{��<S�b=�:��t�O� �J����'=�]�< H����O=յ��c7�
��<�!=��c��ǻ�m;�
�qn����6=0�=t/Z�ʁ�<�·���=��ǻ�0=�ج���=q�c�WS�<{��%�3������j���2<��;v:$:DxQ= �~�-�%�*�;�b|�<3J���=�e@�":����껥������ �'�g�Z=�d"�� =�;��ϻ��
��%�9i=zI��Y���&=R����;zm5=��j�,�V�*�伶��<�^==m���!���F�7<�>��/Z=L�=I4�Ikx�)�z�C�ʼ�ɀ�7�&=��;�d�L<1�@=��<�#6���=�)��<��<ot"��mh�:�A�C=��'=b�h�C@�C_�K0���n%�� �����A�-�3=[�����X"���;�$�<�.u�S �r�$=��=��޼{�7=d�F=yW<�"&<X�v�.5N<�lP;��)=�k=&��;��o=MЎ�K�����!�%=ź����t�eBܼ��=w�;#�]<�YR���=<D�߼��=�}R��<gm��H=s��;�C�=v4�<��m<����'��;k�9=�s�<ew%�kE��� =��ϼ<�o<�/�:����?��O�K�hj��q��	�n�;=̕��g=YP�B2�<S5��=�,<�U��i;;=�ͼD���M�<|��<?�<6���2��Ұ�<
%C=G�=?�p=��`ܨ�$1��I��Aw�J|����C�Kt}�\N�<�o= ��=�j��P�,�5��<��:�Q��-[`=i��<��Ż��K���T�l�Z�~�x<?F��L�l=��˼!X�x:�<�Y�O=Z�,Z۹��1=����l��<�9�<�Yܼ���<l� = ���B�	<VՀ<�ut=��$:L�Ի0@.=�e�WWr<
a�OI=��5�;zC��=n<7�&}+��	�`�1:��\߼'���D�<��<>%E�w+���E=�rL�󩜽�/��ӊ�P��K䑼�,=%�ٻ�|7:��d=�a�</=�˻���$<cO��J1N=i����1�<E�����D��nL=n�S=yH=�3�> ��=��R�ݲk�F��TB��`��<�2=�a=fh?�b= Zz;�9��+���-Ӽ�����-��;�m���t=������e�ܧI�YD�<n3�,�B=�u�=��~<r���bȻL�=7����7�Y�<�D	��	��~�=M1ȼ=ri=�����n;"���W���̼�̾����<#�s=?��;�?���w�_*��m= W�;�=AS�xB0��e��м�H���<[���]��3a=��3��:;=uB漨�U�a�����u6=-�;f֍<�n�WG<׈=�#�ׇ�AN�<$	=?�w��k��dBF������R=��<�)�<��R����� =)R'����<���`�<������;vJ=3R�;�@_�s�=�^�<2�?�)�ʼѿ����<��=���&=؃X=>)=�x�=��e�m���_:�a���=Cy&<"o���<�BS�>�
,`��$�N�Ӽ�7o;��?�B�&=O�!;��kۼ��:��Ի��4��8=��4�4�o��J�<���<raK�6t2=z�b�;�4���R=�a0=�d=ns漩�J�J����ݼ��\=�����=���6H=�T�^��!�<�c=�=��49��\=��.=��i�4jr�dM=;��<�4���^�u5�{8F<+`V����<fpk��&�;�����0.=��ݺ*�<�������Ȅ��c+��Ս��H_����<���s;��,=^.��X��,1Լ��A=��5q��\=�5)=�:9���;<�g<�<�>=�#\;P��<S~O<�Xl��]�Yf��9
�ĺ�u��<c�=�^�l��;���;wy���K=Q����MrK��5&�G�=��ּt꼘Ĳ<d��E=	�Q�p-�<��,P'����<n���gh�k2W��yv��X7�.��S�'=���*_�NH<��k=��*���E=?�r<q�r�tN���jg=P�<�(ļI�\<P0�O��;I*G<'�:��=Н&�c�q�TtO�^�=H�=DC=�ND=��z���<5M�n�<�S<j�D���c�p׍�>��ۥ8=sէ<�/�H�_=���<�r�<�����8;��<NU?��Ҽ<�]�<��8�j�<�zj=�$\��8I�]�1=�c�;
U�;��׼+��<1�<,ϒ��ꐼP�c�&]>��M�v�a�v��,⻼ ˠ<�5���E<������;�L=�-��ר[=��2���M<bQ<=Jʻ�;�<��+�����Ӝ���<��ռR�2���(���<��K=��^=�˚�iƙ�(�*��L	����㟈����<Q+=c���VV�=1�Y�B�u�%�a��X<��d������f/��= D�<u�ɼZ�:�*[����<��;	š<���<J���q���� ��BE�<�g���菽y� ��'~;�>ݻRN�ٻ��*}}=V9�t�l=�.{����<9�5<j��;�ټ�<�.=E�R��r����<�2��t��+�ؼi��;��<z�!=�*�?Ι<WAG���ܼ�ׇ�8��<iټ�%߼�3>�v��u���9(��J|<����*Xv=�hX=�<�3�:�9=w�=Ɠ��/N!=��[=��^=��93-���T<;�_=������:=�`��-ż�D����#=B���a��팽x��n���x�¼TL�1<�G�<���<��k�S�t<�6�	��*��:.=����e=�JW=ʫ:�uU�;4i=������Ö=P=�{4=pe.=��5=�.�<�;�<�d������U=�����<�2�<c��=qB=q���7<�;��S=������<��=��� �;�
�=�e���8=��ϼ��=	c�<0i��y���Ǣ<k,���8����<�9=q��r=.?�P`= �F=	N�z�%=�G�?8�$xh��<]=P�}=��̯5���=��컑�G�'�̼W��Z��tV��tμ�<����qR�`�< =�	�<�Yݼ�z=�F =��s�u<j�<_��<��z��D+=�=�1vn<�'=�)Y��ѱ��5~<ض�<��<��Ӽ=�;=}��r�<�;�<��W[���»�����v�bFԼ�Bs� /��@!�<SR�;+��\
y<�p�z'=!�h<d�{�%�=�QT�ok�<I���=3�=������;�~μ1�?<�o?��]=�i=9��������%D=*E�=w�<��/=kJ���=�"<N�p�G$�<�s;ɼ���nk<��@=
e�<�T"�
�ؼ���(w=ù��	�A��Ĩ<�a��un���⻝��<kX�:�<��+S�(gG=��9=X0��x�\E=D���7�/��	����<=���k�</o<_P��ts�:H����J���o�;D-��,<3����<�@j<���<nO�]D��!u�<�G��[ڥ�P��%F��۴��r$<8U<��3�Xr�;��Y=��9s麼V=7ܼ,T�<�T��Z�;�@ۼ׆=��&<�q�;�0�<��^�֝�<�k=TeӼ��d�`�<f��<��j<��=)@�<+�;=���<0u=���<bW=ڡ���55���W�ϙ<�nF�qĕ<U�<���<E��mb=�y@�ߊ=��2<�1�`
=� c�p7=ڜ�*���6<Uk�j�
=q�<L���(e�}n�;"A��,� �c#�<�񇼬�1�#�9=�^����'=b���X߅�s !=�����Ƞ�t;�<e^}�����Z�<_:�G.��|�b��=2�;3�+=ȿ�<��<�=7~
<�<=�<��k=��c9�-����<��C;��o<�Y̼?p�~��<��_�Aq�<�y���Ļ��-���<)�D=J���1=��<-!��[:	�e4�<uI����06Q��[=�<�tӼ���<{x5;L�Z�{�=i�׼!�V<@(����D�A8=:v\=-��p����8��=="�]0�<1��<Xd=q�r�aa7<�����<�U-=��3��g<&� ��wc<����~�<��Y=��<G����am=$G`�T�A�k�Z<��]��Q�<���<x�=O=G�B��w��{� =g�7�+$�qL=�\�<Fl];`A��F��<��s<���;�>;=�O����8U��&�)s
=����ސ��J��:D�	����<#�>���m��H=���:��A���=�C*9#�&�ަ=�}o���R<��:�sh���3��E�;�l��^�<�f=������<c��q�='J���z�<⫠<� =N�<�=1��=0�<��;�Z��_<�|==��<[t=
.b��a;�N=�+1=V�=�n#�AfH<V��<]�_<�W;����to=�Ŝ��L��^6��oD��@x���g��x<E���WE����<2	1=�Q��ŕ=/\%��<�=��=B|m�S�M=��ݼ߸>=-XJ��o�;���<��i=d,�<�<����AM���=�v�<T�
��yλ�'�<�i�=���<�J�<�\���"�9�<�J�<I�=�>л��n=�&M�
����p;�VZ��B�f��jv<\���ش<q:[�y�<F�u=��;=�#C��u=yї:y̼*}�	����(+^<�h;�����۸��G�gˊ<<-�C=l�W=��C=����}�,?=�A=��<�Q�<�$
=�����[=��Ǽ7�=x֢<��%<�s��d�6'=6bx=��=�3ټ,���N<{�U���=��#��\D��Z���<=|f==Λ;M>M�p�Լ�Z˼�j=hj>�+/=z?e���;�����n5='Q<C��;PO==�z0��Qy=m1�<��<��9��3=02<K����m8��=���Յ�Z:[=��-������<D�=�.=��˼�"G=���<G-P�0z<��e=�$���:����n=m�v;�gN�;��:ED=��ؼ��<bp���=��-<��� ���\W<�R=�f�1T������W��ެX�Sa��*��a�=뭌���r��+=��U=�$v=��m��L����$���'��]���D�Q��.=z�e�<1-��D�y=I6<���<I^(=���q�;=0��<�=6WN����_�<�y�=d4�=_m<�,���<B(���d	�]�g�����R���)���~g=l��:�/$�|�=��vP�V���nRg;_��%�=��;$�<�<���ɦ�:"\�=lu�<׏�����'Wu��n�<3�\<g�=Qн<�|G��=*="�(=� 7<h�h=5W��;z�C��=��Z=��t<�|�<7ˊ�uX�<�����-=r؜;�a�3ɼ �*=�c<S�<G9<I�=ټQ��=�<3��<���ͼ��d�̼���:����g<�{�Oc���T�<j�K=��<-���D�M=W%�<|�|�᪭<(�T���:���5=q6����=iY�A�<=sP��x�K�6[μ�K{����Z�σ̺Z��<��L��_��Vh�7�M =�)=B�=�E��+(=���<G�Q�����Ṻog�<"�{=Nw�;��=�V=����%��<�g��������f<���<��x=�>n<H㲼�=<Z�#�u�g=�&=��y=��=5L\=�H =��N��Eʼ�E��ۈ;<���jfj:Q`I=쏲���y���'�Pշ<���\�<��<�A��e��<m�a����;���'<ǳ��?=0�T�)�=��=��V=��I=gB��,:�� �m7=��<�';=�yN�S�,;�!���T��ֶ�+n7=`:z����L=��D���a=d^�&s���;�"m=W�-��H=��<��;�H�ܼI����<lR=�F������$D��3i<'V =�i=O���	=�{�<��I=�v��w;U�O< �c�F��6�I<Bq �"��<�c�ҕ���w��;_�=XQ*=84[=`_=���<f�� �4��]�;���B�$=���;��t<�>=�jz��7=�=[��kY���p=�#�ۜ<��滘.=�O<�XF��_=B�G����4D2�h�ں�;�A<���Ӟ;^|��=��<�@(=��мs�4=+Ӷ�����^��5U��Y��<����8���Ĥ�<�7���<�b�<0�<]6V<�&=Y5d��Ȼ�v��<}���"��<ށ��Gb<R>��|�=p�2��+7��	J��̛<�P`;�@=�1�b=�^��h=bJ-�a��7�J�<�\<�<�2��3���<" ������6=�h���=	�>=����`'�Hu�<�� ��G��W�8�l��<FA=�_ټSF=��u=��F�f����d�;�^м9�|;D�0�+�M=�a=�|[�<��=E�����=_���Ē)=�n�<�������<��<�.=Bmt=�<�.6�Z�M�i�/�����<�d3='ۍ<�R =��a</䑼w���,��;���<r���9��>��<�/[<\ߺ
���O��[�[�ٖ%�*�<Z<���F�=FH�=��\<<�s���ٻEz���=�M�b���S=���<dρ�"�Ӽ�,=�yD=���v%��a�<�d��|l��f�:9Ҹ��%,�<0C����=r'H�P��C]�[}+<��=�|U<��=�%�Z�:=�<�G�3���}����:H|3=�1�<��I;9y=�\;�oP)�<�*�)��	0=�p�"j!=�7=7֏=b/w=};��9إ��#�<�O��L�<� ��\\.=A��<Q<ػ�ve��uN=�v��Lr���o���,����:<�ڡ�vW����+���=T��_Q��P�/v��^Y�� ��&=K�:��R=Cv=.lO����=o���{��Z=<�=¥i�R� ��b$=��:�}�;�3.�Ɵ=�)�)ZK�c�z�@['��S_;��z���A����<�6G�4=��<�l�m�=�D?�<�<��S=R�5�����3<W��;���d.�;��
=����:p,=��y=Q�{h��,ͻ���<�E=���<��<�9���x쳼�8<gw�<�B�ɼ���Ҁ�+=9qZ<�@k=���<Ũ+�|�I<��<(�&�!+<�=̻�pP��O��s<x�P=�Gi�2�[୻��2=$߼.�6�|�J�=x�<ocb=?������*��a���V;`Wp�L�<M<�_�Ӽ!�L;uj�Sҗ��ă�i����[9�d�;=,@�:��,��Mû�񻼵�u=�i�>~������"=��#=l	:��,=���VOڼ)�ټY�^<5��;P��:���<Ԏ!=4���{=�[o��A,�����]��e���2�<�Ҽ���<�������<��;'���P�� <�!L=ʰ��jJ��mO=� ^��8�;5�J��`�<���<�>=�=��0����p=�&�<c�=-&=�ļ�� <�+t��O=^W@=����]/���w��S�;p�;':��R<g[
�qS+���>��� =8�*<�!=�(�Ku+=�ݼM?�BP0=>�<OI�<��+w�<Eӻ4M�<--��Wgs���=�׶��#=����s'ۻ����a��;'�;
B��f�<�'�<����$<;M�Z��<y��<Ά���=<�.�=y��`W=���<"���t��?M�2����"=���<|�J<�|O�vEX=�.�<���P��<J���Z��0<��<��E���h���+�XK=|aH=�~�M<;��o���<j���g��<׃�;ؐ�;t:�<�\1<ɺ��)�<��H��;�=~V=im��|�"<=|�"=]�K=c�<w?׼��<Ͻ*<$���m�<��<A��6�$�|�=Ҡ<��`=ז1=��H=G=�7��{��:�<�53�І�<�)����B;�`����<E����a���c;=ڍ'�m8�(� �h`�<j�<u�f'��-<Ot(����:Q._�}Gm��$��w2�L-h��jD��H���\�p�=߉v�L}�;<����<.��������?�;����E�7�����(�;��<t|=����'�k;a��}��4�G=�=]�,����9���W� =��<=�cA<g��;\U�����;�ᖻxr*=�r����<�=�$Z��Ƣ<�DI��0=�rC�/[�=���=���C�T=�����<{�
=�������9 �׼�7=��+��o��]�==5�h;Z	G=�1��X��<M�ӼU�<Ur��Z<*=��<&X�@����R"=������,T�<;�\=i�<=�<�=+=ˤ=��μ��t=G�[:Oi<�H�<t�<l�s=�8��<�l�<��<Y�Q��&7����<f�S=�L��4C�k�߻!ͪ���ŻTS�=�"���b=m�=��<���fl���/����j=i�h=��j�xX�<����q����=��=h�o ���?��&�a�]<�Ƽ��1���l�7?���<NU�Ikl��B��<��E���*=OR��,'�<R�� 9r=鶔<�w=J�o;=p�<�=��B=�o�<�һ�ۜ%�P�<c<��DY�`]�=�+1���h����<���<�M�};�=,^�:;`<`=��{�<���Dr`=��e=ZɈ�����Tk�v{q��q�:�b��l�<˫:=�z缨94�h��	���?����<FX ��ޚ:�������I��ꦼbÚ�xn=���F�ȼrp��m�#PU=��.��Y���x��������'%=�V�<S�%=�G�<�O�<����ͼϼ"�L=���<5=P��-����uZ=t¼'R~�rq'���=��+�B=�\�#JO=Ʌ=	�A��1��K'=�(Z�m�<�釽��E=M̼<\/Y���I<�D=��=���9=�P��j"��/2�<����l�<j>�񝒺��<Ii�ʮf�TA�;��c�_@�<,Zj<�Ω<@��<�a=��,<��,��{A��۬<е6<h8H=I|�<�4�;�N��R\=�C�<�1%<�	f=:{��~=d=I�a= g�;�F��1��/=+�E�<����	=l�p<~���<�4<a�87=M��j0=vr9=���<�j!�n�M=�3=J��<h�����;�o���H=ľ��3ɼ =��==��3\����<\`�<a>#����<X<]��A0��l���נ�)d]�/D��@�<�_=��U=���<��T\n=��R=��A9�#k<[5v=�9���<R�/=ێ#�N�׼��_=F���.�A�`�r�^��i1=$�1=�����j;�死q: ��� =�����.<���	��<5�=��8�l�:�%�;�D=��u`@�VG�<em���?|=�扼��;�s!��h3=1H�%4��/�u������&���&�dy=<��F"�<�8���;�&3;{:�;��<�m.���;_�<��_=�_M=r��/�<��u��Tl=�w=&b�<�*���ݼX��!<E����<"�6=�|�� PX<T�V��jg���=?�����b�X<Dh�__�<���Q�o�� :��;����P�q�	=DGs=��<�s8=��i=��r�\<���]3ʼs��<��b<����B��~�g�r�=^U���{���A�<�F�<k�=��<��	=�pB=��"�J6»÷j����"�<�b;<�U|;�7�;��=�I=x@�.�D<L�<��2���C��#=�sB=bh�����.�K�ֻ��Q���̼�m&=Z�o��~���"μ�=�=Y�;QTl���=�V���m�Z��<���Y�i�.C��̓���ۼ�Rh=���<ȯûp��#F#����g���ܼv�
=Pս����<.;=�m��&�=�E`=cH,<:������ih�L�/=߭�=P�/�L�<{,>:I~Ӽl=����1z=�Ǽ���<Y8��qk�NSj=Һ+�V���zE�~@�1I:GQ�<�5:�P�;ܱ�<�����=�>��\��<(��[a<W��_���2= �Ҽ��n�=*-�*oy�W'=F�ʼ��b�?�2=ETI�4PY���5=��:B=��<��;z?.��.=��g�;���<ܡ�<��=5�`�Т=}�,=ؼr<��B���=��\���?���-=�H�<Q����
p�p���V���	YL=A�=��Ĕ<n���X\P�}TC�J���V=�-6�D�o�}�#��G�;�U�Q7�<�Ӽ�#�<��t�K+ͼUvH=xh6=��<�=1�Ɉ�<%�<�����%p<�Z=��o=�6Q<m��������u=*�)Y���𼈈�<^.I�rjI��,=#tv<��W�={��\�4='&T�g��<(ر;�G�F�=�=�s��ɼ�v=�d�����;��ۼ'VH=*{=\p&�@+<�<���(�<�L�ٳ=`:�; ߫�p�һ��<�tR=v�==v�<�7<��S�/����-5���J=�"ۼ�����I�Z�=%���3K<X��iq�����;��ּ�ˑ���(��Z�:�����$=g�`<d&���%=�#=�i=[�2=��i��Lz��K=I�6=a��� ;.�;��j�i	��cZ=on2=/"�l�L=�W���`:|-E=[�_</pE=װ2<6�h�}KP=����;�A���\<�_=�U��.�:��0�vi=��˼�=��|�R��tf�M�=��M=NK+=oqG=�w��a�=���:�qI:��;9:Ǽ��mC�<�k�<p�:G�]=�u=�e;9&�G�4��lm=
J=d��;|��BA=g=IL=Zy��)�<㸼�	%==c������h����~B<7P�w����A�zzd�݀
���ƻ]pĻb�`���M��~B�9=����=�� ���A��U����#�G��I`8�d1�
�=��_�י�<M���q�y���<��k<��&���l;�dD=�v���=pN�.i���!����;#����:�b=�wݼ�7A�`�,<�]?=�y�;�t�<��R�O�*�ֹ	��
=m>��B�= ~�<+���n~1���=��e���Z=��<=��м�)�<Ƽ��	�^�ٻmX�!Dr�%*O<�17����;�3�cr=f��y�-=X��xD=�ŏ<��ƼO�<�-�<i�=�±<<�s=��_�{fZ�(X�;ԁ7<7�����;`��<��Q�1��R�`=�Q3=�y=DX��<��ie=�����<��<"�)��1һd���W =@����P=�1��>Ｇmɼ/�c���m=�;���t��W(Ƽ@ў�g�:=y5<];;ʏӼ��ʼ����g���Y=^�r<p`����Ӽ:�ڼ1�<��L�46=�#D<���<��N��Av��Ѣ�|�v+�<wǼ��=9�4= d=<���<G�d�pw�;�^�j(�:�4޼�(I�h�5=ն���[=�=�96?�-&=c�@����4�T=&Ξ� �м�3����F�;��;o���yz�Q�6=�bF;i�O�`v��g�j�K�0�ij�<Ǩ</�<3�<P�!=2�b���� ���U�Լ�n#<�
��	U�qJ==��ܼD���ǟQ��?=��L:SS����"��Q�<�+�
�=`2�=d�<���Q�N�:b=3@�<��<Ex�<�Q<�:����=L9b���=�YK��ݼ��Ż]�w<�6�<���<�/��À���c<ODv=�cں�C���P.=��2=�<��i<���<� ��������<l�:���<�b9=��5�E�=H*��)X��u���$� =x�=a#3���t����ׅм�g�<���<+C�<_	���n={�F�|=�Y=e0���b=�\��ɂ����;��鼒�%���#�%�)�8	�<!�8�� (=f�#������u��;�C=;Sx=��<�q�W�ȻX��<�7�+���q6b�<	+���_�q=���L����W�"��T�<��,=>K��=@�<�[�<��p���=�� =�.;ۇf;�Z���y��s�e�m==��{���V<��<a��==�]!=��=��=�n�<�
Q�k�a<�%&��Q2���,�"�<��r�[�<J�<1%=2Ǧ��P�-�V�W��-7�����Os�<��R=��>���k=G���z"���<����'�;8�?����Mu��kR��
#��I��';5=�6��� 5�2s���|���;����;Ò �Z�<8�W�-=3C_��H!�S�):� �<�2�^*�;Y�2=���<��N=%�3�wq�{��<_R=KF=�5=�q���A���<լ�{�����r<�W���8=�I$�f>=7��]�<��7�^ܩ<-�=���HV�b#Y���G�r·��0ʻ]49<�2�:��=�ǘ�}�E=�L�0�޻%�<�V��a�;Ȏh���M=�q <�ܺ;liU=-m0�+��<�ה�cX#=(�`=!=�?Ǽ&�=�ގ��'����5�"�;v0�(���=T�6=1�N<2v3;l1"�~�=�Rm=�(<�H�<�,R���7 ���)��	+�e8���v�<���:ҴR=��f��x�8p����������j�6.D�N�<����x�Fj��g4��Gf�B�6�u~q<7>i�S���mݻ�
W=v*����A<gm<8=N䲼KB��r����8�&��2=�����e+=�y�;yHH�� <Qw�<���iL<�i�m-M=��v� '=��D�@Q�6�I�<�TA=��=�/��ǔ<�X=�[=��D�I��Wν�A�U�D27=p��j8=��/����QY��el<{��<��=�OI�{�9�#�x<'V�Skżx�c��\�����W�<ן �/W4=&/���D�n�C�MI�<%&z���"��<��<l�	���*=SN.=��8=`'�iĻ|�:��0K��1ݼ16�H�s��Z�<q8=��3<I&F��"=���<S��;}�=?�2��h(=�==�o�/�u=y�W�з�����g������S=�7�<�<-�<6D���H<͏T�G�ٻ��O��==�I�<K�=eX��Y�k�+��F�<h9�<��X�n<��3��h<�VI���*�,䨼~c^��OԼ��=�a=��f=�iX�``<�2<��;�;���e���a+�~��W+�,�c=(�!=A=�P�(y��IH'=���٩F=&f^�X��y&l<����QH��q��a�5��,/�n;�<�1�<���<Ӯ����<��¼�b;g�K<���<�7�<3J�<���;n�<l� ;�,/��+=-�	=��=^<}�m�(M�JZ̺Ĺ�<�B�(�N� ga��9>=C����]+�]m��#����y����1=�p��I@��1
���<��A:����.�<CGG=+=YE�<Jf<��v��O<��2a��b�*�=��G�ʟ�D�,���S�*�x<)��<�=�O-;�L�;��P%�<�
��O�N=	Θ;j5C=FK�<�[�<*�=��<r�_��7�r/�:�.��r�=K�
=��!����d�����:��
���m�� �<��2�*��<�[��
�;SW������:�^^j=KJ*�[[=O�%�?EW=V��;9�$���x;��'=p#ż�1=!��;����A�<?����R={���c��% ;i�;�3=^��;�A��f=T��s�d<�3L�ٸ:]+��T�X�XPQ=�A�VR=!�D<��5N�\�=�L=�~�'��<я��RU��<�6=�w'=���9�<Al<�K�<�<yX��_���(�"���=
�;=i���#���a���!��Z�;v������<��N=6\�<Z_ü"�b�#�k�|�B���E��=��Z=��_;0=�;(�伞T5�r�>=f�<�*	��U�N��A�u:�����B=�/x=��$=�����;�;H��{K�И��@O<tJ��j�Ӹ�=7�>���r=2L�<�v=O^2<D-
����\�;���)=**��7hb�H�T�w����<���Zr==KK<|`e�F��<�z��i�<�_2������<��p<	;ϼ������\�����u��;�9��!=N��;S�C�c�S=�<�Z�<�);�0��;=�m'�Df3�B���=���:�[�
�*=�l޻VQ<b;�<
>k���0=ȃ�<"ż?/T<͚;�5=�L�<�`ڻQ� ����Iu=0=�Y��'M��=%=+���H����'=wcx<�=��:��q�<��9=X0{��v»?��;���<��<xwO���Լ�H�\�ﻲ���q�<I�f��`W�����`��;$=�B�=]������O!<0,�;�ꝼS�s��	o=yFv;j�ޱ��z��ӢB=�o3��=�Ie�B�=���e=��=r�8=�=?���4��k�;��<=$�X���(@W��~��l]���� ��F���+= ��⺼3�1=0�����k<2�E=�n��'`A=��=���z�c��W�<�~��s�{:����������<Q�<Q��</��;HmǼUD����<������;�r=a�@=�F��n�=�H��.}�C>E=��H<�h����=�"�i�<�S����j�!;ıf=�]=��<D�<�o�<'��=�PD�0�$= h0������=ݸ�;˷+=�����]<P_G<��I=�4@<��漪����$<}��<+y�� t]=
='O��&��zd=Ք�=��R�����l=� =��M<0Ż�����=�;G�!�%=8�+=뾃<Ԑ=��<��(=������=jPмN"�<㰗����<J'9=f��;3}��bFR���d<�^C�=�h=�l=	Y�����u�#��;`��
 
��D������1=��;��><br���-�:=�F�]�<D��<)�=�q���K
��z\=�GE=҃�<��a�<�0���V=��\<Z��8��4��R��?�;���<��U=���m�g<��t��c=���ړ�<�G��=˦L��k�<+(����;m��Y�<��=%\��U����=�</=c���(ͼ�X�<����l�=���<��I��?�<~�_�XNS��<`����,=��_<qIH�J>(=_{T��D=�<>�T=�A��9m�<=�0�D�R=�TX���F=g/������	�=���<vd�,���gZ<��<sq?:M~<+`��S==:��W��8=4�<3!q=V�/=�����{�DAK=���<��$=�� ��}���#����<���29I�)9�<e�i=�����??�毶<r"k�� ���s�`
�;+Pu�iDU=Ǫv<�;�*1S�����X�P�(�?�8�[�G=Z�!���-=Z��<U�}�z֫<��=���?���~VQ�3�g�v�H=��<CGA��G5�y=�O�<�$�<�%�<h�d=^����<�ܼ��&7<;49=q��<%l=(0�<5�����<Xyq�v9,<��p{���<
�t<�� ��T��U5����</U��?V��&=�{K���7=�GB�B����8���<sq��-�
�'���=�<��<ሓ;L����g��M2�Z(�<�ѓ<u��A^�;y�Y<E�s��RH��(���껲R3=ʅ9=�!=�lr�Ј�:x�=?*[<��7<P�G={�
=ȅI:��;m�r�A���	=K������N�ɒC�L�<�H=�*=d.�</Ic=P��=d�9�,�O�3a��n̼C��T+�:��P�e+z�[ʼ>E�3� <\�o�,��<�!�<�7�H�"ņ<ۚ�<|�<�5���=�rD�z���%!������[��\����k=�+<�`�G�=)�5�H�1=bP=�����S�=|<f�!=X�C�Yvμ͂=,S��=�ε;�#F�Mg��b�<�a�>q=󏄼�6=4I��E�<@=ټ�iO�ƥ)���=��2=�~x��}�:c���j=�0,=�+���)�=��;�=<=���<��F��E=���<��6<�_=���<8V���=��o<���,rY�u4#��-�;��==�{'�_��c�=�CV= X������]7j������2���2�<���<_��96=�|e� 䊽F�p=?'�<v{��%��<��6�I\u<ТƼ=B�<�_g;7n ���;¢
;��<i�2=X�F=||-=�yp�����<H?�o=[Ш<f#?�O榼w��oe�*�+�p>�1?Q<�A���R=nYϼl���� <��=A��'����5=�=7����q��g%=\����ڼ��e=ą���Y��Th���^=o#=�J=��K�x��H}<�̇<)/���>=3�N=�vr���<CD;�?��E=#�<N,=e�
H弞�H:M�R�<nʼz��;�c=�<�ϐS=��{=�e�-?�<��0=z�Z=	g���_=4�<�u<��y�_�6��'x;��-=�Ϗ<sd=d�<��k�<M�n���
�OfH��ӊ<˄=uC��~�}m�:>("�?�=��1��Ǻ9��7u��Ⓕ�u:�'�d�%�%������޼�k�<&DZ==��<\! ����<v��(��'v<�}_=ށ2=UAT=Vy�<h0��n<�f=���2<��M��|�<�ü�q��6����}����<�Wn�4�c�K�������<�!�������ր�R�*�1x����;S�&�v�I;��ͼ)����`�]n�:��c�?G���:V=y��ES;"��<�u?���]�t@��1�3=�!C=��<U	-��Ӽa *�# T=��}=���9w�<1�	=_A��P/߻����\Y�^*= 	��=�;3Ao������`=D�¼��>��'���-=��f�7�b�;ZP��Ad^�{����c=VN�H�0<{����YK�0'!=��2����,�=P������ڬ���s�T蒽�n���I��%\��nT=
y�<�Z��@���N�F�@����<�++=8��=ɚ=��;kD��-s=G�뼣��<�~s���<��;�}#<�uS���1�M�$���<l�(��%�<��@=#��<]=4�c���C������/���/=̿d����<�V�<��>�h�4� =|
��=՝	=�Ȏ���O=L$K�?]��P�<�W5=z�q=B���;�_|�<�߂<�/�����X�<RB=����n�;�2�<ˆ��HN���~鼖=�=D�<@H"<���#=�g��_=}��w=[�A=N�<~=��@����8"�<��Ƽ�i=?^ü�=2��<��<V�=a���f�;��<u�<�k=�=Y=�0��d"�t<�V\=2+>=yǋ<s��<��l���*=C�"=9AY<@��=Kf���>4�1(ʼ��<d�.=��<�<�z�=�e�$�<�0�h=cka=�ܺ;؅�<>�%=*�绂#�<��;�R=��)�S��'�M=��� ��м���<��u<:��:xs(�*�'<v��< �r�1�2�?�`<2R=�S �����u|������<Ұ*=�2:;�#='�:��#=�/�<3�ؼ��);��6���̼ы�:�;=V�=��<��v�<�{�$c-=�5=)I�������<���w�Z=��4��»���Q=��<��\��@w=MP=Xtj�>�A<׭(<�%S=IF�<w�=Y��<r����=�u�w�
��a�)������<eE=}�7��E��f�
=�([;�x'�BSD���w�%5�Q�K�f�����=�ڽ;���Z
(�Ə�<�d�<���;��~<*����:��1����<'�b:�<P� �G���
����ۄh=�bG�3�r�Gg{=�&;W�<�ǜ��C=���^�:~f��ư:ɫ!=�>�;�E_�N)(���;^r=� !�n�� ��� �k<���<�f�<~�<3�<b��%n<� =	�=�f�<l�Y=Z�w;�<Ã?=�@�<.��qs޼��5��U+=�{A�.[�<)��3s�{�k=�����<�� =�9�s�d������Ƽt2U<d/+=Jt=ߡ�<��K�D�9=U�u=�o���#=��$�T�r�ٳ=���w��<N,�<a�.�_Z�h��;�T=��<ͯ���$=�s;�oD=5���թ=���	�
���ۼ��f��9=�=�O�3Ȫ���<�iw���,�*��;�-���F�+w�<��=�!;!���u2=��V��'={��AP��FR=:�^��=�L�<}�O=}�ἡ3*=�;6��03=:�׸�5<�=Ä-<������Q=sVy��I���Qa�4�չ�#;�fr��_?;��3=I�UA<Jq���LD=܈h��=�FS����`;; ��P�� ,���o���d-�ۆZ=۞t���?=b��?�;��<�!=�q�;dk�&�,=���TA<�H����\���f<�:-�N��#g��F�=~%#:\G�<ɼ|<�^��XP���;<	��E�=���<��;FFZ�r�Q�;�5�����<��i����<��S�E��`M<�� =��$����� (f�F��;�Ss=.�<�:��U[;�I�k�м��:s�R<�1�ݨh=��=^2�<�CR=ztf�����)=|l�;��;Q4��=�D=�Ju=�O=�����v=�� ;Ē[��UO��H]:�<���z��F˻r4K<�Σ;Q����N��6=.1+=��<�N�<t]�<�-�1����ݼ�*H�.�Y�!�B</NB=	�<@?�<�ʩ�m�缤R=�c���)�:�2=T�<��
<HwԻD���S��s�N�H=��=���q�<P�=2�h��a(��;<�u}�� K=^�P=_=I���<�K�g�	����N}K=S�h�� =�?=b�;��V�Xy7�<UR�v(=R��8� F�&�Q=�H>����X��<E�+<0=��A����<uA)�ΩK�&:�<�e�;�2����_:<`�̻-�9=̖������k`j�
8{�����%�<aM�<~Z=T�<�&�7y1=��<o��<�}q=qgY���r;�,=�E�<�kS=�4Լ�d��3$�WGS����<!ki���	�DE�<�.9�'�@=2=��;��;t���J=�������R�<�(�<z�<�»���N�N��,M�~Ї;`5=?���t�=�과TE��U��YӢ��d�5I�<x�z#C=d��?�鼳\-�
���A�O=b�@L=D� =��}=�G=@�W=v����<O�q=#�� �<J�<�1%����IϘ<0嚼�=q�<�P=j�8=KT�<܏B��B���[=��ɼͧ�<��R=��:�Ч<�C:�l=Kg=�M4=R��1�&�X7
����;�Z$�Ua=A���4=�#h��=R�&��������E=�潼��`=]��a�Y<U�@��Un<�mU=��=�<t:�<$U�c�@=-�<��2=�~鼧�=�D<j=��9���.=�w#�;�2��5$�w�'=2���17�z?���N��;=.H���Q�;�<�������d=8�+�v���G�6b=���� �.J�<�5��ilA=�#��
�g=,k鼒o~�]�=k����
也c�::�0=�������+=KO<���;S�ּ|�;�c<��D��`���Z�;����E�:
�;��N<;{=h��;o�'<H�`����<�@<�6~=4�=�J=��b={.4=u'�<�f%��:������ǔ9=e<���<ѩ�������1��B~�(�>=Ve�c�L�۴��uy'��^L��q;��E��j�<����<$�	��l=��3=M[P�k$z=�zռ��<��e=�{P=.9=��%����<Zh=x��<F�:uN=���/�T�<@R=\x=O↼�K*=
��,�T=V5��� =c��9Ox=g�ü�ֽ<�f7�96i<����<�:nRZ=������HD���f<g�ƺ)f�8Gl&�v�m��{��@-�D�<u��;v�;�%=�	<k�K=�gw�'"=ث��!��?�ZY��s���UĹ����QT�'�7�m�J=����pY,��'�=�Ld�]���A�h�>*�`c�<F�#=5��<�2�<-i��Al���:�ı6<��a�_���׺���:��v�Y\5<kEq=�]o���<�Xc���:��˼����~Pϼ�G=.�-�(��O�=:٤<��=X1V=D�Ƽ�ˊ�o���Y=���<�Y�<�a�<�&#�7t�Dp�<�t��� d=��<I�<����H<�;�=��$��� ���Q=��ռ�U�01ʼ�O=���<��A\=�u��zg=+��<}�;�(�e��M%=���:�ϼ/ ;�`�<>CH�����2�l�dP�9�#�/�ȼp�k<.[K<� =�i>=Ru�<�4<�ZH=Q�;�đ�<}�<���8d%=(�d���Ir�<�T�dO"=a��������<)�L�*�&=�:=ear�7=l�h=�l�<z�����;hKr��<:P�4����H�;~�<?�＄=�<��e���G=�I=,��df=�����{!=4�"��	=`"-�;l���W��*;Ә<�������SM=�+�<͊g=p<C<�1<�{�<�B���Q�<�\�<l�=�5���Y�mT<=��ûc7��iκ���<Z��6B���g�@�<��U��64=H�!<��+=�R��:��<�/�v��;�q�=�#��C=�F��;=�,=�������[��<��<=?=K%�<��t<P��}ef=y��;ZeԼ�AY�4�8����;���;�eb��c<��<��6<��^���#�);��<Ř��¨�n�=ĪG=�+}=����=Zh��y���L�<��+��KY�Hd-==�i��z��i�¼�93��K��K�X���<%����2�K�<�yo[=H�!=x4�1���ڃ<�-=�%��e=��<��~q�<��浘�4�4<��<�<.z�?+�R{<�1B=�=�7w<�+'<a�?�<��统�����^=�(=�[�<@�@=��*�P�E�P��<��U��zD=�?[�w�B<��<N��<���|$���y/=��0�vcD=R�;%%��z�<�ü��<HH�����Dқ��C<�AH=�����J��%�c��;~j=]�<C��<Hwi��M=�h4=IF�<K��;@��z�<�W߼Y^=֧=T�ּߨ���p=#�M=;�=��B�=9=�S�=� �;�=;���<z�������?h=�Լ\O_<��<��	��a�<�'��=DC-�X=��<;�<I�Z=߿<��:�{a*=��@�؆�:�[w�
�����%o�vV�<��k�p�H���_8<ɮd=�,�<G=8��i�<N�a=�=<�ǥ���H���������<��Y��$��n�!�J�	�.\����<�t������_����=��#Z���K�<��\�Uv��n]��9;��q�a�l��e�=�-�9s�Ƽ)�̻RG4�Q�
;7=,�;%*����I=X����%=�2B=A��<�%�;F'\�Su�1�2=���9==dd�<Z���l�{,�kn�GE=}8�~3=��i��dM��]=�'�5H���=I=�
�<�BѼ��;{!�<,�0�H=S�$�{=�h��� ��Q����<
�3^`�~�m�7=J�,���<���\�<l��oH<�-����<Ϥ=_b���2��г���J=E�<[#=�P���G��u �_z
��XW=��\;Y��;H�<�b=��==̕f�z)7�8��<�*=�M��ɍ<f�_��_��F�<�(=m��`vF<~ټ��6� OC���<��\=�dԼ��z�nK
=�2���S�ަ!=6�=X��<�黣#�*/����3=p<���e�n=#�J���ͼU�=g<����;�0�;4>R=r\��)!�����<��x=���Ϥ����$<�t>�_��<q�A=N�<=��<�.K=�w =��=���<��VF�<;b���=�<L�~�Q[]=uC�z�o=��'��M"�T=�l��χ$���;򦐽��7����p�׼�A[��	t��e�=�%�Ʃ���a<p�９m>���4=��(�=��M��G�;�b'=��*Hk��6N��.h=r�<��P<��\���W=���@*%<~{b=�$=֠o�`E]<m�]�7���=�n�;)�ϼY	<�8�X=�9==�ݒ�s}<)���%<X�p=T� ���$�S�&�</�=ڠ;��S=�bJ��SH��=���T���h��~J���=N��K0=�u���S<
��<wM!=�t�;IV�}.q��~=��<��Ǿ��5<H���T꼶I�<K�f=ct<%}�E~��b�<�M���<���[�zU�g�.O=��1=�x��+���="/׼W��<�vn=]]+�B�\��&=ꜽ<�Ǽu7=��	<5O��!�:O'��|ڼ����؈�Ӟ伈=�O�<�w�9��L���$�!ч=e�<�(n=2��p�<��_==�R=��8=h8=�K�;�dL=��Z���.�i��{�3���a�.I���Z�3=� ����e������_=�h�<�+��6y ���%�tcT:�����,�wt ����9���;��=J+��>�<f����Ⱥ&:�<NG=�l<���<�1!=G^�<��l=p��;]/#<#U��J�<x��$�T<�`<��)�;�������O}K=���<�!���S����*Z<~l_�n*�A�S=��p_��ئ<q��805�=�k?=�|��F=��=C�#<�m9����Ynq<{➼�.-=�F8�?�O;�����==�vq=��-���=��=t7�:8|�o==ߺ-=����=Ǐ[���G��G����<��?<.�k=w���L��j=q!m=v���: �<�O�=ڟ��z=�W#=��f=(<��km:�<=$q�fg<<���XL�<K�=��+�Ơf�BtS���l���b�4W�<uWN=.z����Z=d
.�����lAѼI]��`� �W�h��!K����<��D�¥}=�&=1�?�30�gn���v=��v:&=j�V=Zټ2�<��=�I3=!P�;M���if���q�<�0��dN=��� =D���	:�~=�iC�E�=�C,�޴=�a���\<�>6��B��=���<E�=00<E=/TL=J�=�$=�����4Wj��AA�����\U=YzZ=�r��<�P��}ɼ��=�� ��c����w=ӎ�<ոA�E>�v�W=MJ<��<8�O=�A<�C�:��
=�ϭ<]𢼺<i�X�U�D<>1<�c=���F3���;����E�`=)�<�$���7_��|���L=^�3�<�=z��9���iz=��=Ց�K0:�]�;�nO=�B��W����4���=��=���;l��<;�T�ы�;##=� H�����ãR�fjb=��
���<�R=�ݼ�ӯ<숪���=�[A=ޔ =��=��9Nf�=��;�=���G^��<=VO=D��.�G;�q��荶��K�<��!<!�.�]�G���J��V�<B9Ӽ��=��:�.<i�(��(��[==暴�d�_<B{!=�&=)�z<\XO�V6s;Gp�<�ԯ<,�A���g=�v�<3�]�{�����<@�<W�S�ʩ+��3=`K��L��W=�/}�8*ɼƖ�<�i"={�C='ּޠ:�]I�;� �/YP�Y�����5=���<gn���V�����x�#�߅�
Z;Q�h� �<fU�<�Z�<葼���I���#���ú��<N���0S�<�UU=���<�N���:���2=E(<�N�<���jDM���e�=@¼ۯ=���G&��y��<�<��<��+��]1=� =�j��l�:�Zc�<�T�Wb׻�x�: ���?,�)�
=�h��d�Z=k�.�ˢ=�yŻW#=���<�A=m$�=5��J�=�u�;7����T�<�ڼ�{9=��U<2�=��)�?�һ]%y��u�m��4��� O��ݥ:��Իܣ�\ �o�/��J�<�pg��f=ئ�;��<@n�6[~�H��r3;��J="�L=�~�<��̼�I/��wU=�@�}�<DV��j�;l��"��<L{=�m=[�=hmQ=o=ޢ�<��ab7=�>_�F"�:�(�<<�$=��M�(�r�<��=ݢ��P�kB=���<.{?;����ҡ��X�i<k�ļ7��7�N<�M=7	0=Le��^�^�X����ռ�J�<�t�<N�$��<�ON���Wm=*�"=��V=��e��gмB����<=|���=�¼{*\�n[;�x"=rɼ�\ ���o��+�F�?��|�5=+��=＞�< O;��*��e;����*�<�w�<�����X���8��n#=ܭy��^�;�&<=C�&��]=�gj<]�%��y9�#���3���/���<v�;�y�[��<E2��آn�n�F=8<==Ƽ�Ύ;}R��2H��F�r^]<���;WU�[���[�i<��<. =���<Nk�ǈ����w<lk�<�[�NkZ<Aҡ;V��;�[c�k,�;�^G=ލ�'��D�<�=@r@��ʉ��&�r���-"<����d0���R���P=}7=�w�@0�<�,�����E
;���_}=�[��*q=�jA=7G<3I7=^�~�ˮ�M]<X�<K;�����˴:��;��$=p��l��;\mK=�Z<�R�:�v�<��,=�=4��8���y��<C=��ۼv�ػNb�v�/�T�ǌ�.���X�<�;=n�;��$=���5���_��/Z���%W=hڻp�"�i��c=ő;:@8�o�<S���TA�<C�<0�q���5�E�"=���<dCn;��f�x�j�9;��s=xv=��N�����ߖ
��)��X����<-M?;�Cf���w=wgz=����T��v=�����;.!�����7��/����F6$�Sɗ=��P=���=-=�=����(=߬A<��_<Ɏ=u��=�λ��Bg�Ͷ)�;]5�?��8'J�0Y6=n/F�X�=uJ=֎l=����������b=I�Wd`�t.�9��A��������a�=Rd�<G;<=�� �nQ<'��=س���D��j	��/=�c�iN=i]8<�pt��׻?v<�<�QXE��Ү;�է��v;bS=��;	=<�	�4W=��=T���L=�uG��»��j�	�;<�ּ�K=��=q|��gj=Nvd=�:�Sgѹe�z<�u-=r� �V��<�2=�y��q�`A]=�K=f;E���f<�){��ld<$���[���dG=˼��O<��;U�= ��m=Yb�<~%I��m�<?F+=�P�2H=��~!=u<X�=H=�?�<m΁�!wU��)3=���)�$�ĕ�;c��<�8⼇:��<N�=����svE�00��{�&��Q<v*��+59�A�m=(H��k����xT��<Q	|=�;x��#�<>\$=�^�{�\=::�)K�LJ����R����/dq={�M�+�����B�[������)=}�=Bf����;pڄ<��1<���<?v(=pɼ-B�("=6�.����<�]0=�<aa�;����~W�����@�:¸9=
���!�^�'4q;�-лm��8ͼ����!���)���*��ܒ<3QK�(ܳ<:=t=��<�G;U�E��H�;�F�<� T=*^Y=V��R=)��e�����r�*���=ܴ<a�=~4�<3�
�����(f���&��"S=�$;lOc�5!���3���<��9��==B�@�i���(x;��<{=<Ի�֩<l��J�׼(�B=�{s�$����
=����q\�*� ��O=�"��ב�Q[Y�3�-�(�&�~nj���ka�"?�<��F=Z�༜�8=*=��<qi==�`�'���m$/����P��f<u�μ���������q<�����?=q�=J<������<Fv�<`5?=l�==�Ͱ����<���<��E� l�<a�<�=K2=� u;G�0�d��\����b��<i��<O�:�b���O�DP�<��`���h=x����5=|��<�ҼO <��$=��3��AG<�G��;=�}R=`N]=�\E<݈/=�=,�3=ǡ)�G���`�<��r� ����ڄ=|t��%�	I=eF<i]=�D=8U��y�����=Q�n�\�z�ֺ�<��ؼ������rF=�1k<��<������h�p=<m�<!�|��0���Y��zV����:g�ʼ��(=.(��,&�Q�<��<QA��K��<������ü&����NI�����ѹ�eT���=���;OdM=ī�=�8��Rͼޅ�<�8<�U=��7=�����wG�<�6=6!���C����G<#E�<�(�;��Z���R��6��^;�hj����N�k�D<��0=�ռ�;�ʬ��Vݼ�݈=���3=DA�<���<�� <�����&=��<j&�����v7@<I_�<���<�a�<]�:=�z<k���"�����F<����W�	�@=�չ������7�TC��\ ���P=���<"k�.0���@=�d���}<�d�=��U���<n==L/`���#�����ޞ <}��<���g^６�v����;�:�;J�<q�%<b�l=��0�<%`�=�*�<�} =6��ϴ<�W=��
�= <K�	=�](=�]s�%d<{J=�|�(� =�s��Q?`<n�Լ�2�=�\-;��,=�"�;Ae;���<��kD���5=�<�<�5߻��,=��=��=��,=$����<zl�<��C=Ct��)<7��I��E: ��<��A=��L=��<����4��#��š�B�;kJ������{�*=��	�У��)#�<�����~=�E���D��y:���<��{�_�W
4;j$�<�Q=�<�0Լ�n����;0�I�	|��e�¼��0��t�$���VX\;��<A��� �����K=�҆�i��<�.=��F�j=Y3��W���{�C�}�3Z#<��ܼ�B�a�v=�i;�)����x������<5}�<s�ݼ@��x�@���F��K�>�X�Z<$.�;%�b��'=l�P�=c�<Y��:�o<��<������JN��� L=�J�<"D�&a=�U�@���Vļ'�<e�<x��;$��<h�!���J<�Cs�?F��/=`�Z=�_�:��5=A�<*�<��+���N��yM� ��:�w�<�p��Z�R�>�=�v=���<�e�u�
H<��U�[OL�c�&=b>�<���;�.=_l<!Y����[<�O�ۜG����ROt=Eʗ���<
����x��3�!�H=�U��C���;���(=���<�Bt�\T�<r��5]=BR�~"���a=o�U����R=�x(�����\*x;>���ڼ ���>�;�a����;*,���<KF���=Q3-=�=7��M�+=9�����~���Su@��P���ɼ��x&=���H�<���~�����g�K}�<O�0=ϰ�������Q���$�F�@;E�7�)Z�)�<�?T�3$E��|�<ȼ�U�z@g=��<��,�������[
=m6)���@�*0��-��<g�
�����w�� ��I;�:b�B'�}�\=7�9=!�/=�7����<����/=�6͏�#�R=�\C���B�<�7�CB=�@�;��
=�x���/�,1��g��sTM���ùNk�j���s)<�0#<��$=J��HM==�G1< ?s=#� �8,�<�K;V��;n8Z�W�ܼ�7�4dN=Jz<��.������A�5{<�Zݼ�<��7�D�;���Q^��Q=�So��{+=2=�<�]f�jH�}�G=��켩�s��U�H�����w=rb:����=��� =^=et=��8=	l���<�<�<<�E<ޫ7����j�<X4X;��<O��<m�6��>8< �H=ɨ����ɼ�&g=����=(�;:��=�q*��D~<%�ǻ���<<~�k=Ʈ���>��=L<����jH=��G;o"��*�:^�.�&=��!=ΜB<1����&��ܮ�>Z;=�a��7�<_Y=d��<*b�;�,��t#���w���B�E�ټt�<}Q/��	L=�=.��U�F h�3�z(�<zPH=�����!+<�u@=9	��'��f��U��]Ҥ:kׁ���7<q/F=n�;@��{�G=4�;�g�L=uS�E/\<��j<�i]<B\M<mDL=�dU����<F�.�<���8�쐽E�?=����F��Q�%���9=��-=oE!= N="\3=Z�'��&�������<S�6=p7���;)����$�������R=�؍���E<[>=R�2=�u�;I�<��w<4dZ=I�J=|�r��< �lfT��Y[=7/=BS���Q�u	n<
�ڼ��x��1X=���=Fb4�y@�<������<~��;J=9��;b������+=��=\fi���<����"=�h���%<t�:��|;�<���G$����D=D���=.8=�������Z�<�$C��\1��~j=�k���=0E=j����ǼߙE=�6�~yb=L��@��<;=N!!=}��$�~���e=�ҼttT=~�(��oD;}��G�=�(���漡�=�O�=~�ͼ��"���]=�Hp=�Q�A)�������<d4I�˔/= �<���j�6=h�b=d��<E 0=1��ռN=��A�f�'�x��; �"ݸ�ys�<��<�-��67�<��@���B��G+��B�<e�5=��8<��U�ci�3E!=;�;��=�_M9���=�d����c=j�U��μ� X==*$=�����S��fW=�[�6$�<���<��+���=˞����r�?O8���=ԇԻ�G�<1�-��N��V<=�X;85H=Ɲ:�+�C;�9�<��;� �.<���H�d����<��U=Y�<��2=^�<ݵ�<��;��=��=$��<��㺓j!;�=;A��gOt=VLn<��X=t9�;�_P=�O�<�|���t;�
=��O�"���V<��.=r_��qU<���<W`�ti��m�$�*�=�Rq��sf��\/�m�<NZ�<�h=m
a��a;���;�R��
g��I~<|���o�<l��XR=*�V~�<r��.%����<p�=w�'=WW=�g�<��[���<��X������ �m�(�y�.=��%���=�>��c��<���<y3=��X�fu;������p<cvJ=St;ك��������=�������r3������߉Z==��_:dټ�/	�B�=�(��l'�w�k��=z�=�~<���T�v=����qخ<�F���#���<`�<�pD=;^�m�S���/��;��=�gR=��=�6�k�r�-k�]x��#�<�����h�4U��v輢��yּ⯼��<=�����P<�߃�wE=�d#<3+��j��r��������^�<�W&��>꼋�_=�C_<f~<���������6��V�ϼ�;=�*���Q=���;k����<�3�!�N���^���)��n��UU�<
�O=�҄�* �<���<�<#&<kGT��~1��@�z
8=���S�����7�<,�=9���#�<P��;T)=v� ��^��+�I=B
\;��=��F�Rׁ<��8���^�==Q�l<ԇ =R7=��g=&�J�E=��<]�߼`��<%�<�6=�4�<^W=&���*f�����;�켉���޼{X�I�%<^���_�%=��=f�;�ߛ�%�;2�:=��C�O���>m������+����4��Gۼi�=�2���\�9�=1`�:>#Y=V�5���ۼ�	=t(�;�ٔ��B7=���<�+(��L><)wZ=��1��=\�=ea=r�Z��t�;�y=�<�<S ��3=����&�<J��;"/�"S��O{��ý���;J�:��:�<�#>�N=|c�<��<�F���a.�}��|H=�hP=�S	=�=�<��&�h�=I[�<�C;�nƱ��+��NsƼ;����c=�&N=	N��)J<-�*=ۛM9\
�̜�9^�S�@�\�!���,=���<��<9KM�z��<P0(��X<��B=��3=�I<#�r<[���ϸ=6h�h��<�+�<���<Gl<�rq=FD�<W�t�X�2&�I��<�
��d�W���a= ����+A��%���<B��n�	�lh.<��7��ͼ!:�l���u<�qH�Gvx<ċ��mh ��	<z�T,=��C=��$=�]�;��d��n3=:P?��b��_< [#��L=3nD��DR=Ȱ�vE���������;��λ�/^<g ��c�F=Ƽ�<[��<�O���B��_�<e./=i� �D��<+��<���<""l:f�v<�Ѿ��_�;�Q ��K=�6C=�Z?�|�2�|�k��a=	�`��#x=����9ĝ���1𔽈�<��"g����T=|Y^����<u;W�9��3%=Q=��;��{�Z�F��i;ە��yռ��=uJ<<Z�;-�C:4e�<h�"������ɲ��j= ْ����<{�Ӽi�;=����lh�F�@=�G�<J�C<,�<����"m���0�+6P=:t�<ŗ�<�	��ث=\��<�=�<X0c<�m�,�;=*,����LsP=8�8�U��<
~��tۼ�;fD��ځ�{�;�̱<�򽼅����R2��Q;SĄ���f�����!=��W;�'N=���;�<�<�_�<�Z|=�ǉ�лb����=�y4�����C��<�z�=��㼭c+=�%;zW�=K=D��b�==��]<�׿;���<@�<�����}=c?,���.��I#��<�e�<g|<�;�<��f<�+�<k�0�;�<�Jd�),6�;Ar���&;sB=�:^=1�W�/���+=��;9O!<m�]�*�,ER��nQ;L�组2��|w����~�:��h$����)jλ6��Q= O�	���Q>󼝓-��w[�Ł��`�Z��(��e�=R��/��� �;��,�� ��Fo��!=K�A���&=ַZ��	�={-s<���<�*Z=�i�������9��=�V�AH<�H�A��g�<<~�D��a�<��=.�o�{��<x�U=��V��P�=�v=��3�t�5=���8�����ּ��)=xQ=���<@��<�Y�A
m�e�l:��=������<��=�2�1�Q&��u���<�=Ż��<�мF��<g<�?�4<(��<}�P�7��w=h7�<�8�;�as=:�W=W�9�V�=f�;� >�f���a�C=�����<����������<���<�R=�� �����;�"��ͨ���d=E����=�El���m�8�[��%w=�{ �Yw	�p�H=B�����;��y�\μ�2=b�X�NO�_D=�B�<�[,�4�=����!�]�T=�C��E��	�Or�`�/���n��!�]�K�c+����=�j<�=�(���A�<g~�<H�E=y!F;��R=����̣3=�`}=��ɼSȏ<ʍH<�n=ț�<WS��n��<į�q-�=Sf�����6�����:!F=P��q�;�w�<�o������={��<�æ<�^�<��Q<���;�3��܍<q�U=�7���c�{E��_üN	��t�d"�<�;5=�w[��f=��t=����l��<j�2=;��<��=i,_�򭉼��R�bC�<貼�,�<�-=���;�뎼�4=a�弄x6�ѳ$��J��Y�[��N��=i<�B=��=�M�<$�����a�V+=r!�<]�;�l�r�j<!v|<[���S���N=\j=k6W=y�<�a�%ڡ<�Y=&=?��o�k��"��~�Ƽ�m��-6=�3�;G�s:� ;��,=���=Fz&��@�=�h;�a�<"�H���<�@뺧<[ż?a�<��=�b)�˼D��<>`+��X���	�hr=�|=
׆���=P����������U#=�oA��J=)���	=D0/=#��=O�F������y<=:dK=-�?=�LR��k�<�d=�𫺿 =]�<rJ_=�ܕ��p=(�y�g�%��J2�?��<�B<�r�.m�<ӡ�<��<�\a�_�<�<Āp=x !�ކ"�:�M<IS�į%���:��5��I=��n=�F��0�z<=�f�.߻�<G���<R}�;dX
�q��<K�3<�����o����9��y�<��8��i����<�'W=Z�g=��u=T�b=dCM����l*<t�L=y�;��;3Qr��r*=ô�=ː=��;=f�®�<���sa=PhP�MW��a�l=���0)J���x��	�<,��&��<і�<�l;͎�0}��C��<*]L�UE<@���qL=���<%��<���1�=B�^=$���d��;���:��<�C�<�H����&=�4���n<9��;\ִ�+=--F<[�W� M&�v�~<��<�.����<L�g=��g=�%=!�g=�.��b�;r�\<t�D��|#=0�0=r����2>=V�9=2�Z<F�E<���<�=�w�p
<A+��<f0��>=.[==��^=C,��Gz�$-�������������|U�<D���JǱ�3�c=��(��<-9�����</X �T����U���!m=�=B^� �<[<�{�����狟<.� ��|l�T	 =ɏ*=�b�L?	=��=Q=E(��u\�;��;�5b���=�q�bk=(=d����=�ߴ�5=9u���l%���<1]�<�Q==�l�<\8�=*Q='�*;�=_�/��eM����Z���6:��G=���<�3H==G=\XR�<�<9D<Φ�91+/�IG�<�<�켈�Ҽ�=V�
<�JQ<�.}<n�<H�B=WB�ъ��j�<Z�$��(ܺb��!�</�C=b7��@���{��`��
=�$���<�!w=��=\1o��F=��<���:�2=[�9<tj=�=I<���
��<;7=ҋ�X��<�<_��8�<��<�야��;/nY���+=.ռt/y=��O�{��2�6�bt)���<��߼P�W;4%���T�P�<l�G�b�<��%=lH��ky���;ۖc=��黆"I;�0u=*bR��c=a�>=��)=�#>=d��<�<�d�}e+=/)����O=�r�Rh�<F �<�	�;��8:�$=I�D$��o<E�H���<ne=���<*�=�m�<"�껳���+�a=8$���6Ѻ��;ߞ�<( �<&d�<�P�<�k7��ڻ�E�W�0=T�~=��=��;	:h8Q����<��i��?�;!yC=�U
<LW1���J=ʯ�<�|��J����j=!Ҽ̺ ��
��H�<�m�:�=��<�M�X�=�+M�-4�<%g ���6=�w���ώ��B��LI=��+=0F=�"�֜�;�Yt;40��lk=.[=,N=�s��lB��F�;�:k<�s���d�<��	?A=�	=���<O
�<9u���V�Bx�l<�kD1=�7P�bg�<L�N=j\�;i�ѻ�5<��O�C�=M��/(��bD���Z=Ŏ�<�H��K@<�Jk;��W;�@�<��+��12=~�S;�'
�K���fA=�����Bmz=S]G=uw�<�T= =�s}<�����E>=��P��F޼n�˼=y�<=����ɯ;�&���)=��A�=~��3S
�F��<�7=�5���Af=�rG����<�w=���K�<=�7=jz
;I����Y�+=��<�4�l=Z#2��2�<��s�Ln-<0+<�{���9+<�~=z���𮋼�ʨ<�;��G=]I=	{�Bh3=Td�<oB$�$%=�aWʻ���!�e1;=��K=Ƌ�u��a^=z�؇�+C=�3=��G�g=��%=ꭷ<�lE=N�ܻ�l=ϛ,=j{�<��h�a�;��p��_ ���c��k<Tư<��<�1��<-���pϻG�<�f���]=E�<ca�S_l=�[=��Y�>���YP<2`J=�\�$�A=�!�<=A�NIC;���_݂�8�=~=����GZp=�/5=�~C=<%=�K�;�I�<���:�Y=<�a��ց��d���1�<��2<ՅF=j�D�=6C=�u��� =�����<�=�8y���?�˾�@^-=ԩݼ�◽��f�X�d�{�<��K<���;��@����חn;���������=��
=Y��<��"=r�F=�k�<�`_��=�,@=uM=Y�]�=���G�Ժi����p�d�����<�,����;�2%��f'�n"�;&z»�5W�fW#�`�
��և=JV=��<��3����<��>��,=��=� ��O�<�'�;qf�<n<y`�V��$��<|=:.N���l�8R��>=���t���6��<�5'=�wV���4=���<1�<@��<�PT���<;��q�<�r= ��$��rW�7m=3A=��_=&j�;��"��Q
;-�#�|V8���{=�>��-=6-��X���i�=!����O=��S����mW=�=N��<~�k<>=��v��0|�8H�=KQ���=Uiټ?��?ţ;��e=�u�a{<�u�<�< �B]���=Bޓ<��*�����k�:�yc�I��v1(�;�\��y�<�N�<^~#�Í!=�^=o�0�����bĻT;����0=�{���\<~U=}��������<��B��v=%�M=�/=�"�Sͫ<����#K=5���^t=of��i��<�r���p�nU�<�1�9d=�<�
»��<C�6=P2�:���鱃=CT�\N�<�_((=H䋼�S?<_��;��U�3�V���<�h�<^��H-=�����
=�%�;�xR=��伷x���h"=i0~�B"4�`g=j�C=������^=���<�]z=�%=
�����:�v���-���H��+;�$Z��f<`C��L<�BƬ��̼�=�?�=�i��Hּ����<�2=�N+=�J�:׭><@�R�� ��S�;��ʻUd��㰋= �6�V��ۗ<�)�ἳ�=i�<T8��*/����]=M�tá�5�����<����ļ�3�<M%���=�r=��C=�^]<H6��0҉�k�S=qCT��9q� �M��� �w��9�4�<��+=�;= ��<�oF��+ܺM�=h==ጼ�f�;)-�������Q9=�D껐1ǻ%g���<��0�W{���{�u������)�����i���<��=&º2F���^<T2=��<�/4=�;�:�<�qS=�j=$!(�R=?�1<䝔<u�<g<��==i����&�;k���}6=]t�;'1=\�L��^</=�7;�s��<�j-�q�<���:�j�H"]�V'=��;�P=��=��=u��'=�#�1�K����ּV�l<c�<켦���a��.=�y�2%=���<�P��`�x=M �<m�<+軷d�5|�<��0�l�ݻ판����Dl\�`<�<�����ջ�'~=W!�~Yü�7Y��|Ƽ�M��J�<��W��;h��U��S��������q<~�ha���v;��F8=�c���+K=���<^�>��=>=~�<�U�;Vť�N�=|�t��T��L��g��([x�Uٸ�S*U; [/;��N��»e�hI=�=8\����O=(��=���<��$�0�<�L<�l<��I�[�/=��p���1=�Ѻ���;Mi:�AT)=�b�����<쎶<t8=�<`��"��`ȍ<�+�j3==���b��qa=�ޥ�Y�4�Wn�=\�+�R4~=���<��G<�>�q�;�D7���_��!=V�-�X�u�X�1���Z=�J=���[0=��5�g�F4�<��=ty"�94j<�F=H[�<�^�w����9m/�<T	ԼH�_<���<��a� ��X�<VB��-��A�]��"��@7�͈=td.=Ѐ�K��<`a��*3���8=�C ��悼[�=��-=��<�/b�ٿ��������8��v􄽞P�^�.=)��<�M���t=��=�p׼�`���q�s\�<j���PW==Y��󐠼��j=h�k�j�߼J�M��d�yC�<F�<�ak��A=�]��=���7�θM]i��G�����&@=�r`9@T�;����@#��]���|=�ۼ'��^V&=�!W�M��d9*=����0����|l=Be=ul������%=iq�;.\&��r_�-��R*5;mɪ���<- =�e�<j@S��
<���<�Ak����<�jE�'��;�Aϻ�#̼ׅ<��b�UXR=Q��<T�ٖ��^U=�F<�^�<7���
�;=��=+�¦=l�9=��;���  =�W=&U�ٻm��=l[=5(�;�b=K�P�&�e<��=��V=�xP���'������� =Г�<����;���<���:l	D=$u�<M�<l1=T׸�F��������]�<��9�)�����q'=����[X=y�����=/�ﻢ�;�"�_=�%,�����O�<J�*;O���=C�=��ȼ\⭼.{i<�ڵ<؈4�lJ5�q�0�:���&4=�l�<���<��;��=�<�{�n�P���<���<����bG�U�M=�UD9̭G=6�d�.  =1�h��V���v=��D=�c)=~���?��K��XvK��R9<t*����_�[=g2�<����w-=��<?�E={b�;=𺟪����<NN�:�.=x d=؃9=2�Y��7��<j6\=�6?=FU��ND�CQa��7=�S==Z\M=��<�*�3�[��7��W���=z%f=�<;=4����^=��E�����=L�;�5��e��lT
=uE�<�q����'=�F�a>H��<2<k2==t��Z�[�^��EK=��<P&��>������q�0��<�;��:c�&�T~C�W�=T�#=z}<���+��N|=����+*�>c�<Nө;�~��e/=�|#=M�X��=����0=��c=�i_���)<�'7��z7�k��W�I���;��i:�J+<ig �|m��Ƒ�A�H��_仈j=��<_�<
�=�3=��A��-�_��<�]�<b.U��H=	��;i�Q=>��]WH�L =Bj7=Fּ�-=RG4=5L������47��&�=\�Ҽ�$=��t<�-R=�Z=�R?=�=�<�(=��j=�$s<���<�QD�J��5x��RH<��<Q/;��W�;�|Y=T��<\����d=�0�<��D<E�=�B���[R4����</�{<�M=��i��� =!�;ֿ��<:�ʼy� ��T
=$�� �S�̞(<� ��k	�5Y=`�u= �O���<.>;�")�;�/9=lb���;�<��#�;Ԏ�����q����;5��٩�<�e=V�'���<��9�'=eA�<��;4l$=fO��Do=1)<�](=��	=S׺�����m�$=�{-��~}��6��{I��@L��9�<�UT;�9=�8�:�ڼ<���A��x{�=ѫ�:��:<=9P<S�Q;͘(=?�-f�<�8+=h�f�p�<2�\���<��<
�Ø(=U"b�Mv�<Q���8L���<��'��| ��������<X�K<�⟻c�$=�`G�Tf���[��
6����Jn%=�=���<E�<�]J��� 9+=Y�̼�z��ְ���=�#S��4��%Ӹ<q����DF����5�E=o=kc�2��<��;�����$��;缍�T=_�3=N���j=?=��z�[j5���<h�T=t]=v�J=a�:=����=n0�"'u<`� ;�<v$i=�b =	ɽ�%��<�(;3��<�z�<���<Nj��z���6�ɼs���3j��5u��$�<��ټ�����u)��"ƼC/�:�2ļDY�!=
5};5N��B @�ә�=FgL���1=׎�;�P�<�5X=�Z_���:Ra<��u�f*0��`�x^-��}��mټ��C=h`�<��+=�<K�l=k!V���(=m+;e��<�4��aN=�2�S̯��*��J�9K���Բ��e�?���6<ч{<)��X�\=M{��4����v#A��h�<A
C�8y�g��5b�����v
�5����K�3��=4&��9)��=�;�<[��<�<,��P=l A<e�t�z�<��1=q�":d��r�:�z=����=���<.�S=
ч<���Sy<ry��Lȼ�*F=��7�ky"=�=:��?=�A9����<�
�<�U=q4��h���B��5�t=�
����=��L=���<Ȓ��W�;�L��*Q��Ƚ:� ��� ,�+��<f@s;��:=7�i�	�4��7�;l%/������=9�򐼻�d���<oh��C[<G��B���:1H�<�l]<O�&�d=�)	�@�3�������=�*��)�<	�G=��6=�M�/��r/=�鼣=�8��l^<�E=+�����⼽��<��h�U�;0��<�J=%��;[|q���};q;=�V<��!��Z;����<�,�N7=�1�<P�Q�\UQ�Ǌ�9� �o�;�<E(S��ڥ;:�=���  �aP�<��==v�{;B17=�H��ֹ<�"�"�O=��E�!�U����,,>��Ro<b�<��BC8=��}=}�I=����;�����<7Ó�����ڐ;؇��Ӏ<_cP���< �(���A��G�KU�<�恼�z����=\��<i�2�������<n�]=a�:3��
�u�x	�I�l��i�<���(��]9< �J�Z���0����H�/�OH��n�<u+=~�j;��
��Y%=���<=�v=��Ƽ��;��w�^%���T�(=O��<�k1=9�Z����<|o�;w�?��I\�sS&<�1�ٓ<i唼&�<%�C�:��m�򻭐3�P�Լ\eԻGJ̼k&�:(=�������\�.��QU=Q��2)��2�4�a����r���&�<�Ŧ<���HZ=2�q<'I�;X��<m�C=��pڼ���<\7=��h<�6<W`%���R=0V��08=�Iݼ�q˼H��3��<˄��=&�}����-�;jv�� �m=}�)<����<�<_s��~���D�LV��u=4�G<���=Nzq=|y��-ټے(=���<w���!���:<���i��;�.`���<HOG���:=m�<�d=��<a!B=֘0=^=<��3=����ET=_�5�g�==u�8��m=���.���� ��=��~ �<�L�<C��<->=��K��/W<���<�Pϼ����1����A	�<�<�I=��/�3�	Hn<�^��m3I��D=g��;E�=�����S:=� =�,�;���:x�Y� <2�f=R7�;=NY=�1��ߦ<��&<KK)�܉�<��6=�I� 3���>;Q�<?���#�<��f���=1��O:������aq;�,�<�r�<*�|�:�"6�6^�<�E���;؜�<�?=o�3��#�V�=;c���Y���E=�ﭻ[�❉<"�F�^�7<�˜���=��o���z�;ixü��U�2=�����A)��O7=�UﻎA%=��'[<�"< (���j�&��֩5= �
=bF=�<;�P}�i-���3=���:@��<G�$=���>K�;��V���2�x�=�;r�⮼½-;��i������6=١g���&�&�<,��<1@oU�/�}��D=;tʼ��Ѻ>���'�W���=��<�3�;�,>:d�<�x(:;#��ӌ����<���e����}<��/�'4��Rq=�Ȅ=l��<���?"ּ��<��<�(���jI;����f�&=�7�g�$����<[�!=�1"=�y��D�<���KA��<��;���n=�����g�<��<Zll���ŻXyg=WC��̼i�s����<Z��&�n�HQ=���H<6=R]��ɇ<�n��*�=D7���;JS�<���;HN(��P=Ɍe�o\y=
d</��OZ�:�W=�s[��=�L߻L����� =j]�<hѭ�;PK<zy��D�/���5��H���H=�mf�:�V=��:�B=��U��f���B���_���<��<?'��hw�<ā�$==xT��G,�<�|����7�C���Ac~<}:`�\=j_м.c�<��I:>�/��L��6L�<��¼\g�]#:�'<���=h�,�o�λ�p��3�CD$=\ڷ<~.`�r�#=�����?=��\��G=��<�>W<�c�:B;<�<[���"=4���y��d�O��ˁ=�^;��&�{�u%=j>5;�X��)��P=1Z�;�5:=Bo�*��<0���q%A<u��U�L�N�o<	�=�>��B�#�=]<�,Ҽo�-=��X��D=�9�82̼��!s =u3$=�EH=��x<�2�Ꭶ���<~���ݳ<�z=��3�~���tC<Ug�d�=q�4�������j�<<�ؼB�<[�k=�t���X�t�k<�ż�O�=A<�P����W���<��=��=�AG=�s��̘x=H�#<c(�r&=�)����=b�H= 2��2G������Hc=�� =,F�\�O�sF��6LT=�l�<�Z�m=2�D�=���L�G���#�#=���cz=��6���J=�D#����<��<��S=��x�:�7:��;� =��x<w���J��Њ��\=��U�*=�/c=�ԃ;��2=M�"=r�%<�5=R�=����H=`=�,�<�f,=;Ln�2����}��$�<�R�"L��=</k����=�YӼ�α�s�����<+��Gn��������oTi�754�[7���+��H>� v����A�G�1=��<��?�_�̻ ������8=���<�EF��"�;�G-<��=l%�?�/=j}��=s�<�8��ۼ��9�{�X<1�1�}*���A��D�:�;=?�����#�c�^=S?��� <r�=4Cf��#�t�Q<\�?=���,�1��du<�ϗ=��==��U�n!�<m�K���P�u��YZ[=np���F���G=�ut��#M��M/=��.<:_�<��<}Y����:8�F,.=gR<��L=�-=ӇB;�a<���b�=� ��
�;.��<�[��G�<�m���;=����=e=Z��K���:<!:=�<0�NbR=�d/�/� <�O=$���l4f�����<�Y,<�O=
ZA�]!=@�#<>��<���<�� ��β���/;���;+�)=X�j����	��ˌ�bD2<��|��G��:����W�d3��Ơ��z�;�p�<��<o�����_=�1�gG<�d<޹�<X��;�<x ��ވ;��S�vPO=�<��K���=�	��8��/)<m�V=�=��������<9H=H�O�<�09=.�<�%���!=*A
=� v=V���+D������<�P=�eS=��;�����<fmV�L}E=�(=L�z!�<�[�;c�bc=�V>�䝓<��)���?=SH�<Ye<��'�x�L���p�N;N��L�CD|=I=<4e-=li���v�sC�2�S=2��v�;Ӫg��!s<˻ʼ�F����<����c�s�i�w=j�u������*==���;J��FZ˼�?�?�D=�c=�S.�.��;�@�nx;|�_=�#*�1�K�����=+�3�#&�<��ļ��U�K�)��8��g'�<]�]�!E=)�g��N/��S#=�~<jc�<��<�K0=���<���<��=��=<��U�2�D�\��o!=�R��µM������<��S;���TQ��G�Q,(��L=ܲ@=U}=z��=��h=a"�<�L<�r9=����r;����"��E伴䦼�1�;^��<1�мQ�:;�b�
��I�����<��<�-=�N=G�a=�R�-KB=V:s=c��<��<H�`�M�6=��-;�hY=t����]B=�A�<'/Q;,�+=y�����:p�����<�[�a����;���=77��׵K�-�=���<E�=�'l< x�<��/��PZ�v+X�Z�c=���<]�W<�+�<D!E�l�̺��c=��1�R=��:ִh=]���n���0�aM=��4<���<��B�ձ��+���ݰ;��)�OO����(7 =��x]E�ha�#��<q�#=-�H=�D���:�|�c�@�l=�-����i�� ���<{Ƿ<V|;պv��?˻���<��1<�~Q=w��;�(ռV_t��;�<��9<����F=i��:�4=b��<����S|=#�ͺ�i�q�S<��6�_��<�t<Нa��'���.<�3$�xZ��<��?�5	�;���=��[�fv1=�*�:�/=j��<�/���=�>6��4=�u	=A�Ѽ�W���â�wҿ��g=h� �Wf����M�+�<sy=�͛<ղN=:F=�34�� ���� :*�J�9��<|�6=-4=I�<T&켡u,=�ݸ<�M =�*6��7�=i�i�ɥ�<eC׼����X�3��<$��<���	y=:(ʼ�G����=��s<�=#?=�w� ��
.{��_⼅��;��<�Rv;#+?<���<����<0/�f�U�D�]'x��4�^=�<r]�9MOw���i<ִO��z ��X=�i;�6G<�.=-=�;��(<
�=�� =mQ��ż<ɼ#����i=�$��7<L���}�<���#���
�i�;���<ݽ�c�v��e���1�Cg/��s�<C ʼW��yMe<+��Z�<��;� ]����:8�=��d=C��;w=v�L��e���#@����;�-��Vy�҈�<�`�<�=���X=��9����<�m<���s<�o[�;}��&��=q��<wڼ�,�<�z@<���?]Ҽ*�켪"�<1/�<b7���,=��M�6�x�a_�<0�U<������<�Gs�z�����J=��X=�j�4�`���ļNf^<�ݻ�f=��y=��D���<�3=�K�<&G��c[��CY<_���^d#<�+0��V�Ԍ=ce�:s9��pһ�/=
�0�z;�s����g��Ϟ��37=��#=��=K�L���<>�;%��;�m�K�^�D��;����:�:Jx<L^=�Y��)�ټ�ۖ<�|�<�	�m\=u��S�=�#?�4��r�,=R�c��E�y7�=�� =,G��[�<�#�<©���j=e�<�4Y��~�<��=���^��<�k���T���D�K��=0��;Ά<h\p=2�?��<r;�T[�'*�:g� =$�X��6<�Gм[����� ��Q=�*F=�%<�;�<�%"���=���A=��<j<b6N����<!�Լs=��<��J=C[=��;N�߼�������B���L�%�&_=���\���<��<v5!;ll=�r�9Is�<x�.��C�$�7=��<S =��g��v��j;X�ٻ���<��G<{Q<��^=��=�V�K\���ul:$4)=J���`B�<a9μ�[=����YC���â�
�5=e6 �b�=o�i<%ߓ����<�J�< �H���m=*L=������u= �i=d�t_;A(=/Ac�E#��ݐ<*iU;R'R=�?�<y�( =+�Y��)�=��=?rn=A����n<`�<3�D�M��<|\�;&��@=9���<��y=�=�׼��2&��r6=��L=� &�-�t<f�z�w4=�]�;�6=����8U�:��N;|��?�<�2N<q���4����=�#�ڻ�~�;��-=m8軮�5=�4C=�(c�w��/C&=�`����C��AG�Y�/�}YJ=<}F�4^q���U=r���ἱ�N=9`D��ty;�#r<�4��iu<���<��A���<���:�Y<\�$�=�D�`�<>�;i��;\��<��h=�<,
s����h�n���<����0z�4�:�N�<�2<����%J���;Z? =�f=�����j=s8<�=��F����i���:)�<�-�/�<��F=ƈڼ�%<x8i��;�|P=s��<7��<tE[;��߼��;�|�<l��<�| �)n��}=j�%=5#Q=UD^��bu����W� ���<�r�=�FG��B�����@�<���'1E�5^�<�Cg�j�B�{<<[�)����jg�<Xq-=��9=�MX�J�<*� <�4�;4-V��hZ�$�<�霹t��ONT�H(�<�.��F1�<H4�<�ˤ=���;h-�=��Ӑ����<8�J=���;*��x=�-�;�8*�� ���|0;^)A�a[T="2C=a�=���*=�F����<���<1R|����<pM�V,�L[�����n�<���<p:=qZt=M����P�L=��d=�%B���=�=��<����	-=�J˼��<$�;V����<wJ�<|��z^=zHj=��V;��j��GI���+<D!�o�2=�Ɯ<9���<'=�_=;��"V>=N=2��8���N��:
=��<F�<:�=(;�`�<��<?�=��=���C�ȼ���=��rrx=�@��2a��ȹ����=��Bw=�M#==�*�<��<ݼ='9�<ft�Z z����=�<ZK=�YO����;j'C��3���E=��J8�Ht<t�'=�3=����'�6�"�:=|)G��=S=Bfv=W�+=�=r��X��8�<'X�Xɮ��R-=�+ܼ(��<��[=�{\�|2�<��@=XC����d�HE���u<F��Q:��h)�<+3K���L=�cb<�d]<��*=�[�k7Z�����ǐ���I�+�$<,=A
D�Z^=������<N�7�~!Z=\��zK��}:9m�<�G�������������#�<��Y=f��<)�=�ˉ<&�/=��W;]ڼMF5�-�=H7=��+=.瀽av><�-����U�� =,�r�J=���:�u'��D2����& ��X��A
=Ư�<�=�0<4�k<�'<�={&L��|�<������C��5��؂<j� = |�<d�<d3ջo&<u��<W8=̡�< fZ=�j�<_���5=�D=��[�I=V�O���=��J=,]�<Ț=�xq��l��^�9�����(��@�ü���<.�V�Q͚�`�g<��d��wJ��l�<�����Ff�$�\�<N~=��F=��;m�+)�2�!;��K�.�<�)�<�me�ԅ@��d���<v=��;J�h�Qm(<� 3=H"�<y̅<M�O�*�ۼvLݼ,
伃{ι
*=a�<��<�Q�<�Z:�ƙ���Wu�����<��¼����xw=���<��������;p=�>=TBR�.Y/=��C��B.����<��m�"�.~H=��=�/��̧�۳y�����c�<[-!��aS��&���"=/��<�P���-A=�k����<�{;_�t<ZV�<��<M�*=�v�<(�X=9�ֻt�d�V��<M+=�+�-��<2�ݼ�C�EA�F�q=���<��='�<iw-=|K;�\���b�<�X�@L��q<=�WS���=�i��+�/���ĻJN`���=9k�NcE;�oL=�JR���==]4Ǽ_�x��,߻��<��n=�7�;*Qd��a�<�.���n<L��<E�ż�t><��Xe�<��3=�E�<)N�=R=}��;��=8�񞟼�=�s$��2*=����!=K�9�0�Rk���	<�_<�"=nS9=MF ���:=�*=07K=j�r�#��8��=o,��3<9 �:J���K�;롖�g�l�*��<^��<	H:��Kl�d�=��F�/Q���=��=���<~�<8b�;�{������ ��f2�}Gz���������	h��q�����<����5�< �z��)��*��$i�=�=0;}�N=�pO=�'�����D����=�-�~<?�<��;��C��/�<j��<�5�<�T��q<l�^�sE�E�;=�ߌ<��:���<M"a��GA�R�N�]�H��W<��H���9��*H��.=�����E=��<�F��xF=}�<h��?��<�P��!��MHD��q����=�������vv*=�J(:�'=ǉ���-=_-/��k��'޼d���Vv-<l:��Ǉ=����m=�9�A�p=��CvL=�]����I=ԍ�;n@���3���2<��e�ׯV<��ג�=�%=]4�<���<��R���U<f�C<c�'<:�<��<�cs{=GJ��>v��W�<���:��<غ,<ؐ���0�<A�&���?�������}���=\;K<�.�<m�l�%?)��J�\��l=7�;,\W��P��'=�����a<:� =��O�ׇ��Z�;,6�;�h4�@h�<��0�X�<��<�E�<h�Q�sP�<KU��|��;���v�<G�;=0r=H�0=�$=1�;>�%��T3=;���><���<��'=��ؼ���<�6���?�FR=�5�Y���a=�!=;W*=j?W��M�<^�<i%k��o}�N�m�󱯼*�3�Ȼ)���=т%�ڊE�{J���J���,<I���
��<���n��;��	�3i|<��W=��;�f*<�p><.b==�x3����@�I�P�s�4EI=~Ry�گ{�U;==>^8;�
B����8=��=<��<�\��AW�H$�������<j2=�֕�	�a=Z���3=�␼3Ѽ0,��ƃ�u���b���]=<
�<:!#=��L�,I3<{�<�D��>�;��׼���<fE������˻5&=�E=��:o	=r��<T��'�=�q�����<�I�����;P =D�����]=�ϼy�I���<?�<��<:����Լb�<X�T=��Z=�rB=>c=Ac輪�:�
'=�h=�up����<||Y=Hkּ�p:=f�ۼ��=�yv<��=`@�HB<�d=)�<�jZ=�72=v]?=b����q=�9=��<d�ؼ���6�=�*=�(�j�=��">=��>�(�<˴�k��<fS�<�K=uǛ���<��;mI��y;g��@i4=lp���ލ�iC�8��K=�{<�^�� �%�VM�3�<jF=:q)=��Q<����\��A�$�&�0.��S�=��!��JQ�/��B[�<?�{�ڗ'�R�	;�u��D#=5�3��{�[;�ϼKn��7�D=��L<ʒ=����< ��<�P=.*�m��<P�:����/E*���<��1�g��<��o�t.>=��==�5I=@=�l&�B=ۼ�������(=��c�{{Ѽ7�;�����2<�9=�#����R<�^L�Dr��*I;�t��d���,<L��<T$=� ��á:��I��F�M9~<��=b�7:$�<:F<�s;�!eA��	o=sY���t�`X`<(���x��g=$bH���
=�!s=��`�+�m�Oh�<<eX;5�g<x����0=G�[=A��f���0X�Z��<+w�<��0='M=�{K���[=~����I<.�M�(���)�G�2�&�k=�j���w=Ic��!M��\F��E�e��< �;���C�;1�<�0
�ʤ<t�<=�7����<�9]<p���BF�n�3�����j=�EB<�$��<s��<�����<S诼��.��y�6��<.>����<e4*���L=������=-3��wl�;�r[<B�Z�T��:]�<Ӯ%=��<��W�ԆU=͎�<W�4=�z�<K�t�ˍ<�F.=��i��:Q����5�����<��I=��ϼ�2g<�Լ�̼��T�}ٌ=�=;1��<t��<�jW����<�8.=���<����c	\;9l�v�$<_�A�\&=#Ѣ<�-g=	�'=׻�:!ɺ�v<F�4��(L�����7��ZQT����<y;�@==�'��=�;d`3<�� ��M=M)�<�+����� � �e=K�;_�#�1��z�n<��<�v�(��<q#
=�='=��c/H<l7�<��<��m=��G�<���+���?>�3U�<���S�=D�����<}�<uD0=Zt=���+XC<ɕ�����w8�&<�9=}t�&�X��6I�7���Ux��I"=�Q�X@�'pU=E�d�K�j�SK=��<=8=,i�<[q=�,м�&=<}�d8����7<��<�!�<t��<P��<�g���Y�4A��t=��k��h=��j=�=�`�<ܘN<���(*<����y��;*�(<�lW=6��m��v4:�!�?<z3	��$<-�X=u� <���<�|+�{�;b<=�
�`=b=�=P#4�9������X</,���G<z�S<w9l��;��p��G�!��L<H��<��,=�����<˚伮\��g�<x9=}��#_�q�X��u�<y\��@�<�ߡ�a;M=��<��=:4=��g=W�,�p�3=*|H�/�� 
�=�I�:˧<�=����=='�<��.=��[=H�=N�8�V,=�� <tz��R�Y<n�b=�Tl�/�D=��I���K<E=^$c=;*����>�~C=�k�
<��,ń;~�#������#��0�;쓏;��z=��=�_G<P�����K���#=u�ͼ�5=�^c���=��<�%p�8�<kaT=NG=4Hg���6=��=E�ż���2F��xv;(^T<�;�:��W�.��4�Sa=+��38=�cļ�[�����V�:<�"K���;=�}�:���*<�R���G���X���>�u�O</�:X/;T+=Ud��鞼)�%��0��z�:��
��d[�>���Q<��C��jT�?+�<y�<=�45<�; =j[<d�=�a<W"E���2=�H��i�<�Ȓ�y��*���s�#%��������*�J�<�����U�<�̧����L�K���T=Y���tw9;��<YFA=_�(=�	f<3�b��Y^=)!�<	�r<�E!=��0����3�\��<62m="�,���ZZ<��<y�����=�;�v�<ȃ9=c�����/�-��<==�x6�azY=��/���<�4�.�̺�'Ļ�=�lQ�YO�<q�$K]��<w�<�+,;�#I;��+�r����$����TY=��<H�:=�4<C6~�O���9��u��O�|�E�Ό� d�t�}<��a�~�E�����<(}B���==���H����Ώ<a�v.<R�=��Z���?=����E<Qd��:�����;d<=���<�=��)=m�
�[9�����<�瀼%:��5�<�Ҳ��眷 ��<W[
�闁:w�=4^ۼ�S,=��<s�@(;H�=�l=��:h�\=|�`=6E<��ɞX�}�!=�:�<���<Rٯ���s;,�5=�T�<�_=B��;�S���*/�<�._<=�WS�)=P]�8��~�ro��:J=0��S䰼�o���-t��� =e��<a�׼�3��TѻO|Ƽ�5=�9=��q���<�W���o=�_�&�{=P4̼��K=6������ԵA=au�r�Ƽ�& ��'�̢=��A =�V�Z�񮘻]��;'==��)<:�=�h=��6�Qq)=b�8=ϰJ��Ch�JM�����+�?��<��-=�N�<Ţp<��B�i���8=]���G�<�<)�0=e�;=�h�	ߪ���<��Tb=�H��.���f�<i䌻�S�I~���л7��;$cA�()J���<B�U�U�8���I=�P9<3�=�	�l��1��{����lcR=]�0�f����%�<|�ݼ�� ��]G=WUc�8�G�~�`�.��;T�C���6���'=/';�60J<汐�F�!� <�	6=��;�ݘ;Yڸ��Xd<0�3=��ټJ�*��4������s?=��&�3�M=G���[Wc��vJ�$x�r� ���b=��N�~�)=�uN�R05=����XS</�<�uO��BZ=tX����=1����<�)D=ݽV=��<M)%<��<�aE=�{��JY@���f���;�� ��������|,=���<��<�O���j<�G�;v:�@Cf�~����I�.�Ϳ�<�?���&=I)=̋f����;�q!�^�A���_��\0��Bʼ����Z=ǫ��<�W=��<����<tË�!�
�')T<����;!<�;�޻4���&�	'=�+�<�f����G=�Z����<$��m}�s=}�D�oZ�0;=��f�}w`���_���M�X�
���<�UV=��~0!=���<�)�<1����]�<�qH�O]E<L?<"7=*�&���9����!�8����<�֮:ǭ�����<�PM�o'6;����=�t��$=�MT��/�<^F��N�<�Ә�ϰ�b �<G��<�C���<i�=~��<D6����<==�M=��=^������<.�=[�A8�T��K&��=��<)N���q<��B���/=o6�;s�ʼ[=�`	=��<���<�o�;�n���}����<�6���M=U#���H�����E�<�jP�AbG�,fr��W���N���<��Z<�	��5��7��<��;�������ў,=�s=;1�<#2��چZ<�P<�i�u�=�*=Su�����<��<��<��=�E���9,<]��=;=���9�ؼ�Eκ�-!�ͿS<Qh=w�л��<��:��G��9W<-W��u�<�ٿ���*=8n���?��/w=P�R=w�W={�~��=��<��P��Uh<�[=	#8=���x��;��C=��E<�oB=ư
<5�Ƽ��l<���z`��B�;]Q$������@�1~?�G'=�C<>�Q�r|��12�<J�:'�Ż\9�K7��l�<P1Q<�4�%��;���<:�ꯠ�h����[=�=���<ދZ<��B�"��;o�<*�<N#<Q�[=�j<e{�<'<༬�9�	�����<˕^=+�;�Sdv�Q��N�<_��<K�;��q�l�2���l��8�����V=7��<�	�g�<�A_;{��9��W��{�<bBj=A�<7&�<��	���\�kHi=��ʼR���4	ܻ �i=�,Ҽ�sO������0y=9Y<A�@���d<=�;��;�'=��^�;�B������t��̼�O�b9&��=�� ;��=̹�<�Q@�[�<�"=��E=�a�=�;=r[=˵Q�B=�d=�8�ߠƼS��=u_�DJ�<�S�<�ʝ�YJ@�� =�#���l��,�a�)���=;��<�Z=XUм��P=/S~=W�<ɵ��>h����;׳E��z���IU�}�;����<��(=�0�<!C�<��ͼ4�Sc� ����5='�;��-=���<c;����=;B�G�]�4]�<�=k�;��:2>A==={��<}�;<�<w�8=xO��$��<�^8<w��@-^���B��� �!˘�� V<��:!-=�n������Î%=��&��cn�G.���Gݼm�<�S��$6�;�4�<�.���9���> b=}��<�}Z���=�J˼�� =ߣ;Ǥ<G�%=�q����;�#9���
�&������кm�����(;ü<�,
�9"D;�Go����<��=;���t��<PL=7�=��J=}�y;�?q�6p�H7=eM
�3�������=����"]��1\��G�;��S�_=�^�0���G�<�`j�.�=��;;��<m-�'<���U;=Y�ļI��V�ļ�q_=y�=��1���<�J=A¼���<Os��Z=��u=�Ar<'�t	�d��:��$��B��Ir=��#=K>_;~�=�e	=o�'�x(��2GF���.=ӆ=�iD=�ʧ;��w=��F�떅��[<R����<�B�<T�:��)��8ܼ6�
=�$�â��1�<wwD�*H���U<ػ	=�W<�q;���<=3�;�S����<Գ�9ӭT��.��|8=���<� �<��c�x��>�Q�4�����j�{b�;������=;�/=Ў��z�ͼ�=x�i<�&=��P=����7�=�yu�<��]�Bg�;�=�Xq9)IX=�EP��Z<ӕ�<���<�g�-����Ю4��/1=-�=X<E�²��b���<���<�Q�A6"����<��;\z��`�(=���<�>�i)���O=gEe=��7=@���)B�<bMU<��=I&�;��-��]���OX<Xa:#bͼ�Di<D=>'7��~/��^�<"\ڼ��5������?�x�d d=x�<s��<�
=\��� ��A=�C��&��.�\�l=�9= i��W
;�-=!K����S䄽�I�&�Y<�<C=]&=�� < �;ӑ5=��S����<��;|�'�\���N�O�v���͋;K$s��4A=�Eh�u?������hБ�%�)=��+=���<x���,�<��/��L�����J= y����=��<�G��m<�w;=��P��Jڼ��ܻ�1j�v�F�I�F��<�=�%1<��(=8�4���<��=п.=+��$�)=���;MP���<l�<w�t����?=P��<�����<��;<�Q�����<W5�;_;.���A��`��޼��!=���x��<�	�aK*=vC=��;��<����(��{
��ј����;g��;�)�7�� ]��eDZ��g�<��'�6�ܻ��;���<q�<�h<��&="Q�=\\�4�˻J��:�
<�"߼6_5�\U�:�%R=@4��Tk�)��<�i=�X-=��<"4g=!��ΊH����<�_��w�<��ܼp\7=
.�-,�L
H�D�<H�a����<��Z���J�Sy=��C�x!��p;�w�F$ =f:�,96�%! <�1t=6T
=��\={�<�!μ��<�-�<�if=5]=�� �j��<�0�1L�?V{�o����ȇ<��<?P���0=��c=}*|=�	�<:���2�i==�s�<�y<�L�=v�;2�9�&�7�a��2l�>֧��B<������X=Ɣ(=}�@=�ބ=��=<�!)�o�N=�"�$��<G&������k�<=��x�z�:Zdż���<(�"<՜,=A�\���Y<�L=7'��3E=
��0��;)�&<L2����H:G=�Ϡ��-T<�߼y~=z��<4��</�=�}��<w���.=�6-�!�=w�4����ЃS�I��>&��hʓ��5`���PPK�l�]=����R_�<��<f4 =	�=�;ټ��$��+�<T��<)L;�ri<�֢������<�\�<��\=?K=����G���;+�k= WX�l!ۼdr=�C=���/8N=.�T1�<��E=�ڊ�4��B����q����;\��+��c�<�Tּ9�<��Q�҆
��q���b;��b�<3;#=�,e�_~�<Y��<�/1��@���ټ���=8:Ս����;��<�^�K�n���<���L�j�(7�Ɖ*=
5?<�-=�S�U�=
�)�"�=Dԧ<~"=Z�L��s�;	>�A����3�<;lS;A�<�
<A�<��ѼrV�<D�@=/�E�[J(��0�j�v<Ό=��ػc�H=M�L<G `���"<9Z���V=ann=�Q��Z=�S[�#���!E=o���sU�<�  ��*����=8Y=�>�;Χ@<��?�����==����<�=����A;s��<�=���1�<��#=���=2�#=�r=��=�F=q�:��a=6=�#8��W���?��}�<�<��<�pK��+=Q��<q��<>�ʼP���W~=
$���zQ��RN=jb<�F>]���	:'�#=�Mk<~�����i������2��r������<?2���=7&�4��<N��}S{<�@�&��;�b"��;��2��T���&*�fP�;$�3=?��<�.N=I�<�.�KC��SE;�Z�O�!=� �<S'����}=N��ʤ=jHx��;g�������A=h-�;�g=�J�i�<e�)<�땼�����S@=A�<����p�=aq2=`�b�`�+=�����<tK�Q�1;����y�����q=q��Y!?��*=����Ab�<(4��뀼R`�<ߨ2=h=W���9�u�༐NV��(��XR=��h=�+���U�i�Yڊ<n��iW-=� м���A�F=�}u<�<:�2<*���<\$o��A�ƶ0��Q=$V)�!����.�h�{���"�2��;]5=k!ϻ�g=�%��Dq=�<Ӝ<�*Y��˅�
�ӻ�*ټX�=�xT�k�Ҽ��!��@��f�f=���<��j=��H�bE�I'�<��b=.T�L�˼k��<p����+$� {�О�=o�=o�=`ג�N�<���;L*l=��L��ʎ�� n<��
���;a�=�Bk��B};��S��d
�^3F�R��7	s��ϼ�޻�ٛ�8!5���ݼ'i�<��#�[�-=�}�<��z��;�7)�!i��X%<2�F=���Fn����e4��"#=;V==�b�2��=A��<B�3�e�?=G�+���9��Bк�e���)=�,&�7,)=�"0��˄�\Ǽ��I��/=�/�'.H=`�=�F=������-<�#������=��W8���e�8�2-!�^�b��~�u<!=�g)��L=rl=��=�=�;�f��.di�@��<��;=��L���<$�����1�����G=|X�<�v<�����L�H�5=��H=%�|e����L=�1a;�'����Nzƺ������2�V��z�Ykl�dt[�_��<�S��K�!���+�?Oi=2Jļ�oN<��;1����Ʈ��Ɉ;}����;》������<�����/�2b7=�U����;�E�����;���j�ƻUCԼ�o̼$�X�S�<W�<@:,���<<DZ)=Ǭ��A=�Ȼ8s"�/A�<Եx�y/�<�=�Hi���=ײ&=��;���;$$μ�ԫ<Bg�;��=���<r/G=.94�a��;L��\Bx<Y�\�����V� �퍜��| ����d����~���=%t9;�����2���<���:p:<��!<�x�<�3�p�
<�.�<�?=��&��>=�C1=�r��<��_���ɼ�_�:Y�'I=��H=Cɼj���<�5�<A�F=g)<�:r<��D�B�<~�L�$&-=B� ���:<�Z/<g���I�<��<��t�걼laӼ�,N���S�o��36f�-�'���3��P=�p=J<�)=�?=CA�G����;(�=�����;�Ӡ������J_�hb8�TJ=?T�:�c=ImX�7�[=0��<��
����<�P�ܷ��*��<��=��	��R�<��<*+��?׸�r��<2?�<A���J��<�7=9�!���==�7=y��De�;��I�}�b<HW:�iA����<)&�1g⼴rV�hd=�)�<��lYo��=�p1�mC�<y�`=�Ҽ�;�=_�Q���C���7���k����7�8;a�:���Y�<�8: d�<�H=��H=2)����<��l��i����H���tc�Cm�<R��<#u@��;�:=�m�	( �ABc<z�#�!ܠ���;(������}��&<c7=Sl�</�l=xx;;��
<8ɼ��Y=����SD;��U<� Q��i�=Ѧ�����;��>�;������s=��=� �<Г��9�=�l==8�:<T����S��^��^�>X�<�|I���1��\9�xE�E�F<�>�'3U�]N�<jZx=��r=�Fx;.��;Xq���;�ݥ�9�n�zo-�N~{�$�J=!=��<��A�ζ]=�y"=���<����C��<��B=�U=��F=x-���;�&�<��<�8f��)=S[l�	͠�L�%=�0=Q�W����<�N=�	=l�M=E;�	1���=�h-=J�;S�#=tU��2닼r����<t�;�j���\�J�%�B\8<�Ƽ?�<��G=��m�`��鵼����D=4k��ge��!:�Y+=4L�3��<8� =������2�>\�HDǼյ�����
�=��_��b$�wZ���?"=�+=F�=mE=�S=����]=9�S���x;r�k<$߻�f�ຎ�7=�Vf�H�Ǽ��=eM�f~K�a���Y<_�<A@�=�����S=-z����]��m��E�=<�d���L<�&7��	�v�
=��ݼ�廅%�;�ٕ����<��q�K�%��y����p=�
�<��¼��A��t=L� �J�c���;Pv������,��F���P=%�R,ؼπ���r=L�U���0�~�	�j�ق!�+��<�������WL3�'�T=�g-�{] ���X��S�;?q�釴: oL�S�+�	�;S�ʼ��_=�屼ǔP=\2��o��|?p=^H\���ɼ�8k����c1ݼ���<�^=�w<U�ɼ��<Fe�q��<::��?.=~�y=u�<�8=;X=Y�;��Hȼ�F<9q��R�i�	�a����s����h9zl�<|J=�-%�+�V�	��<���<��<��P=]�<=��<�?<u�S=Xq=%Fx<ji�<��q��GN�<_��L�?�	����ݻ��"���<�
�<c~���j~���F�B�Y<({�<�=�U�=�y]=�3��r<R�<�pH�ro�;��T=�-<X=�����X;q��S#<�~>�d���;sJ�	v-�7�
=�C=�!�w��<r����˼^��<�\=��߼���:B���>�EP���{��;�Ӌ��������<9��<�o@=�=]I���
��Q�<�Y?�ʆ=-�̼���k��8=�e=�Z�<��U�<�J=�]<[�w=��6=�����<���<(���A�<m4T=(�M=�j�<�W��[E,<`�S�i�-�WTJ=�_:����<����+�<(����l=���<=s&=�T��G��CX=Mo�;�X=� �;x^�t�@=�e�K�+��1=�w=&0<{�=E2N=Ǉ�<�8��p=P�
� ��<���(����"=�.ż"ME=`�<�̡;��D=|x��]B��#�;�2����4�=;˻V�����<�#��gT�<�V�<#�9<Rv;�5N=�F=:�-���8=�[=wk �7�l=��	����<5C����;ld�<&B
�����2�<�[��7=�Z-=v=";�ܠ<��S=��`��i<���<;+���C=�U�kK=�<ἔ�ݼ
+<�!N��X9��%�<`�<��+��&6;��1��MS=���;��#=�����=*ZB��Q�<q�:;��1=P��<ϙ2�m;�<�� =hu+=e��~j�;�Ǽ�Ƽ�����z~<�b"� ��<<���� =+0�9��M�g4�Y�K���1�-�X�`�ӼԳt<�T�e2�<
 *=R��_P<�?=��T��O��C�<3��<�i2��4=�<?��LW=����+�<M�g=:
�<S�=�/�;��<kF=�3!���N��Ѽ�-=�>q�lVL�����*�6=*�o�Ö4�V�<��a�s,�wX��e&�`�0=�Y=m��=Zc��;7׼��C=�u�aU��2�=�<"�=�p�<���<:�Y�����'L5=@���V=��4<Qj�<<�;��9�=�V�<�"/�6�&��-���w="�q����V���]=G9=a'<��}��������t� =�U"�vu���(=�L�<�X =��w<�����=�'��8���_���Y����<l�<��+=��\=�|D��w��)R=LY�-�ns<�\��CDm���<�(�=8�S=�q>��p0�����H<A���	=1��=�yͼaξ�WT};9�ļL���%�$�:=6dB<Ҽ,�`==o�<��	���k<�qS=��4=�����< +�<;n"��+�<i!=�Z��<+I�1�K=���� �[=C��<���^�C������~�JI��o����<�l���=5{�me�<�c��,�<J�<ڑ<4押 �"<2�R=4�=l
���*,,=�,';O����N�7=4S�3��/=��3<�9L=Q�j=4?� a�<��<Fi4�LJ=	$5���<0�M=�&��=FL<4�<��
=�9-=�V0��PV�	_�����:��/�:��h�<)(�7DK:~|	�~�_=b�=n����<���<I�=�a=;�;���<�,<a�.<\��<�OD<4�ܼ_���;��<4CH����<�x�M����k�&F��=hV�;{X=�L <w�<Y�^=�<�)�<X�8���Y=t���
=��O�~�.=��R�����gK�[�O=!:)=h,=�C��Y�<�M�<9���唄=M6���<�*=�=��C�/�;mf�<r��<�i	�F�<�Y�� �<��Z=�,��6=��0�'�]=������=L���$��U�̼OJg��L�<�@k=e���D����;poI=�o����ϻ9,=��A��3�<�AG�r=���FO=H6�U�1�Mj��=��<�%��=�2;=��\=u�����_��oN=�ĳ�w��<�A�f�i<�^%=�}
��ɼ�b�;B�;A�<,G��ge�<�]���u=�r0=�����:��^<Q��<�BE�u��<���� W7��V=0�'�am=V0���>=|LH��<�޷+=�q�=�'=��R���#�eD��΅=�����μH����Bw��K�<��ü=�:�J.=3�<�p(��yp<���<�T�<r-�}��;�=9���<��7<��<Ϗ+���ݺ�2��� ���8��r=<�S=�޼b8���^м��>����<�k�ф��69�[����h*=ۯ=��=��\�3!<�j(=��=�v��k=��@��m�<!�S=~U)�
?=���������
¼��#�/'=T=>�4;;	/����+�M=�p�Sּ�v;��<9�M=7i=H��&;�~�8�~�q��˳u<`�c=�U;��j=���=�`^=r=z�3��$=N�Q=�"=
�@�WI�<�&<]t��3EE=ذ��o$�!y���a><)�(<�?���=X�G=����{n�4X��r;��G='�w�T�<�����/�(�Y=�;=�r�V�/=�x&�z�X����<�cj=�3\�����<���=�Lr<�:�<b��Ä�=�����=�^Y��N��؄��N=�^��s�j<E�ļ��)�{���ge;�����f�>=HB�<�;K��<Gy=->];+�/�0==
���<`�n��?E�C#�;��<>
5��G�<$u8�w���� =A�
=Gg=mz�9^�H=h�¼do=r�/=U�f=O[<Ԭ���U%�C슼�ּ6�&�D<�R����<|ك��L��j�Zlp���;��һ�!�<����	���+켃*s���'�ҫȼ��Q��P�P/�<L�U���; �<���W�;��=�(��Y�=��ջ1`=38^<}@:<�{���h=근^�ѹ�;��==ы��/�v$=_�=�<d<T�I=F��<����
j=qd��\������he=�?<��ͼ��:��;����;|��-¼�z�<D����"<��<j�_�Y���ɢ;si=к���$<tl��Z{�������&tz=/m�M���gI��<*b�ҍ8�T�ʼI��<H�޼B	8=+G5<��N;��ͼ��H<�={�;F.μ(���y�Uo=MF>�55�t </sӻ��<�'=6�"�/҉=
g��=3Rٻ��=6A=��=`8J=z�V��?��,!�=�����������Ǚ<��@�$���g=�H�b_���_=�����G=!�=V������;��N�Y�x�
*�<��<clU<@/�0yd�|�;}���P;GC�<)VL�.�8=@�V�����9��<��3=��=�l�<̳����;�J�o�1=�1�������&�>�h<*��<Q����N�V�H=j��i�$=��?���I=p�K=)�<�ֱ;��S���=�A=v���)Tڼ!���X��;�B���s�<���<�_�<����P�<��<:�+��[�=>fE��|<�9���S��;nҀ��{��:5=�]��Q�8�K�O.��M3=�;=Y/���a=^E&�4��<a�z���G<�*X=����<��<{P�,�=᡼y����[�<��;| ��K����j���9a=FUX��(-=捻Ay�P0*���<�gm=��_�4+=�?)=}��MD�W�z��d��D=1!c;jg\=���<	\�<-��<]��!D=��#=�;ĻN`��'�y<l��K�'��=R��H��PF4�~@&=q{��}�N�ż�/�����g���T`<HCH�H�ɼχ<��`�w/<�c�a഼�Q�|�p�,���֞*��` ��e�<��=���%�)<�1i�[O��Pz��98���<ex�iH9���2,=U�[0��ʩл����8=m1=}�߻������;hsB�5�<�<�ġ:9���_��ƺ��i��=�;=�-S�s�W=�>���<���<�HJ=_Kf;S�s=�{C��ԕ<���<Z�a��_��5����=q��ڴ=U�<=g�P���(�2�<����J��G���L?=�ۼ?$�<M=���m���==2NP=5_�;}If:���	�r;�<
�Y=G�3��+H��#?�5��,*	:��'�n�Ѫ�k�ص^=�#V==�=s�h<�Yq���<��)=�_��u<��Ἃ��>$<=U�L=�I�o�(��$�<#�9=�0=>��I��<�F-�����&</=�4��l:�-H=���<�"<<VF=9����F</���7>=�)�?�����)<A���}t�<�d���(=�%N;S�>=f�;DHH�}O����S�j����z<�K4�F<s�'�n�޾�<��s�-=yq=��;1T�<�=��U�S:�G	�	�y�W�#�A%=Y�⼶����5=����-��U���\��p�Ӽ(����<[L���)���=�F=�24��}_=|�C=�].=�`����^=�a:��;=S8%=�8x=D/=�8l<���RRܼ�X�<޳�<Z�B=5��T�
w=~�<�/>��'�H:�<a����;|j����м�p <��P;3�8=�/;��3���n�z�μhIW=.á<IV�<��<hB��8ɺ�m�<����*���=*��<��n��N�1%=5xJ���><8�H=H�����:l,9���[�r����=�����~�t}n���3;�m=7�,=*�s=�塚!����!�̧O���-�T�V= ��<}Pu;ՁR=�V��R�������[��w�0y���A��"�E����8�|{<kr������<ɖ�<t�t��<;LP.=����<&f��:k�ͼCD�< �����<���;O�ּ<ƒ��3��i!=ЛV=�g<D�(<dA ��m=Q��<b��<;pv=%jk=E�W=1�c=7��<��#=�K�Q/�<O�M=��<,���9�)=Cm=?� =3�=G��<S�=LX�	�ͼcm7�����z�����D��<m\D���=ĳ��&ẗ��<WXU�D�^���N�,�d=��t;p��������!=�G4�	�<%�<	o�r��<BtܼL��<�0�3��<<�9�FM�<Yo=�z޼%���:<���<�1+�W�V<�bP=FG�N"X�:=22p<�� =�4� ��<Z�L�&�Z=20�4M=x�8�$��<�߄<�<��f=�'=wc��0<�=TU=jϼ$�������%�R=u�<|2��a����<&�,=`�1��H<Zǋ<2���$;5Io8��$�C�=R=�`�-J=}�.=eF�:T-��,U=��V�6X��C�~7�<�/q��{/���<f��L�b=�Si�h=;_)���h��1�;�$���<51�EE<��_=�0U��'<���:��*=R�<8�I�8�w=��<Ǹ ���:=�_�ԅ3=�#Y<�\��E�6� !��S�ڻ�XE�?�=H�E��@/�/�8=�:�<G�*=8� =�=α.=g���E��6�<���_y<��S��,<��-=�/�*�<���[ɷ<,I�<��޼�+>=2�=L�X�Rx�E��<'�=������=�
&�uS��F
=��b��5?��Xh=qu��$��5G=��<Ay<���6.��ä������a=T=+F�[Rz��C�3��:<-=¼�l=�*=�?=��m�f5��#�ɔ�W�<t���Z��5��χ:
[W�4�5;�[���`�<�Wչ�{�<�=O9�;4=\+���=(��<Q-�.�3=IO=9��� �s==�j��e=N=>t=�i��c}�-=!��P�<T>�A�"�
Iv<@@��<��ك�Oc@����9q�<��A�>i���J����=��+���$<B�K<lvR�+� �AO>� �i=�P=�o;Σ	�y�C=P�<)?�<ܰ'�A/��A�<�D0��J���*�_o��s1)=
��<�'Z��B��:=Q	]�3�һw�A=�m�B�%=�;��<E�+��~��W(3��e=�����<Sz='�i�{v<�17���7<v-G=�vƼ��=��C=��<"��<���j�5��R��AK�<��'<J��;��<6�j<ƿ�ִ�;&����Ҕ���:<J��SԼ)���+�9�D���𼽒�<U�<}�=�B��%=�=`��<�?�<P�R=�}><���Q�q�\�{���<����T	��
=J�6<�8̼.eC���H=�C\=ǧ���=*�����s<=���X!=�m�;Dk=4�Ƽ��&��r"=7΂��
1�BI��@�<�҃<���<=��k�hF);w�L�Hn=�/<X�i=�S</�<��M=�*s��b�;����!�<`�=2�7=�Z=bO-��b�=�Y<�MA=�LF���E=���<)�����=���;�G(=甇��<I:���E�[4�5H2����<�(_;�@l�{d��^E��]�0=F2=/�1��X����<��4=υ=��t9=;�0�%ؼI�f�^t<�e(;7<��B;�L��%�4��+(=� <�$/��Pb=0!H<��ϼ��j�jS�<�*o����<�^0=��Է�ؗ:VP=+���SY=�Va=:���v7���=E��<��ϻƂl��^	�
���dF��G�<f�ͻ��C�(�=��H�5a��wK��>(����	�>=y�����7�rRx=�-�_�
=^o��8�c=���֔#=�<Q=JU=���qю=����'8�9�-����<%R=O����[�$�/=�P;g\�RGx</l���Ŕ��Xü|�5�a�-�`�� ʻ�c�<!��<"N=��;"y�Y��<��7<�闻Z�b�Z��i����}=w�x<��\�\�3�)��<�L���I=�h1=0�M=�7=d4=+3v=��;7����˻�J�(\�<ϓ�i�����T<��R=��<�>=,�-=�� ;��Q��}�<��9&"�<�� <�Z�=��<)$F<��=�����	E< ��9�o�i�5��9s8*=Os=��<E=9�2�
�#��BĹ�L��y�<�H�<y�v=)�U���D=PG�!�ؼO,���=ˠG�UB=W*�<��i��O��uB��.(=�����;���ᨦ<�1�u{�<ɧa;xeC�D	h=��#h���Q1<\��oT`�<��ND=R^�H<=��6��D7���:�>�'���Y9���oʼ��<���<�=U�t��|7=	Q[=,�Z=%��<O:޼�J=pu����<�.=gz%�@�=��<��<��=򫍼3�c��ܼ9�#��������k=0ϻ�|�<��'=&m�<�\(<~��;���~HO� u1��T)��-a=@� ��s�Q��<gy��d=��`<p�6��F�<{%%=@8=�	�U�/�-F����=E{7=�V�<��<D�ۼ8�<�R_= �a����<Wyr�2$�T9�8�<ە<�d�<
a�<Z��soɼFR�]4=+��<:;�<-�
�1����U+=�F�;�+<��X=����Z'=1p���~�<�g=^��<Y�<�2�<ɛ{<��R;	�=�N=Y�^�i)�����;*�=�լ��=�$6=�<;��2�����)�-=]��4 ������<����;G�<X�<U�=�m==�r���� =%E<�r�9��/���<r��;���;���J�<;�f�ڋ�<M�j�]�0�{�d<K��<��^�!�M��B��S��.��<t=�X7�?�I�0��ˈ<��M��[9��u^<����DC��W=�B�,���cL�t�<����_�*<�$=��O=Ԃ�<��=3�=T���
�^�.���h���<?nW<Ȅ=��@<��=�WG�R4=��;�}=�L��|��蠼,���1a=��W��@= �<�Gg><�w*�/�8�!i=�Bd�U]�<�ۼQF鼽w�<��{<��*=vi6;r-�h��1���	���xD=��<XY=��<(o���ٺy�!=�uۼ��=0OQ���a��"<��<��@��a=��<�z���d=`(Ƽ9P��&0��¤#���v:�MH���n<����W)A=J�8��7��xI<)�!=��a=b���� =�46<�|�<�7��<w,Լ�BR�/aݺ~s��Dd� ]�>��<?�=[�T���!���<���:g\O=���y��<�͎��s=;U�Y��<E*2=��a=�ͼƂ��g�>��3�<[W[<����*=�v=�;�i�<@�<	=�ie��b�@)�>&<�q��C�<~-q��PZ�w���B<^.i=�L=t*=FM�;�

���s����<���Z�=��<�8=�����;"�u:M�I�� H=�=��4<e�=�	�<OH�O&�<��[=&�U<�ǡ<?x�<�����`<J�U=��β=���8�xV==�@S�,�M�����C]�H�3=й'�V�a���<��ϼ�le={K�;�*�gF߸7�<����!=�7�0�,~���G���.<5S��|�=��H=&n+=�'��?><}�=� �;>�W:N[��D=��ü���;_�
=�;#����r<Ej�=������q��2�l�4�汷<�r<�:�<=2=�WՆ�j3�<�
�<�5��ݧ�;GyQ<�?�����gE��[~��S�<	E�,e=x:�<��;�Ý=JU2=x���<���<~��<��<�VD=��J=��B:��<��<�D���.h���<�
z��ʖ=���<\fӼ5l�<�x���]=K�<=gኼ}�i�pu�<dC9����<--U<�x��^�<�H0�=,�E=z�;�Ya��D�<�T+�Oi<�ϒ�(;Q=��<i ��U�<���<g.�`t�1�b=�@#=t+�ަ={�<�3���<�;��Ԯ<�{����������&�<�P~���P=оa���<(=v?<�9�%�=��[� QT�9W��^=&8(�i3�҄S�/&��d:�<�<�#Ѽ���<W=b���Z꯼����U=�d���d���<�%���$;��<����G~�BE`="�<�s'<��4���*��/=k[�<����F��~�ٮ1�H�5��K5��[=ٰʼ�.N��:g�oe<�[A=�х=��G;.���Jt���&�5SB=�U=yvy=���;��]��<&�oB��Z�_�P�+=z�W��
+=n�t���:<��<AB���O�<9zQ�e�߼<�8��X=0m�=������"<3�]�"0a� ��?/=�[�<g8==n���~=��`�V���ɠ���^<t�(=�`7=C�p<�f=�y�*A�l�;)K��3M<�3�B���K;�;�ؓ�&����^�,^���d�$G	�}�μ���kb}=�t��m�Ήy=R*<�k�<�$F���3=\�e�=}W�;E�N�/��;�d�<?���Q=��O�ļQ��R�c?=@���<�<�Q<y�=�����~��w�#@��<J��o>�>�$����;Dt�9N��C^��ޖ;Q?p��c��H!��Ms���+��P��U��<(���e� = �&<DK�!M�<��L=fǼ�r�� �����Cl5���ZZ��Y͂9I�����V=��+����̼��ɼ�=P�-����<�W�; �a=
-=|:^�@Y���$��H�����<r�C=�7�<?1���*<R��<���i��	k�<�(�����P���h<�t��P�68<��@����=�<]�=�Z7=���<e�0=<��GX1=0Xv��0�P�)�}üy�<�Q��5(=�m=�W$=�%M�:6��� T<k�b=��L��!?2=����~=����}+��=���f<Kxm<ByƼ������X=a��;$�4�p0� n<��<��r=�=ĻK�B���d�<��w�;��<l�ֻ��`<G�<�xļ8Oy��TH��x=�z���F=�F\=N;���9�f�=q�9=��6=��H=��%�P�;=���z,I=�׼1��:�C+<�-	���P�V����[#=��E=ՍK=_<}b)���<���q��<֦.<��[����|9�<�ݼ�)[��p��~!<�r0����<��(=/ػC=
�D=�� =�W�7/�����ei=Bռ\: �G'=�������<B�;WP�;$<�Ť<w�M<� =�@<��'<�vL={!_�LW����+���=����P`<��<=��<sR=^�.��a�Q�;�h�\��KJ��׻𞕼M�;z=�B����Z��)=�Ǔ�h�<��J�I��<2�o<��<~�=�&�=x2n����/��q=ëq�~^a=��˻k�����<��s�����-�#/=M������� ������8C�E&A�g����<�' 8=�g�<u���/�'�f�Լ=��<�}���=�p��u<�V=I<!=��
�߱�<!6=o2k=���+�;[^N=@�A=��.��_��A���=�V=�*4=H�A=��:���~>��Q�����@P�<Elw�޹<��R=ăʼ?�<1=��L=��<xNF=<�<�;=�+V�_l��"g�
>��8/����;�9M�`�$�(�=\H<�%�<�p;o�ļh�C=�#漹�.=��o=�_�X��<��+=MYV=)�O<\Tȼǡ�<�欼J�T=�x9�h<�$=�&����Ѽ�0
�>����Vc=��%��h��pa�;c�/�m�I��f=�P�;x[=Lb�<�����ig���<�_��z:��"=�ܻ�:#.=A�d�s-=�1j=�!���F=�%=��=��)=��o<���<�A<=��<Wp����3=_��; �=f��<��s��<M�9��=�"���;�2�<�t=�u/�8l.<�=2i�VX`=�a5=�;��N���=��6=-h�<-@H<��e=`�=��м�͇=Ls7�)����C����@�[@��BZ=��w:�tB�:v=�M�5�W�
�����[���{��mm=*m9�,:W=�I=�Vs<�F�Z��<�a�Y�a���C��JP�o�J�/z��j�<s<dzM=t6���8a�z�<~4=&�%��$=�;R�I��<9�)�
�� JO=�^����X�<�E��w���N�[(`���S�f7=�;]��Qm=�*˻�G�Gs̼U�)�w�=�X=�	�<ζ̼Aֻvb��إ������T�k�b=3p�e[Y��E(�k�6�z��<5�_�\�<����2)<I^@='�a<$?=��
<�����\�;l��=M��<���������<2�w�<��m=m�̻��9�-��;{��g�V��ߐ<u�8=���;�5���(=�h�<�߆;�l�;V.*=���f%<b�!���O���=�J�F�R�s��;��
����<^1мRT��BB= �j��<قC�w=��$�;�bd �����)��L=Ԁ=�<s��=V�,���|'�i��<��+<�c+m��>9����<-6=L�<Ly[��<O�ؼ��=������g�i�U�	��+j�bg�b��=(/߼JAH<O������;=���; ��0����;o[:ħ�<v�X=%��<����FI��-�;��G���X�6����<v<D�@���l�-�n<��9=`�E<%��<ʢ= m�<�K�;W���ӝx����� �9f��b�!-���]��X8=�E༒�ջ�d�ѻ=r3V<�'�<$81�K�t=��<�;4������<j	��y��s�9������0��%=��;#y������k{�<�A�;9�%���߼�?
<���`�=� M��.�==��Wn�1=�C��/�=>� =f�=�R=�(=��i�y�.=���Й	={=��k=n=�<*q����=[+Ǽ#����a�=n�+=�_:�z�<�u^��}���C;�4�<��1�� F;�fG�E=�;#����v,�n�<��W��:a�P���:=|;��]<��p=�'��7�=*˭:����El=R4<m�q� ����j���<(=���<M�m��T�n�<��A=���V)�0q:�)� �fqW���(�'��;v��<n��<Q5=�І=�1<v���A�R�qR̼�.��A��E�$�MT=3��4�$��h;Ǽ9g=o�<o����P=O��;5�j=��.<Vi<�_�<;6I��C<�<=�=���<�.��/Q�n���Y�� ��<����$=�-��U�4=�<~=��[�`<���<����A�j�J�tt�<���<g>=M�#<c����6�D6�<���<���f,=��g������=v�ռ؆�����_�P���4=�O4�n<�'=X���==F����|Ļ1��<�43=�/D��8��5=�ԼY�7��O=�/�E+= ԫ<Aj�<7� �b0�<ךg=$J���S==k8=��[=���紺�7[�%Gݻ,/.�1 ��8'�����Z߼P@7<��-BɼE&Ҽ�=��~�)�����<2t>=��)�"��z\��*���[��<�<>�u=?�=����vn<Jr;��s�s�o��"�<f�9���=��8��g=2�;t8=Ew�:�!�o�]�<��;��=�Ғ=u!=,m��RFp=!$�<s�~<��r;�O<.G�x�<��<�#�<L2�@�V�
̟;@��iD=�2��s%Q����ǉ<���4�<%�A<R�Լ@�G�e!!�}��"�_����=1G�G��h�꼛J�� �=	�<�@u8==�*�<�
=���=�<b�'g��4=2�м�ނ��A;:�U=��:��læ��z7�N8���,�<3$<�rT���.=����f�> =[��<A:=��Z��>��[p�y��,�2AR���>=̈u��{�<ϼ!�����5=R��=!l�� �<�<�<���<P��5�<�I=˘|�%��<w*���i���(=�Y(=�<c�$�K=���63-=����;�m��	�;'���`o:b�<Z;�<9>=�4��wlv=3�`�rj�> R;>��
=���<���"����e8��*~������T=YM�<�M4�{hI��D<=Jp����<4�<g�y<�n�;AM=;:�=�y�����<�R� _���b�?=���<05ǼSUF���<�%:=qŸ;�9H��<[�8i ��=9�`=�lR<2eb����<���� ��~�;�6,=�mx<�v=�K&�Ĩ�=Pq9=�%U���'<��3�RB���g<�C��7Y��`���b'=�\�<ʐP�;��;�����<+|�;��0=�j0=��=K�	�p�:=֑8��/��a���J6=�R�F+e��Ag=��c=h��<��{�
kC=|�C<�jq�37üi�;舊����F�<Y�����}=5Wܼ軇<5X�<�y�/y �*)Y����<7)��V�,��<Uz';��=z��QI=R�»�W{� �@=������;$��<�~=���;�k�<bV��B�i���<��<U��<Ҹ�<����h�5���?=		=6-+=|n4���%���<�9��.�]3p<�x6�Bؼ���èz=���<i����><��<K	=_��<!��<-HA�S6�=a���#�<��};Lҵ�Hld;�1�<@�=i�L�I0=y =]@�:�o=�|��j��ˁ���E=Ѫ��I(=_��;���<��<@���//�<\; �٨G<�=�cU�lo4<���= '=ѹ+<�p,<L ���F��pH�y+%<);�<�)��π	����<�}=�Gi=��i=�K<�v2�	4{�񚼪@���X���A<���	#=�eW�T�5=�4�;"/����!�cB��vL�:�r(���=-�v<�AT<��&<�be�Sͩ��񪼐 �a��:�����<�7<]�)<1�=�|� �:='�Y:�i;�*><�f���P.���T��P
=#=�^&��>�<i+����c=�� ��u<3��.��6�9���<�e���8`G<��<~q�� |�ǔ�<E�V�Uh�<��=�)���̻�e�s�伕�p<�R�j=�&f=�=̈́����<��ŬD=��ʼL�5=	�b�@��"n=���j(<�ܻ��<��L�!7C=�Q�<��q<�j�q�A=z�<D����h<Qּ"z��<�==��P��?w=��� w�u"=�M~=�����d�<S&</ ��n�<)!N<�]��v�=u*��P�q<�/���'=��&��F�c��s����;w�h�Hb���t�-h�&:=�bC�V���+I=	�@��=׼��Q<�c���<7!%=D[L=74O�N=��K����c��uT=r�
��![����;F�=h�m�
X�<	nF=J��< ���	��<ƴD�}^+���=k��r����.�=�3�坛<i���Ҵ��^�=B\=)�<������L=Z�i����Oȼ7"�<Bol�Q��t�;�T=,r��ml��PK=��I�M���l_����;��@<��< �;�3Q�5��<`㻉�D�S�׼�=.B���ހ<]%+=�)�=!L��
�@=��<���W�=|�)<�G=Y"�<C�8='��%�l=��N=<=N=r%M=�[�<�ts��L����7;n�E�<��;�M&��W<��=|"
��&�
�����(=��"��0=�V���O<��<Ɍ==�=g���=��
=���<�;��K�'C�xP�<6.�M�<oS�<�Ԓ��nY= ˼}�<v���@��=K#�;܀�������ʼ����N?���T��m=���<�%�ù=�^�<��;=sL3=%�^=�X�Ӫ�<���Gwռ��<��*=s`�<��N�,q���M=�,���4�=�@�NZG=2[��BΨ;[�;=�Z�� 
��"�@��C_��(S�>f�1#.�G��<���;���<m`��%�;}��<]
P<�z�o�j���<�=�<�!=企�
��T1=����]
I��D=�*=M2�<��w=�� ����<=��;��;%萼�t��i%����<52ؼ.^=��-��70<��+=�S�<ݗ��.������;���L=5�
=�D��<��O=��=e� ���@�ؼr�<|�Z�V���ʊ�ND�<V �;����E���Į�*�]<k"=��?=���<���D���=e�<!�&��̸�/[��w�[=n!=[A2���c<[���H�p�r&�<�w<��;���<)�]=�n<���<:�$�PBR���<19v�K>=��W�a�O<�r���kcn��X�>b4=C����U<AM��;V����<�͊��V��=���`�$�XݼA�v<_�<x�h=��<|+T=���<�}�<�\������g��/)�F?=�����Q��"����i�Q�P<�&�<0r���ͻ5>ɼ>0���Ѽ"�@=��V=t����<��$=�:�94;�<������-��][=�"�Ǝ^=�`<ݰq�tM=��DA=���<� 9=#�<�fY"��<"��E�Yu4�z�;�6v�m ;�YU�X뿼��:��K��������1@�݈�;W�<��%=u꼻V<ؗ(�^獼C�=#��0�J�m��Y��(*��:��ܵ�<���/�cvE=84�m�<�� =2b@��c=����E=w�ڼ�pn����<+�<v�<��<�!9�#;�H=u�y�^+V<�R�<zb��p��.�<�%���z���8���#�;��ȼw�8�[=�B<���-Q�<0�H�+ܵ��)^����;"�`;�A����C{��K7I=_:<"]i�B/�<-`X<p��1��<;Az��\n<j��<l<<Ua<{�M<�:4=S;�<�� 8�&,�ԅ��;&��2;`�^<xa=����	T<K-����^=ѷ]=�?��������zd=������<����2=���f+=�+���t�<v��<-���M=\��<��A�6t���/U<B'����ϼQ�<(�Լ�&=��U<��7���<:��<ڙ��K�ڼ�I��=���U�r����"�T�o���c=��<tR��5���h-=���L=4�<1Z�a�R<Z)=��#�l�=C�6����<�D�6=o� ���uL=7ͫ< 3f�e~s=5�;���X�2=$=PX�<4:�;��<������1�<�.=.І<6ɒ������<=�E�μVv��M�/���=��O=+���	<변=VS)�k٪�q�=�?"��|L=cG=�~=��1�ͬ!<��="��\=��0=���<.�A���o�_�d���=DW=m	 ��<�">�8��;�H]=�<}+��@H�-<=����*��E�a=��<����q�%�#G�<���7I�4��<5BI��<�V�/�%��@�+�;�(����C���Y>�)�=H�k=^X =@
9=\�8=�;��KX�6c=��'=A=�TʻF'9�EѼ�]=���<v\;7µ�J��k=z�=��<�z�<"i�0E�<LH��99�<������B�|v:��R㻴L�<(����1���U=B�+��#;6
=�yvr����;]���tQ=����oO�%�=<
��V����;4���od�O`|=I���u�;M����)=B=�^�:�0C�k�:=�6S��'N�k�I��<A��32�tLK=x�:�)��oA=�4��HD��pX���� �X=��=H�߹_��<H:<�45=������cR=�n=
�k��T�<�hX�PC=�a9��m=�V^="�<�)�Y/^��R�;N��F=eQ����q=�u��I�c<��V<}�d�t���7L<d}�a�D��FO��5��=���=�ɪt<�\=]Q����</��<,e\=R��<�,m<�s"��ZB<�w<�\q�y��<�V��\F��LI�;���i��<F=<����"���E5=�84�.����h=r�[=��<:�M=T3�d��Gk�(�W���������<��.�+/<�����u����+< G�}����<�]V����^+@=�H�;���<y�O���c=z�N;I=�h���Q�L�:�~ ��8Ƽ5-?��y��['�}�`��-���k�;z�=+���e���P�;�6=�:绣Bs�FZ�<���;�g=�a�<ً��Ƞ<],	=��=�'={s����O�b����6=�-�)��<���<���iڼ��N��(i������)<�� =�{�;�M���9;� �+�r̊��G9=#I�;�p\=KX;Yz>�|��uF8��b¼c������&p�<��[=�,��!�<���=���a��;b�)�z�1���t<�� ���<=�)=��%<U�:��μ�E_=7&���#=F=���;��=y].=ݨ(=  5=��_�"0��9¼&���R������$�G�t�=r�:=��<��H<������脼�n�;��2=�p�<��/�:�T='�⼑ٶ:�@=!F3<�\=�T���g=�4y=Y���м�]��������<bvμ�F8#�;�_T��'=���:�&P����Ω细��<q��<Iڢ��F==qsZ=��N�����F�0b!<B'7��=J��<�W?�~�=� ����/���<�4�<� =�ld=Xh�E�	=nq�<5��d9Ź	_T�!�#=Cg�<�e^�.�8�\�<JM�<�x�:Ϻ<��<H<%j�+U���<�{���;��#=�P<zx4���*=�e��j���|���+
�M���%M=찒<@Ci=_�)���=<�,���8W��Ea�R^�;�;#���D�ȹ*=j=�3�=;=1�R������o=К��.�B_�<��j<	�ͼ8�%;x�����\��,���w=prټo͹;fb�<#o=���<�����`�����h�������=`4<��|��6=M�~�y=E4}�A�T=˹=c�j=~R�� �]=�T=��=&Ke=��8=��`<�,��:=�<M��v<V@�<úd�=Q=W�=^�a=�nK��I(=j@���<6�#<?���d�s�<��<H�@=K[������#�	�����0��!c��Ǣ �#�<u�;uƏ��#���?G����=�ļ���� �X��I=����;�<emQ=m.m=([R=b����� �0L���v��P5��)�h�<]X�;�G�<�v������C=��L���=�c=<N�<��2���;���<��1��a�<���<�>��P=>�<~�=徏;�U��Q�<ZXɼ��T���ټyZ׼h4�5�#<��<1����ѻ���<G�ļ�R�<MzM<�đ��sK�����Ӿ =~O����<+�*=��=0�*=�w�<��<|E��]���<�E�㼝U��@jV=x�Y���%��B
�P�Y=��׺��>��8�<�[�5�)�^��߳_<w�I���m�^���<�żH.����ƻ�^�<��w<�Q&=��;��;�(!���=�Ë��<Y�J�W�=��Y=�oj=�ݾ<3ȋ<��B�r��<��ټy�üjGy�s���<�<��V=@a]���<M�<}i�;!�^�D�E�U�~<Ь�<Y�\=��=��#��2�<0�;=(��dm<�]`<����u�B��<)%=e��[0H��輇O���<�����';��Ѽ$�O���r�(�=�+y��ي�<ڧ�:1=[f4<KW�<c�`=�=1.=�|�<� ���<ێP=���e���a��P<�<JY�9UU��a#��a��0ļ��k=�U�<��,=6��~g�Ϲ�;#��y=O���=t�7=ߋ =C]���Ę</+3�6���b���)<B=1<�	�}����^=@��:��B
�s�rf��0;�39=�đ���m=[g�<�%;I
��T�~���1D�>e��=F�C=�=t��;�'(��E�<<�M=m�<=R������}=�'��a�z�"T@=&ž���l=���<t�O=8_�;�B����9Û<���A��	�<׵+�%8U;!<�l��'
)<�O
=�.�<,Y�<��7��P=�R=�a�;�t�����x�=��Z=�&=��<|��ATJ��F��!=�#����>�Ƽ$޼�'.=�`�:��<?���3�]<�xA�b�x=�gW:C����$<=�&2=� =���-�=s��w�"��+�������<�[�<~��<��?=�v0�t�[����=WUĻ�>�����%=��4�`�?�/�F<U��F)<`� �'�;,s��0鼊-�<�
W���<�"=��"=F=Z!�v�<7d<��n�p�ݼ�?q=#=3��<>0^=��l���\<���F>����<�͕�c���&�<ڙ=��k<>ٿ���"=��@=�-�L��xͼL0�;_�ܼ�8��[������N=�"'��r�<���w=�kC����<oi�=�>���$C=�S�<��=Y��<$^��%���K�sG�t�0=�4ݻ�(������d<�|������,����)[�=<=%���~��<4'=�=M'�<=��E��K&=Zt-���T���<�f�;��=�}"=��B��[H;߿3=�{=܏Q=�+�<@�1��� �+��]p�!*G=$��<�DT�x�&=Y�
=Y&Z=��<�1�`�(=�����L;!�^�->�<o�l=2������:��8=�G��Y*�;iļ�t���ϗ;�T=֫M����`)���S�˜<H̀=�?�< �:M�<�����/y9�8 �<J�=�q���<h<w=�)��~����,�i3�;��R<j;��T3��D7�$�&�=��5�z���nP<�<gZ����<Vw��4P�0#�<�6=Ӷ�:�h�<P~��ճA<
k<g�-��}z�}L�1E�<���<��{;���h��^���[�Q�L�<�垼x�};��_=�1.� -N��$>�!�¼�c\�ܢ]�U�<<dм�[�<k/1���O=5�N=�E�;{�F=�3<�m��=l=��g<9����i=t6�<};����=� 0�8�i��P�@�=�=�<}�ּYü�I�<j��'R��DK(=�)P=���л�<���8=��+<�HǼN�;�	׼��;"n���,�.^=��P=��=z@��3I�_�;����&c+�Ȯ<�Q=��b<�v=�7�? �<�
�M�^=�j�[=W��(�o<yjV��N�P�i=1qC����<[＼%<�Z�=�Y)=?���w����>�)�n��f����.�μ ��] =����E��<U��Ѡ'�m�k<�����;:�ּH�;ʾ���4=��
=N��<��<A��<Ԗm�Z��<�1=� ��X���=R)��f=�-�<%G.�r6=Z6�y�]��=�;��:~�8l!=!��d�ּ�:l<L�	��u,=ǜ\�ڮ1<��*�5?{���9V�=��W=�:4���5cx=@�P=Z�<Ŀݼ��<Y���z�;��=aV�<Ӆ�7��h;:v]���}�G�[��zB��@=^/U��/=�uO�>?/<�L=%EL=+�׻K�{<������<�=�_O=mO=��#=�j��
����^<_*=� ��^=����3=;Ѽ�A��̼6�e�b�4G���� =?��d�-���\�M��F���N�2=FA#=��ڼ_�޼h�v���<K�*�J~'���Q�������w�x.�kTg<�X�=���<3x.=�S�Ց*���=g'k�rRͻd�Z�z���.��<��8=s�,=[���;�=�nx<W���*0��BR<K�b=_E=]΂�Ø*=�O��N�<��N����;S��<���<)�]=D�^=}B�<�L=]}�<���nܺ�r�;�G����^�<nr1�,H�X,=����_�d�5=!/5<cIm<�3G��I�i=+�7��r�@��<}qH�R�.=7S��	���<'�6�7^�<��U<7W=��==�P=+=q�;͘�f�3=��ϼ�P���o=�C�<��]�5�;{_<�ސ<�T=ʜ[<r�C<����vY�(����<�a =<.x��hȼ�N^<Ԃy='	e<ד>���o<jź< �I���N�|Ҽ�~J=X5�j�i��<=f�T=�<@=���|��GI���C=_�x;�nF� o���q=�=�ӻ��໶�I<gR'=ůf:�a%��Q�w4��,=�� �(=;�������*��,��n{=���<��W=��;�z���AE=�s���A�8�Z=SWU��3I=ۜ�tE���l���k�;��=2�~�S^=�ԡ��¥���:�Ai��s�ܹ�P��	Wp=th��uH=�M�;EgZ�W	N=ls�����p��<5�׼�r�"6���1$ݺ��T=��黣�8=�HY��p�<�6�G���3i�A����(=ԴO�:4��1�<�&�>+�;���<e�=@�=��c=9����a=�=���s<�=��T<�WF=�_=Կ�<��J���b�{�Q\�<�,/<��=��4=hm�6uR;9��Y�,=s��<)k=CkM���1=ʷF=�kؼv��{�i=�I=ݓ��к< R=--=~�"���C�{��-�D<�=iS�YJj��_�Dv/���ּ�W��'=gW$��7м���
�;�.=�@���9���"=ǋ�<F��<��4=0����R=a��;��|��<��P������!�����ȼ8s	=��~=�P弇�:�P�	�'.c��$��QG=|�'=U�1����;�
�9�¼�)0=�>�<�7r��4�=O��i��]�o=��뼹�!=m�=���@b'���D�j�b��4� �<�ܼ��#���p����,�$��]֒<��<�/�g�D�/=�5 ��$���������
&=Bu8=}Xl<Q�d��V��Տ<�.�=e��<ST�M9x�nނ��1��k%=S4�Z`J=�*7�|� �ڙU<0��ᘭ��C,<mkO<��N��,=Е<�s�<��V�Fa?����'g�N�;��������A �t�=]ze��e�<Q\ ��$���f=��V=�e�;� �7�5��7=�P��6��� =��<ҹ%=鏌<�8F=5�=�9<v����鼐X=*�<�M=v4g�7&D=�4�ؑy�#C�<��l�1� =fI�.�S���r�'?=qb=�=�'ʻǶ&=y\���%� �8��Џ;�.ǼK�&=aH<D�=��=���<Œ�<�M=h!�8̕����<�/S���<W:	����Cc<�%�z5�<�v¼������<�_6=
-�;2��l~�}<��9x;�6\����7}c<�-&=���ָ�<�o���_�f\ʼW��<��K;8=G3;=�\�'#<X$A=�=���<2�.�Q@����)=��8��L�<O�ϼB	��I͂<P�9< &����;�5����X���<�6�<\>�;)7�*�� ����|�<[�����]�U=XN5���=>�:qF�"�(�;����%�	^h���?=2:��Mr�[=�<�M���<�\���F�[��{W������Q����1/<����(�]=�m=�"<{T��1a�;:�<�.�<"ӳ;�w&�o�i�h�:C]Ҽ�Q;s���<1�u�<��>��D<~c8;�+�M�@�q=OdO=��$<��<�B�;���*���LF=bM4<�R���y@�.=��)�o�J�0!�<�&O�3:9=�{�w9=b�<�>�;�;�!`=  ������ �.in=�u~=�+O=��R=��F�+h�:���1��H؂;~�<��z<	.=<@�<p���p����͝�<}Ǥ<�[�2a2=,tȻu�=���;=cX=��@=\�^<���W�!=�)���,=��6KH==�/�ڼc��<�X�d=x$2��D��R=E`ۼ(�Q��ۆ<�� =��;�^���);=��W<A\���6��D=���:��V=�#����Z���<U�5�-�D�e�q��g��>���8��_1"����<,���ڭ�r�.��a�<����R��:�nɼ�Y�<	-4��v���}��@��3���=��f<������iH�NV��Kp<�I�	=�n���;K�3�y}˼�M�<$��������Լ���� J=�A��=�+=À�=������<+�5��}˻��=wl�<��~�I=Ri���w��Z�Ҽt-�<�L��H��i*=��=1�;�{�<����ʅ��1�h&<Q�S=�S��yP=��d�y<e�<�	,=z�=R�_<J����l���<�6�;d��<
ȼ���Kq<�%Q���<��ȼX.�<�z <,D;�!U<U�=��p=��<�%\���@=�D�<�.����<+/���;����8�4�<�ct=}?e�oH=�9��{�U=`Bp�v�I9UD뼶~���{#=����	1=z���|Z;A�3:y>�<O�5=q>�;���\P=Z���mSD��'S=�ܼʜ�<Q�<&jU��/��`<��]<���<����o���!;�s�$^
<+��<����}j�E�޻� �@RK=�þ�Ku=��<T�a;�̴�n�<� a�t�;�{N��&�<+PԹm�<%Bj<�����T�GA=��w�9I3�	/2<�dۼs��<j5
��^���g<_�B���b=����G ���� ����1�~�-�<�J=��μ��d������b���#=������y�b=7��;:>�;�u�=�!�!�<I
=7.��W���Ѓ�������n�V�斐�N!�]9�[jU=X ��/��o�<KC�<�I��Q!g�ɝ����}-<&�9�c�=�n="�������R[�;Պ��$�<��<�K=y�g=��<������\�J=9N#���;agz��` =�*�f�=�D�;u軟�#=���d��;Lrt;h6=9繺9W��=�#/��U7��uS=nJ���X<}͛�����-=������<6XL��(�<������S=D�k=�m��M�u=���<'#+������;U\=߼��/= VP=Nּb�9��� �K�E�tII�k�@��z=v������]�g�=
d�<�wu<�c���0�<3뷼����'=�\�LRļZA=B�<��B�Ea7��X<=^p����
3=?�|�~ｼQ�%=��<=SJ{:��$=yG����<�tn=	w�<��H<��=�	�<\a=L=G��~<8i��_���/qw=g���ni��𻼌s���c*=�Kͻ��T=hT3=��l����=Xg�s[i=�7�< ح<�x=�=-=�!���	q=�&2��-=z֕;WE���r��x�=��L<�Ŝ������C��D���ǂ<<Ɠ�'7=D�<��8�2<�,�y�
=��s������]�=y�������;�\<�g<ɵ/=�=���<�^�=����5���^Q=}�F7�*�7�*H���8��!��"�a���<̋K��U=m�3=���;�+
=�����L=ڇU=�<GV�<��^=�[	=�k=j0&��&�<�9@�_�j=û<�-�<F��W ��b(�UB��h_="��;_[<j=�����<G�&=��=��-�=�׼.�:IE�&|��<\�p�=��y=H��<�T��mGb=L��<%*���lؼjK�Y��V�!;*=�U=���<�7%�pA<���CӼ�9�<_�������<jeȼ	f�<�o�<�m ��C=����EټW��<�%=�:�<Q�=�+p=�����;�N�,��<�[=j$=���;�w'�W#m=�1�<��*��-��+8=��K�#��5��<�c#=Y¼�^=�Z]��z*��)+�R������'&u�z67=ౄ=�r���t/���3�/��z���=�P^���r-�<������Q2�b�;U� =	]���<��3�:���<��<��4=�B�C�Ӽ���
�g��]=4�Ѽu=�$�:Z��<e�+=���|�&�>`�<\�V=���<�*;��F�&4���y�;���;��<^zټ�V=��˼�H�:!�T�d2���2�<�� ��WR��f����W=?�Ѽ�6���=�g»�"���˄=G���E���=CT�a�H=]=ѩ<��F�3���׈���a��xr��c�:�4��fk=�B?=��0=�f:=�
����3���U�x��;�P����Hp��x�;N��<�b<�^��hA=	h;�Q�;����n2e�&!����K��9�Ӣ�Od";�=�=�&�<��׻9��N��<�������=�k=�_�<���xE;��M��砼)����0=\���=�ֻ��P=����ټ�p���9=+7==�9�<uF�y:���Ho=ɚY���=����/Fg�:�"��z���EH=�7q=���<K^м�B���p;Y�'=�x���vL���j<���<�>��)�=W�6u�;�U�<E6Z=%�B�)�<y�#�;d��&y&=� N���k�\D<z��_w5��9?�C0�G�<�`=	S�=����'lO<_B��b��P9���Ἴ߽����=ұe=�l=��#=C�=�PZ=9�9����h�;�Jn.=�~g��%<2Lü��h��� �<&iڼ�e�<��!v9��	�|$E:�sa��ǟ�{2=)��<��W;�2�ÑǼ�E;=	�3=�s
��)_=V��|^=�7��Z�<sK�n>�KE=q׼� !=qT��(�I=�*�<̛v=n��	�!<����λ�o_=�N+=�o/�0J����<������<J*�<�M����2�[�
�4<i�-��|;��� =B$��-=�=(���!C�7��<�g@��X</�B�%|n���F<˙���H]=I)=��<AG"��y�<�@�'�6=i��<�l�K2�X�:�Î�Gy!�n�����!<��"=7�"�<�|=G��[��	^���s<D�1�bb=Ni+=�b�9P���fN�*_L=��-=�bM=G9�J^����2�� �:��2�0Z=W����R��&�<��==��<���'t<�G�S'�<�n��4��<ɜp��65=���ɸ���)b=���:�)�;h�;��;γ<�<�g�<����M�m��uŻTk�<�4=��9�FJ=Wa�<�I<���=�D���=:R;�8�Y<���e܇���-=
N2�+�A�l�߼��9=0 y�ƙR�u�Z�#����ۼ����Tռ�_�����l���&J=w+6=}�|���?=�<Y�]T�=|�<��n��������<�i���Et��*< �;/�a���y�<7��y=�E���<�ƻ�2=��	=��
���L=�u�=�XN�L:=��E�q�=�Z�p:!�ț��O��;���<=L"	=���<Y�� ѝ�яr��ⱼ?cr=����Xa<�6���
��q�pM�=�a�|�Y=u �;C�C���d=�e�<bj�����`�pB��мJ�<���p2�����<�P=�.=����d<�<�*���O'<��	=r�=��˨<�� � ��fJ;{z�RВ=%߼���=��<|%5�2o�<�B�<�1��O�;\���<���˻;��:�&�O����(Wq��w)=`)��t�k�����f�ےX�K<�ļ���	�X =
�r����>;�c����ɒӻ	2��;=ʿ��:�Ƽ��;������R��<�s`�"�`=:�=P�<!�<�;a >�<<�鍺c���ػ��"=:*O���S�
����ܰ��G`��p=Jl=�s`�:T�L=�d;w�.=1�;��n=�L���{=C��<�9������μ驾9��;�M=kmμ��*��f�G�9�B7�-M=�D=�1�kH�<~҄<wR�D����Ys�
<<ֱ���;f�b�;�=����
�<}f+��C\:j+@�0q	=a'컅�.�p��;4=w��<˻4=K.�ELK=$S{��!��;u��C"=C�H=J3�:���<Q4S=	~����m=n'&�	��=�	�T������<w�=,':�TPN�+CB�8t=�K<78�<�#<�\<���<v��<<5�̖�	����<)��<~
�;�"��L8�L z=�<��hQ�|���}���ڮ1�!��:����Rz�;s=�����0��8ּ?�L�[�=xX-=�+f=�^����I<��'=��=椲<{�<��=�Y-<�1=���-� =9�n::<n�=K:���:���ԼVH�f��<@��� ��C=�H�c��;���*&�<��<j��t,��]����b=Z�d��,N��݀=�[=\��<�8��Wd��}F<�h�;�q�����vW=�}9�~�x�i��2�s}.=.P߼qDT<��:=�� �R΀=�Y�o�6�g7������Z=��9-�Z����<�vQ�ɤ8��HT����<���<� �;��=�L1=F�t����2Ov:�D��4,<�
��aT��J������Y =�:=p���q,ϼR�y���H��K<ީ�>P�<��=�}�<j"ۼt�i=�Qh��� =�c��@�<M>;=-��qNA=O�3�rt���=˰=�O�e����	�9l�=�d;Z�1=�n�=��ú=�-����<}��I�;'&�<��K=�c��p�<<�<�>$��0�x'=$dl��ݼ�N�BL�<I�*=|��<���<�1���=rw�<z��<Nٌ<�` T;�}R=���&�<?C&����<����Y�;��=�����^�-=�<���uT��;<6:�>����=o���V�V�?�ټ������N';=L+;��!={3�O��OȤ<�󗼇
�`�U<��=㸥���ټU<�O<�e%=��`��~n:5�<<�F<1ۤ��O</=�i�;����＆��<��[��� E=��ļ���<"p�<v|�<�0��1�C�<�V*=30׸_�ʻ ��>���\�͗<�lX;�I���4=zX|��j�;(:��q��pZ2=�f�:B�κ3�=���<��N<0D�/[�<��)�ZGѼ�i�<� 8�����"���=�K˻ds=�~>9�M ==ݼ�b��m���<2X=V�>��bi;\�]=^�C��w<���޻�;Q�<ͫ�:(<�J=��B<?<�<�ؼmx{������f=��p=$�Q=!�P�J���-R���;���<�������<E����,m=XQ��:�X\=���<뻆<-+$= /�E0缽�:�	\�<V���$;��<��=֡�=��üT�C��=<9Q=�x=x������b&=��^<�c=����������'=q�+�n��")�;�<�����;�*�WB�ƿP���=�dI<�䋽4Z���֬<7`���p<=oi�<w\��YB=�3�<��N=��<.��<��f=��˼1m������L����<3�6��2�=�L@;��Ѽ��;:�;�������<����<:w7=-L=�s<2�'=*��.�X�t=�o��e��<����6h��o��蚁=t�����<4�+�^O�<z��<n.��.F=,�(<ps��Qx��*$�x��;�
<��i����x/]�-ȼ��<�]b��y<��g��t�<����� �T
<S�N�)}���;6=�h�<ȍ8���=�[�`�;��<(�<!����S^��zt�����+=��W=8^��v=2Y=���<߼ ���<w%s<�_H��'�<Į8����< +�,=�U^�1q���8;&�λ�j�y����6=�z:�r�1;�T�-k�������r��#=�m<<u�#�=��`<%�=L��k�=�Ƽ�d_=���;^��<�v�<���<6��e�m�
9*���W<���<�Q=��C�O�<i� =��7%�<O��:����A=�ܠ�	X컽��PnL=(jg=�,U=�mZ���7<��]=����<-�Z=m2��_@�ž;�-=v�μu�8���Q=uYA����:��0�}N�6p=��(:=��#��o�<
�1=�d;��ng������I<9G?�����K ���f�=d��-=��2�1<?nu=!�D_��2)��D��-ڐ��ҼB�L��<�X=�����%o<gq���zI=HI\���B�]�9<�a9;W��<���j	=���k�D=������:�%�;!��0���@T��1=��=hE;�<�[@=�Nͼ�� <.��2��Ih.=�<&YH<l+�xR=��-<�h$=�Yf�{�:�H�<��$�.=A���yg=��<F6==n��<9��S�1=��<;��n�VG����=�u"=�mg��μ�)K=�=p)=X��<��/����<;>�l5Y=�*T<�伥QS=�S��e'���=k�%�b��<���;L,��>=_�^ʼ�EzT�ZA=�S'=�B��	=+����:�o�_��|X;ڜ=��9�<�n.=��-�aco�������;�R�\kV������"�� =ӫs����<��3SǻO%<�En��!<=��C<����K<���X�W��P"=?uT��ɭ;� $<m����[��*��;{��<�m���w�!�;�8<r~<��';VC��D�<��8=������ <Z����ݻqt#=��V�z뷼��i=z�o�*��<S�c<�ԼY�ͼ��N��	�?x ��᯻}�=y�����<S����ð���!<{�-=�ź�c=�c������b�<+S=���U�"��<�����?��<�8�:1��<O�f=�e��g�<ͅ������@������F:<9��;^d=��=�a��Nb�͒O�"�<f�D=�&=��&��+�K{�qռ������2���s=z=�:�<�Y�<��<�X=N���(=��;�Tr=�c:�^;���<$��<cPҼ5r�<�r�����<�[�;bg <���;�*8<�}�<'$%��:K�^7=�a<�?�<�qF= k�<�:R���<
�^�f���c�-<< �<�*=�Z���R�<�p(=}f&�@�<Þ�<�,f<Z��<4��;�3���+�4���]�t=��p=���MhJ�d��%N=^�i=���������!U�<�8W<�U��ԃ��Q���C<le��L
W�C _=����<�
���&=!��>�<�;�G<�Y6=$ռG<�-��<Ų
�o��<kwD=��<y6ϼo�/�����Ӕ��<i=tq7��[�+=�;�p?�}��{7���=�T��ɷA�_<��w<E��;њ
��x2;0�=-�Q=� ���<��2=�<?=TL =��0=[;=�q<�kA=�C�􀙻pe��x7=��'<Nq���?��<�<�ו<�F;�����U=,S�<��c= V"��� <p�"=bG�<�č<�Q�<Ux�;�	�9��<T��<e�(�j�����s��΂=�f8=4�G=E�P=��A=��L��%=m��bEF=��H�Pns<x�X���-�`CA�������a�����<�mT;���q�<��ټ��C��^=��̼d7p��&�	v{=Z
�i��<����b+;5蒹�O��[ܼ� 3= I��P�<5�񼎶8=M�\���.=,Q�l8<B�K<�j�B�= �<>�ü�?��N�<����v4���=��p=t�1=00�<��:�b�5�U�L�V������=�3E=m�h�V,��}U=��W=��6=�#>=�$?�Z)Ѽ�=��*yA�� ���h���&�<�N=P�+=ЉA;=��;��<�t����U= �/���7��(1�<L4<�*�C�>=��3=�K6�?=�<�|<��"�=	
=���ةڻ৻���I>
���Q�.=:;L�V�:�Vݬ���<")���� �^���o[=.:)=W�r��߽;�l�<xl>=fe���<`���[���r=��j���<1	�<��<�|�Y=U�Ӽ���H]<X�<�����<Z˦<��H�/8[<AlJ�sR�R�s<��g<��I����<㪿:H_�;����2���^=�mӼ��=��r��=Ý0�)9��������0#�p�<�=R=��K�K=�i1=D꫼:��<�S8��Y=(�m�،�<���<8R�<N��<	3����<�A>=nB��6B�b�\�8�:=����P����<��<]�Ӽi�U��ʏ�L6=��qE<�l@<H���D����<�5\�Ӻ��1bd=O�<�1�<B�<�7<�=���<��'��I��U
=�J��<�J�<���s� 7s=�$	=m}J=aE�kK	�/��I�"<��i�s:����<0]��X
=m�*��;�^�;ص�<��c�#��.�<zJ���+���漿�h��ؼ+�)<u���f�=m�4=޲_=����:=2C�E\i<:�Z=b���.�:&��<���Ů������;`Ѻ��%:��4<l-��6��e�$�;�k=P���٬���9H=r�_��EM=bS���˼�K<� ����=�zn<�_Y=F#�=��<��<�2�<`�_<�[������U<i膻��8
=��M����9�KӺ�;�;��+<S�����q=�Y/=��~<�$$<��b=�c=W�)��L<�6.�>�<��=F��<^����y<µ�ֈ��ƼT�&=��]���ּ��=��-=��<����.�"6=��L=���RZ����< (<�=���<О^=��Y�\�=���"V��(M</�=j�K=��;�o�<�0��~s=!�<h3*�M-�Yr&�ܶ1=/�k��<��<4wR���N=�]�<��<P�<�`I=|?�<�ۛ�����4��j�����<��b��G�<�l*=�8�:]`�A�c=iW?�����O;�D8=�v�<h�1��0����������<5DR� }3=Y�<�l��u+<u}K=H�H��7r=��w;�Q<��W�fr� P�<����[�<w�ļxǂ�<�=��J���A�z�F����;&���1J��~<t��g��V���PY��C��&~H��]<��=_��<���ƛ�jb�Jsa<��=�4=�f1��=�ܯ���1���Q��}�< =0	 ���=�����+*�<�sU=γ.=��U=kR=:���a�n�E=%>�<�@�;����_7�|Q�<r�T�$�L�sg0=��>�a�򼗟 ��Ș������H�K��=��<s@Q�t/��!���4�<��
=\=���<�j�<��p<�=u��J��+i{<cm=4c��0��/`�&��Z���<�p�<�b~�l|&=H�	���Z=r�3�w�IA=;��ּ��e;��g����W�f<0!�=�=��e�z=�[�;v�켝
4=m�μX;�3���W����`/=�=�AG�a�M=�����)4=`h�<�Cs��)�<�y�oqV=��6<�%�c�l��(M=/�O����!�;�u<��I��_-=@�i=֝G=�&=�pN=-���m�<3���y�<�4@=��<�@=�R�8Р�<Kw=�bG=xnӼWW=���<��R=����7G�8��<�X=¼!�'<�h;=f�<��<����ۻv�>=��I��i���켖��,Ք��r�<C�P�� �N����jz��|+����<�Z=����
5��%=���V�ʼ�e'�#rW���J=��;p�J<��I��=#$� �'�^���,Z<�m�p�<c�=���y�*��<igt<R�=�\e=Qu�<����K��,�I���������~(<�f�JM��s�1<����Dy~��úH�3=D�<��B�<}<�I��`�'��*�����"_o<������$4�4��<�ɐ�35#=�s�<03
�����R�<֚;���"iN=�̙�����L��q=="'=^��;�p���H�Ea�:m��ߚټ��m�!=�L�<�B���t�ɵ�:0wM<g�<�"=�?c�<�;=���g�;��<��<ǝ=�e�Ј�<Vi�<���URm��@�;
ֻG�%�N�p<@k&�K��;��<�C�<=5X�'#�$W"=��%�d�$�HU׼����}���=T��b>I=ͦL���r����<@�����{�</�;j�*�_=�Vͻ\��<�x<Z�Q�/�)=���(߬;7=4'����ݼ<w�x�<��-�Y�]=�i�;�/#=�n=�4>���w65=�w��0d�?�)��8�<t��<�f==1<�xc<s��<iz&�l#=�N=ܺ(�q��q����a/=��V<���<j_}=w��
)̼�柼����e��OL�<�Z��z\�'H�6==,{{�;o=����ٯ�8�1=6�޼�7�
I=��=��C=�� =��$=��l=-�7G�<��r=���b)�$��<��y=gp�;��1=[B=�DS=�#<��[=C��r�Y�\��<ŝ�<�<w�,�@���0�;6�V�㿼!8q=���<5�w���G��r����n�`�l���T�Y�����<�爼�4�<�މ�yL���5�P=�X9���; ��<u͹;��@=x/=���9�3�<M��<�/��km���=�B1={z9�*����T�����v�=�tP<%�4�4=I�<�D9=;�g�\\=��W=[�-�RC��M����<ژ�<>�i���<Q}-�2K�<aXݺ�O�w>�<��<ۏ�<d��<N�3�bK������GE���<#Rٺ�����<���<��T_w<N �<y��;�W���V=�H!��vʼ5��< '��p���ڼ�]Q=ʂڻ�I��갼o�i=WC�R�a=�w<�Yg=U}ۼ^a=�{�<�01�9N1<�z=l&=
%���!�[�P���"=��\aj����<My�<�Q�ckG=�LP=0lG�$5_��;&=��;��k�^����=w�=�aM���<��:=�o�<-��K �~�a;�'�<��<�*�3Dw�&�3=�t��H}V=�WK�k�O=�I$=��;�"��cS=�����<V��<z#T��L=!���{�<RX�<|�<��K<�6�<:f2=�ك<R�<�2�<�l�<Y�{��F��r'=�)=��T��U�;C|=>�X�ү<h�}+�<��:=;S:�=>V8z�=᭽�R�����=�����<~�;�a=��M��n弎v��/=��b=9�(���uX��$js<٤�<�Y;�����m���q=�$=�ƺ��j�4�L������R�tm4<��<:��<b#+=ŵ꼛L=�:��<'+=	r=`��8y��/~��S`X�ކ��	:�p<=XU=U�\��Q^<�%�g�,����<��*I�{*���;�t*=i�F<޶&�$���;��<�5��ټ�p������<�P�Gr��d�����<��)=A՚�`W=�̇�%�V=}}%���Ӽ��<Ă�;�Ђ:Q��<!P����Ƕ��np�)I==�����;�h��ƃ&��v=�5�<��=^jq=����$=$��<��Q;	��X
=�A�:~3�<��R<W�<S�X��6��QL=j���`B=L�R=<���Pr<��������b��gP��{���׻6Wz;`�̼1����<|= b���� =��Ǘ�<��#�G�<���:���^�=��f=
漙��������;�UG�W�ehd<v����I<��=������=6fv=p�漦��<�9L<O�n��S	=�o�SA.�[������������;�$�;�=�=W7<6J<S�ü����Mu��ȼ�ټ��n=~ō;#���x���0L=��a=,Ѽ�i�J���d�5�s ʻvJ��*�;����Ų=%i<=��R=�ͼU��<��B�w�X=�?Ƽ�ɼ9
G����C�<�d =�<�1��|a=G
%��X�,�$=\[=+;]��Q^�ZW�<��K�D�q�<������|={<	Q=���.��_����=L���[Bq<]<#�����;�W=�-��RN�0�ʼռ�u,���;)=u=]��= �)$T��:��ѻ|U�<��9F)<KM|�\U=��^���<�T��l�>=��<-�[���';+.��Ӏ�.�;�&)=z,=9L��O=�����Z��bR��[;�Rs�Hz=�3<L�5�d�<$p��P")�"I�;�n<^y����`<)C��ȭ��j=�B=��켏'�#:s=�x��Z=7~�<Ƨ�<W����8��]G=i�q�9o��r�<,-=�I5=^�=�=M=RNk�8-�+���=U%=�{=��<��ܼ4`<�`���
<��=A�l��Z���F=-hk�BaH�ltP=���<~G[�	�\<n�F=1���i��<�I�<������_<7]=ML�;{~L���:9+=�a�<}W�<�7$�a���LT=8W=U�{<��<�G�6��<�oH=i��m����;�;���5<u=��<b����l�<���;g53���P=�Ij=72��o���?e�^3)����b#�<�Q"=G���7=�أ�\b�=�����0=h,m<*�<-#�;X��<ԍ���n�;D���x=W�S=Ig6�~�ɼN�N=�&�����6C�ו�Y=���:x�U=@�'c��y�� =��X���<�w���ު;i];���<"aK=@=���}�;�5=dVY=1�<��8=Dc��$��&�G9L�-���8��⺦���#�'=��=�3`��M���_ռfL�^�u;��K=��<urv�҂����>�[�m��2(������.<�}m�?�<��>�O'=���J�=�,t=H������R��̫����"�t�<��<$�e��@;=�;6K߼�����~	={�"�Y�:=j[�:h/=.%�(��<zC��.B=^����;��><�R��dvf=�rF=;Lؼ2�$=��<��Qͼ"�_;�D�c���^�N
U��K;���vZ���<�9=ϼ>9>�wG<�SG��W���=��"��*����=In&=�?=��<��L�m�V�n<X��t�<��C���<�sY�<K?�9/B=7E���!���
���?=�,Z�ۤ��:�%�c��(��|��0L���<���$<�S�^�h;!x�<kB��ܵ�<Չ�<'J�<UJ׼q�u����<�`����=�BU�*<ar�<X���<�d�ik�L��<P2Y��%7���-<�_�<�:=��I�nu�X%��Y�h�P=s1e<�G�;�?<>(׼C<�*�<���SƼ![=�%E=e�C��*=ݨt��~=x�t=�Լ�=�m�<4��%=0���=�^6����<0PO��0�A�1�l҂=�b������a��<�.;�D=��=ؚ[�$��86��<���;판�]A`��dt�e�.��/��B1��Ŋ;�O=�����9r�4�-��뼼%��<;?=�:R=eE�<e�<h���N��pŠ<v�P=Ng����a=H�E��!��`�M��<��+"˺ъ;���<
��<���<��<�mм�^N���g�h"= O�<�H=�H�0��<v,?��J�=��$��'���J=eva�p䠼�7u�(��<fB=O}�Z)�<Hr���o)=��R=�����D=��m��$q=^��<�2�yW*�Y�f;f���!G�<;rP�S�<�Y�<>�F;>��z��x�g���6=�g=��B=X[��	}<��lw=u�o=�?>�h3<�R��L���<;���ܭ�<���;�f=d6=��;��T��Rk<¿�<�
�<��<���^��c2=��< J=j��%N=GW�;�$u=7Dc��9s�z�g�<Kl��#@�(�N;45K=�4�Wh�<���8�b=�E=X����tl=~m��T�<�C=C�^=a�&��l�
�<k,��ݼC*c;;��=[�;!�-=-:漐#��/˼<�xq�7���	.��z𻇹�<b��<
�~=&P=$\p��5M=��R=+q�<gD�;�-=�$�c��m��j=s ><s��<5x����%<���<��>�(]8<�f�;�Q���4�;�rB��l���ۼ5�%�@;��Go�����<�ؐ�y��<N
=)�A@�;$e��K�U=�)=������q�;3_<��<+t&=�ԃ��9~<t���z�<��v��f%=rB�;�d�=��<b�9hi�<cG��qo=cp<��{��{
��Mۼ�����Լ[�мZ�2<
�<pw���&= ��<𮐼b
�@�O<SZ{=�T��Ѷx�I��fy2���<�%<�7�<��g<`[<�h��S�K=��>���l=��|�*�-&N�4	�<}�Լ�<��o�o�=Y�tۼMR/�}�<,�8=��$=�tr��/2=�r<N�;E�<�M=^.U��nm<��v��lQ="W"��?=���#�)<6��<�@��z�(���^�~�4==�S<��B�wܿ<���<
"<��;<������c<X��<ܥC=����T]�r	_=���<�=�8�<)�1=Ӧ���6�5�?=j�=GDh<讻;����o=FM
��{=G@��?��P<�Q���F������];�'D=E^6=�7���9�<���~�6<?eN=�#9�M�&=��^=a`=�fr��<=0�q~�<��v�����
��<��=`V�=���{F��3�<=�=��f��qW��/h<?C�䔗�Gc���3＼�&=��5�5_)=OM�<f���|Գ<)^=S���� }ü;�<O,=��x<� =�.>=�+Y=ZR=O%��X=��<++a��lS�~u��Έ(=�˼s�<=��)=�T���
��=@���똼N�=��H�<j�=�?�CF�<���^����Ͻ<��ܻ�<c���*���t:=��<�n=̴�<����^�<<����L=��O=�R��R�wٍ���;R���LX=aX9=���t�=�=ںGt��4!=�䎽��B-
���A�$U��cO�H*=X=�=����D=9$*�WI=��K�=�:J=:"=��,�Q���É*<�]�<�\�u1���-���~r< �Z;�\Y����<<:r<����G�"��DL=�vc=�>�:W�h;�+=@ZI��X=�dW�ϊ�< ��<ۦ$<��Q��+��"�_�B�&="�Z��:�=َZ=��Y��QW=�H=���#X�Bu�P�1=Qp�k��WU�<2Q=Ы+��k<�A1��ke<-F�*���F�[=�=�R7�W���[�w�6����<OOq=0F��]��<����;=^�M9��=�"=�Lp;`S=��C��L�N+s=�=Ѽ�f�����њ�����W�ѫH�����,<�{�#;�=U*=���<�H%<Q�<b�b���<8�<ЙC�;�</XE��{=YH<��R�[�s��M����{=�%�������4Ț����;���:�Q�ڤ����g���<xR	�&�0<��<��=��Ӝ�#�}=/c=�I�'@���U<��L=唼?O�<4=<��ƿ<c#��l=%H�;0���=/Zy�s�w=�f�d���p��sT�y,1�G��<�5H��~�;��$<m�-C��M�;o�ݼ_����G��fB��ג<�/���*��G�+< �K��;� C���[���@=}��<��#=%�:o��<�$ =��o-=fn_�u��/TS�^$�P)���x�h=ܵ>��g=�[�<���6��;�59�~e�]��:�E=�.L��,�ɔ�;�O�TT=%�f=;S�S̱<?1�<� (�s�"�7�:�5��6Q����}��;��t:����N�P�FNd� ��<���<�"<-��'���B=a�Q<�X+�P�~:�69���λ�P��� >=����,�\�ѻ׵@=�  �T=ͭ?;���;�0��D ��/�:ʋ=�PA�d`�1�W����a���Ň�:��<&i=3Uϼ���;��,==���=ɓ=�ż(^)�И;�1r���_=T�E��~��$��J�<eG�;׼Y=�{Q=�\߻��/�C����ͼ�f����N�u�<��n�X@4�L���$��<��H=�Z���]y�N��F�N�ފ;=�(�/��6t(����=�AO;���<��x<��=1a��H_!=�m�<Q�a����<0w�<1w��&8������M�N�<����]�Å�;r��=dR=�pg�2Q=�p%�{V�<Օ���f?�b�<`q$=ǝ��j���.�R�����ܒ�<� e�	�2��Z=k��;IcļNż��<C�[���ؘ4=H4�w�t��o����%<{4��PA��. N�-����-=�����;�N�;&�<�+��ȇ���z=�T���n���+=�{=��d��C��?)<����<HH@�4�<.Ф�F�==��8��d;�L<�V�;|%=y,=�|s���&��Wл�F.=�Q��0�3�J=��ڼ�`g��׸�k�S��������?=/G=)<�|Z<�g�<�e;��
�kdd�҆�<sR(�����U=UF��M�<�<'m�;?l�i\=)n;��z<�����7�����Gj�p=�<������A�J�=aBH����<ݛ.=h��<���:�Si��
1=�jb=��/==B��B=G;���/H��N�Cs:��H��<5��<f_�<��I���=Ƽ�A��Vll='�:=�UG� =-��9Z�?�D��<�n<S�W<+nI�7Aܻ���<FC���E<���;E=ǊB=���<��c=��p=�9<2KC;U y<��y=4_��=8Q�<��<�ټ%3���|4=J:�g/�<Gd?<�;���F<DV;8���>9=�T�<6�<6!$� <=j�<.���%+�=�#5�d��;^=�O|���3<X��<ϼ�<&�^�<b$�Y�Z<���<,1Q���h��:A���M<��<1��:�v߼5�<��<�%�=FN=����Ņ��Ul�˖�;�|�:0�<�;^0�U-,� �=�_X="#�<�:"��}��3�����7B��a.-�u��<4[�<�=�����Q��b=^�a=��g�����q�}�;�>=�9/�����Y��5?�6�|�ne?=�ޘ<�<Dvün�\��ؖ�C���%v�<��9���I�t� ='���S�-=��j<f�9b�����<函2�/<l;�<^C��������l�l=�޼d�����<�S�~=v<<c[��&;[J=�	�${><<	�<I����b��V='�D��k4;oA-�͇���� =��;�����<#�Ǽ4�=������=���<�S5=�ۼV4N�n�<RY���n����<�I��{ƼJ �p�!��'=�79�r����t�븸�XҞ;�(��/��;���<���<^$�<�l�;g�e<��@��%��.��љ;�0Z���]�T�D=�漾�.=Yg���w�<Ã<�w=2�`<�'／{�<q(=o<mM��@.����v�V���J<� =�dW��O>=�UY=� K=������<���md�c�3�_��]�F���+=��|=�ǚ;�㕼��P=Y���~�����<������+Z���������5=ʏ�<�lV��I���PP=�{���<?LP=��\=Wӱ�1bS:d-%�7^]�6�-��)K=Z��<|!���/��PM<���֤K��\��zP�<.0=��}=����f�'�x��B���7s�)��<� <�#=��!=���<�^�<����<��)���E���{��A:@;cl�� =��뼟�X=�r�<�T<��W�Kթ�A/m���K=~Lp���zpϼ�{;�z=U���Z_�:=w�������1	=V�%�$�ݻ�O=��'=���� ���<G���u�b=x�=���=���<?A��ƻ��<��hE켡������<m:S<@O�'W��=%=����!c����N=���Y=~�y<P=\�q���9V&,�>Z��m�6=Bs���=ߕ�?�p����<MT�;�e�<V<P����?y<�ʆ�:���2�:WpQ=��;�9(�<i]G�WAk=��ż�F<�:���}�<�\��M�[�0��;"�_<g�=O���?�<a2h<dǿ<Y/K���U]���:���s��RN <׉)���$=��%7V��mѼQ�E�\H�1��qҼ�~��:`��$=�=Yd=*
��)� ���E����<�I�<�	=7�7=M�L��-=ϕ��	�,m8=�4�<)\ɼ\�����Ѽ2gh����;ژ�lw5=��Z��M ��<-��<�>M=�<μ�,=�Χ�}�!=~HW�m�v��a=d
H�~׷�36�v�=hN`=�诼F=4Q�o�,��m�;^X��s�<���<70=��<����ϗ�{kv�f��u�m�ԗ=N�<�Kϼt�=c:#�������9�͹�lFk�y�<m��V2�*6R�P4s=�����=]��<Z]�<w��G[��"/�6���AJa�a��S ���<��$�<A͊<��t'ѻ	��<Z$H��&�ak_=eڼSM=aH�<�
$<H�<9���O���ּ�4= ,�<yX��VHm��!伳aI��nd�/6=9��<���-�0=!��<��"=���,�<�ډ;:X�)m����<��C<X4� =*=̢�<B��<�T#���;��� U�BI�i�$�����w?�<�3����=�J����;�~����[�u�s�<"���S�<J9;<q�9=�\$=��W=���<D껬�=��z�1���=��M=@D<��>(����^�=e=��<#�9��伣�a�_�<�m�<e�Ƽ�,=w���=�t=āK=����C�;�R�~2i��["�C�c=%�<h =+.�b)m=sGk��+˼`�3�!�D���<�&�<��D�Uq�9�t{=U=���<C�;OdG�U�&<��<���<f��8��<������:�#�<re�;�(�G툼k�G�_��h��4h?=���S=��<�(q�tyU�[l=-�=��	�����V���wdb�15Z�o=S��<H����?���x��e��Q�;2�<�5o��4=�B�<�m\=;��<�< ߢ<L�N�+�]��+c<�=[e=A*N<g4����$<��=��/=:���t:�_�<u=u,=��>������w�<aA=ΐ�<̷S��a=��e=�;�<�׀<{i�����=�=޼ J��:�b��3��(2=��L=9����PK:¤N=�r����<6�@��
��k& =� C=щ�<��+D$=��o=ʍ��t3�<����;.���<Z$<=���<d��&A\=�S���<Hӻ
R����������Kq�<��<	V��=4)�<�#����2�H<T'=�"���<4 &=�(�9y"=/�=��s<�8=���<q'�;~d=�yk=����f=_�%=�K`<������ͼ*JL�bd=��=%��#h=���;�rR��� ����<�kP=<f��l6\���l�S��1�;�+|�؉;�%�*=����Ajd=�p�W~L�A�0�}�G=��N�E1�>�<z��<A=N	R��*���vd-=a�B��x�<�pd��L����2<j�D� gT=7VM�>��<Q���0{1�}n>���W��	��E���=��<�/k9��{�R	)��L=����;=b���j�V�~<�	ʼ�`;�m~��%=�
�<�qܼ����D5=N���� <�/ ��Ի;l[a����<
��<;Sz����_SI�iƛ<�&O<1���,\�6�X��G�<+���M���������yWV=��<�	=��m��޼y���z����J;�b0=]|<Or=�.ܼ���<�ޣ<cd�s�)=\��<ͦ9= �4=�U(<p����B=0%�;""�s�I=I�S;�5=3�==1*�Чf��O�<�ϼ��m=��+<���<���Q1�ǽټi���� =��<)Һ_]Y=�Q���h��t=��<��F=0�Լ�I=z����/���;	B=h�|<F3� ~�<�:ټ��E=,��ۭ���r:��{S��iW=�TP�X��<��<.�e�J-�;1��[p�;��'���^��1=p77��v=�z�;B�ֻ��;]$㼗�=l� =�OB�ж'=�����@<�H�<C{I�P����F�QS)�/�Լd7=]�=W�K�<^��0S=��ݏC<L)�<R&�*�����̻�M=ЦU��[p�ߥE�:�Ļ��/=;}<�=���<��*=:�)�r<��A=�.4=o� <v�&=���<�p�0a=1B��I����[=�*=�XN�'����7���M�L5Q��b%����<#
��̣<D��J���?����K<!1��.��Nʻ�`�:�F�Z&�<I�F����:��Żd���슼Ε�w�� =����<���k=�#$<��L��O���(:�]><Qr�����<��+=D�����O��<��<]h^��6<� =I}�<h3�<$3��d=�2=%G9�y�-=z�V=�;���<�愼i�T�h�l���%<J�w�<�l�ΑP�'P����� ���Q�}��W �<��i�`:=
�.<��	�5�Ǽt�<=�f�c�弹ʭ�_�<n?p�zB�<��3��U^�	�<=�x ��Z����2=�(B<Q��Y��<a O���<49b�]q<�Mv=�U�T�5�]b=�����X�^�/=f>=ZQ1�/,R=�^;y�[��;��=X��V�4��(�����+=��G�U=�B˼MV=#,?=��9=�L�<�1<�|��<����Ͳ�;<�<p�=�C=��8;����ѓ��T=���<|G
��=�=�P=|��<���F=��<[�����;��=o}(=�"���/���g��f���!\�����Ѽן��	���Ӻ�<6=�=�<@]\� 1*�|��SI=���V��R��"�oT����<�|S=�ƪ� 2=�
��@={<^=�>�@yW=԰�<n����뺼*=���t��;�i3�Z=�<t����_{:GQ%��ׂ���>=�->=��P�C=�� ���,��sz;FἚ��{<Z<)��;z� <�����C�+�=�_����m�=���:<ﻄ����;��/�?w�<��Ո�;0��<c��r�r�7=$#d=�F�����P=NT=st�:��弢f<z<=} ��[�<mρ=�q0<9y:<U���7����ؼ��<�ޤ<O�(��SH����<��^�k�<4rz<B!ؼ:�=�#��D=/=���<ո;�����=:=��/=Q�l=�VH��i=@���}x�ɾ׼q�=:=�ف;��<�����<�p�<��Y��9L=t(=.ʂ=�'L=�'?=,F(�UF,�������]�<�����i��뷼��<�l�<T��,@��Ӹ�x�k���|�_%�<�b�=6�;=V����g<�C�<�zN=%�3�\�=��<���|!=f��=W@�G| �L�ϼ�{�<	����?�G:]�=y��;~}i��C==T�a�[��;�g�<�p=��=!/�w.5�dE���	D=�V(=��<�΍<�j���Ig=��<j�==]J���=!��t@�<��=:Y�<�Ԅ:��2������N=����Ti�k!�����?�D�$0�u]%�YS�㊼�4<��μ��U�5��.@d=;�������*=��C=b���7c=�	=��b�\=;uW�)�'�b�����'<^�7=k<�W�<Y�<�ۣ<�6�<lJڼN��VY�<)}�<�*i���(=t�z�P��;2D=K=ۄ�By���R-�wג��,�*A��7x;T�����<8��<�i�;����D��%�{�jW�:m=�����o�4<#�:����3�	���\<�� �]�;]��<����U=)�<(tO=�w<6B=��uE =��W=�����K0��܈��O{�#�U�Ca�;��q�]�]�h�@=�?ؼt>*�GM=�@�;R6�<�mM���'=���<J�;�`S=j�<W�<k7i���'���7<.���-=� ��w�4��n�=�(�<�BT=t~�oj*�.*=d���
x=M�=F�Ǽ�W��=/�;E�v�a�ż��c;�І�-WT�녓�X�)<�Z</���}�;�@w<���<�7����<|���s�՘��M���=�	5�"��<���:�=�=�V�<!N�<���I)=�]==�� ���	�U�o�U�;0TL��'���<��<}�<8��<iq#��G<��;K#ۼ�Rѻ�ja=]<�ay��5<��;l���j��e��)�n�~ɻ�X
=h��[`ٹ�����A�V�F켚��;r��<��%<�]ϼ?����!e=�l#;� ���'=�rw=�μL*Q�}�;=�<�!�^	��m+�<�v����4�?��<S��M!6��.�����=9�f=+L =��¼�==�H�=�<�8�O�^��_��~�<���(�=�D^��Jm=���x| ��C��̉�C �+D�<�n���R=��\��#=0�=~�=(�������DUv�������j=�.=����5�=�5<��<oە;�6/�`�0=o=�6Z��V�<i�Q��+�;ID��T�7�Y�&=?'���;�M�<vüˆB=�S|���<]oj����<�[0=��<ֹd��^�=-=�O<�SE�S��;������@u<}��<�@����4=cv =��P��,�<�M=��;!��t�����<@�u�����}�,�����#����μ&�=Ĝ�<��#�O�	=��}'8=V�f<ϫ�<<�d=���>�;{ep;U<
�Y����<c~�<�N��BS=1"�����������v�<n�<"`�<u
�<8��<����;=	L�<"=�E^���_���A=~Q=!I��T�<�C�7l=}����#@=QW��$��Z-�<��ĻGv��誼Dȼ�-F=��_<��M��w2�{I��;�]�<��]��&:ǭ��KM�N^�'�$�dO�R�l=O��<����<b =�P�=tT=��=��Z=�H�<�*��B�-�H_Ѽ��<��<)6N<�}[��a9<�x�+Y[��7=��<������U�_�����<��<fy���<!ռ��<�ۗ�z�f�&��]2z�2����F8�Af3=����q͓�;�=��?=Q ˼��<�z=��<�= ��E=�0r<�02�s�"=ֻ"��
�����]x���4�n<�<������b����@�pӏ<f�E<��
��,�="K<|q=3�q��;=�J��J�E��ݞ<�W�;�H"�;7�m*=6v�<r` =�iQ�4�\=Ѫ�<~/-=���LG�`�<�Q�8�E����<����V<9�'=*EL��t<Q!=nt�:������.=��<`'���B���i��o =��m<�e��q���<�E�t���./<qܼr5��ď;-�����=��H�(�$�N�<0kk�X$���ڼ�%=�6=Ũ��f
=�	=�~�<v�;X&=C7��
l�/꼅^���¼��=�@V=`R�z�=��f;W��<a%�<Ӎ��k/�~��$H:(y�<�u�=��;~�a<W���zr���*=U>�<o[�w_!�.�+=^�;{�|���C=�7N��.*����;M��_*�=�
2=�X<�&�G�<�="=��f��j�D�<�P�=&��<���<JCO����<;����A(=��2=A��b*=tY=���,=��=���<-V/=��=�n=N�=�qg����&E	;.Vu=("�=��^��#ԼI[��ϼW29��~�W-<��<��<*$=��}�1�4u=�~/�=���ڜ<G��9�ޚ��Rɼ�eP<��3=�O����V=`k<)��<�OF�������<F��<�(l���7=����as�?���;�d���i�<0�<�qr<6h=�~�;?$U�9����MG=]lM=V����
=k��<μm<��<Pp�;cY��4<hd=�$s��p�<Z=�"�<�1o;�¿���"<��4=�-_�Dzq�^�=~��<����bLּ��.��Y��:��<��d<7�+��<<?=�&;�w�p�<��;=�p_=���&ը<��߼�!=�F3��b��=�p���q�=5��<0�c����C1��8�<���<7�=�rd=%;%��;��?�ѢZ���=L��=#��=��;肽 Y��_����C��M������<׼)�њ��x�A����:��<��3=��,��mP=PvF����cmk��c5=�_=]$K=}ۼ�`�0PF��댼gt���%��Qj�H��1��U<M=�y`=�A���ީ��z��K �;S�=�jC=fߘ;b�y=�VG�������!=r+$=#ذ<󈘽�d�<Q���=��"���@�v�ݗ�<u|����h�WY����<%g�ǅ�;�?���D����;��k���:_��<���<H��<�6�w��<|ݑ<%��<5oE��(�H�N=��m�%Ȩ<��<��<|�i��0�<��:Ư�:9B ����w��4D��_l/:�1<�3=u�@=�;B=�-i=�me�6ƃ�ծ��eg<�������Q8��w=��;/��A(x=���;j�9��*�d�=���h�<X&м4 :�v4��J�����<H�l�ç�<�o�<��<�߀<#^��L:"�&ҟ<C/�<$}���ܽ�@/G��>=�l��z_u�N�U�ٺ��n=yC���P=�ݓ����!=j��<�X<��)�9�����x��w�g;�M)=���<'
�ͣ���7�+v�<�4}���=�&���B<[�	��+���5B�y�W�bfF<*�F�UA�<G��?Y@=Q�&=�b�<u�5=ze=��5���<��0=,�8���1=�\�&h�<�#&=pg�	�=��#�-��=���<U��2�:�1A�	�3=}X�?����> ������5=z4+��I¼�+�=�G�:5CE<�t�<0�����:<��a/�f������<)�]�S3u<d��:�M=r��{�<U�=�.���;�5@=���<�=�<+1�;Wh{=^��IS<S���=�<�7=��ͻ]˒��L�<�ܱ��=xW=gμ��E���)=#x$=;9:���H<pN0=���
^��P=��=�����P�x�n<�~B���.�6u�=��A=%ټ���F7�<�<��T�=�4��k_����<mz}=(�ѼC�ü���<�Q=�Ʌ�m �<��M<'}�Ŷb��6�;���<8�'�W�N=�c�<�l;�Y=��<AFg��˻�^�=��;��<�Z+�Q�_��=�Ǽ �=Ո=��j<��I=i�:,=����m<)2G<����eeͺv�-���U���$=�U�=L.=̀!<E�!=[�����;���"��1�;�c�<X?���U�n��xM��ZZ��s=���=	r=CL�Q�v=E'?�����ۼ�<c��`�U
=Q<ڽۼ(�S<���<��S=����@�O�;����L��>=BǼ��ܼK�`���<��;�9=����T9�8�J�4:=��4����V[h=Iu=K}'�k��`SL�r�뻩M<��)��M�]aM�� ==1�=�� =g� ��8B��(׼Ɏ2�0M"���[=�R�����¿��ۗ�$�b{���Ǽrm<�c<,o<4V�˼;����!��m�r�\<lp�<G�M:��j��="�@�-�=�~0=+D����<'��<�d����<4ǝ<w}2���=&��=v�������4=�x�T=I���4=V騼LC���c��CB=�5<�L���$�g�I�.G(=	&�t_=�}}=�|��RUR�e�Z�Q$�:}+��5EQ=�k9=����#�u�<��<�q�J/U=�2��U�����<�HF�g���Q�y�W��<5�B={���@�$1�<��`��<�lA��x�s]�<��i=̐y=o��;��g���<�-���|�G=��8����6x����P��8*�P�<5E�W�S�&�Z��մ�Q�5��=����r-d�e	޼��n�"�`�`��	�<Ø;�iV=�����3=lƹ;=�<
B=��^=Tj�;HID=C��z8=�N= =�<ӁH=8�W:� �	{��G�|="R����<�[c=�&_=��̻�<�v;�9���C+=�8Ǽ��Q<��Ҽ]H=�&���[=x�}<3�g��u{�Grؼ����D'=�h=(�Z=2W�����\+�s7<R��<{�<������9�c�Q�6�<�W�.��t_��A(=��G����<@��;���R�5=Vi����ݼT�A=�V��
�:��k=wV�<{;��7�<�E=�t1<��컏�5�����,4�;'�=�O�G���-|�0�*��C�<�y,=?*}:n;=��%�c�b=RP(=Xf����==K}�:r��=��C=�|�=�1ڼ�́�ǫ���Z���k=��L�O��Sy� �8�����,<�l]=�5=o���
�bB� |�9�Z�mM���q����gY=iq����ռ���W���"=(�=�0;e�.��=1=˺伜U�<��<3�Ӽ�k=B:9��ۣ<R��<�d�<����3�<'{�;���RH=����(.=��V��;Y�g�<�uJQ=��P=JLE=l2�	�4�h�=)�=\�Y=�V#� @2=�m��u� =^��<_��� a���B=�a5S��~
���h��ds�ݳg=#r�:>{��7*����H�8�]�N�&-����7��m�����&=q�;t O��4���b�:{�T�b{^=+�8�-՘<ɤ��U�;B=[=�E�=�`<���<mD{��C�K�Y=o�O=����r������<2�U<d&X=|��<Hr;��<s?�;���=q�a=��輠���Z=��L��=��>=�@J�'ƅ=2f\���5��is�%G��S)�=md���d�ޢ?�7k"�	�W==?�;���<,�#�=���<��e=��*�@��<��=#���V=AT�<E �;r�0��U:<zBJ���@<zp=J� ��c=7�4�j�%�ӭ��><�ûPLN�|�x<��̻���Rc=�qM��L�</G�<n�R��.(=���;3=	t�<�<SD�;�.=��R�+n=�	s�V
���������%��׭=�	=x������>��;�cF=Yn/�ټ���<<�==�#��/=D��;�����Q=L��<��ב6=�<^<���=�c�=�׋</��E���Gx���Ը4�+=��<�AA��<�p�Js�;������g=��<l�@�i�-�]��D8�;�a�zf =�����<���<�8Y��*�<D]<]��;! 8;J+=�&�e=��[��y�<΍w�mG�:�sg���<Y�y�';�T��V<�\�����ᎆ��4x=��j=�0��:dS<�.����~HZ=�=��ͼ�}�g�<rJ=9�<m�Y=��`��Q<��<�X�B��Q=�E	<��!����\���	�Ά���C��:Լ9���^=���<5P=<l�!=� �<�|�;pݼ 퍼�&�6;�ZQ=;=��μ��E=C��zn�<5��v�[=��h=v����Ảt=,!D���G�<�=�W<(�r9�G8�ge=
A=��=Ȗ�<�����;�_�;��a=��-�cO�<�_�g��<�p���O��7B�����5!��������d�j�Y(P�݀���h�=+�8�S\=.'=����]5�J�5�]�;=�G�<�+��룭<u�P9o���y�<3ن�81��,����y�є�����;��X��B�;��<�l�;js�<y�;8D�F�N�=����f��B��<�1�=�|����;=�d�:_(�<�;G�h=5[�<�.ļn����@;����.�&=�`=�5}���=�x�<�C;}-�?�)�y_;ȁ����<:�W�=kF#�����ۓ��r}<��<n��ɳ?��?B��޼º��T=� J��� =����=�4���<E<T�=E��;���Ƹ?�4��;�У�!��xպ���`�&=Ţ�<g�#=A%5�0=�=%w=�[=M<{Ǩ�9<м�)�<$�N�ڝw;:  ���)=�U�tU�<�]�<��2<�����<#�<�r=�����9�n<e�F�yM�Jڐ<��=@���S���<μK�L���h���)=,_<o�G=9|�"�;��<������p�lչ;�V)�[K��I�@<`�b�M�X����;P+�+9�=1=E�����I=�Xy=�=Q)Ƽ�����
����<�q[�
�6=4V�
�1�Rw��6�<UJ�{켗�.<�r:�*�<O!���<"~T��" =#5<��M�9
�b�=�WH�P.��DA���B��љ<M��:�_�=n��Y&��g�E=q���r@=:K=��=?z��'O��12=	:=u�,���S=	�%��-<T��?�=��w���`)�J+�<�m�<xoQ��� =��m�l�P��pv�J��;
����[!�픐<T��;mZ=#�u<��)=܁I�aMѼʠ����e�*H=��/�)� ��<��ƼŲ���U=pfi�1��<�m�<u�h��#ʼ�A>��B=��4��S�̼�C���w�;��6�A��.�;eT�a�/�Xy}�=����p=l�R�X�R���= ��H��<�,��2��ɸ����zռ��n�6=��I=^;��{=�b�;�2��'n;��<�<�+�;�=hn$=?0�;�/h=�i��c�+�4�;b�=%O��m =���&6<!	��]�1W=�]z�Wc��F�=%�m=�������;N%�3 =�JM=7�:����[�����<'�,=�<8=�+=Qg=��/�_%<0��<j3�2���y�a=��h�6��;��û��<��b=��ӻ�D='�#='�r=ˉJ�p��<b�=�8;;����<j��z=�
`=aؓ�l���H��=�u=%0X�K�r<�u�<9��V'���J =���;��м��=���;����H=<Ȋ<(1;��%=��=�oL<<��< ��<0����2K=գ=j���o =�")=5|N��B�<za��7�ļ�2<��>;߼2����31���6�fN�<�	=;��<��<2�&=�@��U�9=�p���@�� =��޼O�����;��<=�iI�<)�m��e\<<֞<=F=��<;���<�=�v����<��[8����<"ĺ�r7=��1�u��<�(�<��X���<~��<��'�q��<����؉< ��F{4=�L*=܋0��s<o�=�G
��R�~<6���33=8�<�F�B�������\��q�<X�<�¡~��=Tw\�=I<k�+=�~Z<���r�.=��<��5���g��mp����<)�=���< �������H=�d�ぽ�d;�q�<�v=�s
���m�ܼ���<�*�N=�Rd�}Ó�{�:��p�:�s��S<��=0n,;ETۼ��4<��	��\i;��U=+�'��8=���<{����0=�i�!��X�;��
B<eÜ=��G�m-=��m<iֈ;`74<R��y*����7=d�켿T��B�Ҽ�Qq�ׁ�����+�<t��<\��;�r=�r\�gjX=�87=����,}�<�&=��ؼf?�<��= �����P���:��<��=�=psc=^d=J�_���鼍�}�9_�[A�g�m=�M=���^Z��a�+=�܋�i����\<^�:=�`���?�@�j=�'
=�3�<��}=�ġ<��s�QH��0t=�X*�4�x�Kmy<u*��ٻAt=╔<�}༪у���!�W�R=�&������0D�<#[޼��,���;v%E=�x��ӛ<i�a����Ǥ��&!h��=��������g+�j_5:����PԼ0��<���<9̼L��<��(=7==b/<&�P����<a�r��'�<�n�B=�!A�h.<�����tL�;�w%� g(�`� =� ���+��*0=C�Q=����x�K=��R��L0���7��rX=�s���U��F�֣�����{�ӼK�<��ӻ�%�g�<�s5=��#<���s@$��)�<�;A,=+��<�z==C7=�?�k��QJ?�5]_<U?��/=��<�f5�@c&=X���2�0r�<2RS<��Y=��E=��Z=��=`�W���2�����3G=�><�o�<j�=;�1Ǽ��<�u��<ֶ=��9=<O��q=`�:=*��<̹弄<�=>�ӻ&�ü��*=��	=��o�.�[=3M�<o.��)�B�m���r!�;����� =D<�V_q=���<aTA=�C%�N�U�x���,>h<Cf��[P=����A��ѱt��(���=���;��Q�o �<@�w���#N���Y(�����;X}ռ}G(��/N=dp��
};�x�=ی�<X���oW��`�<�L=�+���{)=3�;1�%�=ek<2%=�N�!d�����+�
��ɮ<eS7<vp:�rz��1�G��'=�5<�v���ʻ~�e≼�ᑻ����; ;X�=� b���<����<�l8z�
;	;�b����j���e<��A��>
=�����<�;����~����)�Q�-�8��Qr!��Se=��==�`�<J��<T-c=�M=s�<��=�V;� =V�+{�<�r=�GŻ���<L�<V%�; &�;�缺ݚ���`�U��;�[I��T4<h�=�%=,] =��<�9�<��e�N5=�����<�I�;s�@�')`=A�_:0�8<��0�QzY=WB=0%W=�b+�-��<��< I3=T�<`�a=w�;č7��|
=/�&=X��<w����)=*��<Ou�JY��Ü$=gP=�&E=3�{��{[=�8n���f�[��;.�p=;a��K.��(�<Vq:��@輇D�;��6=j�W���=�%�<��Z��;H�5<��8�"DF����<�$��q,���x��;�#
�斐<~ ˼!څ<�	�b>�m�b=wc+=Pa�!s��[L��eN=��M=��z���L�?�=������<,M�9�1���F���<|���1=��w�<��Q����x-=���;�ƻ��-=rp?���.�ae;�Ho��2�0���|<��b:�U�������;k� �����<��6�I�;�J&�A�3�bؼ�r�w��<�R.=ɓ<gXi�0:,�~#���b=�z��.�G���"���~�� A=����<_��;�b,=�@�t��<�L ���,=])�;X�o+&��B��(���C�<}/ټ�;(��<�V�~uS�"R=��%��<l�S=��<������w���}=��=����ۼT�A=�����l/=�CŻ�U=D����8?�V<���K=��1�.��go���H��&;El^=��ڼ���; �<�{.=�**=�;�����:����˼�.#�K=n=&�ڻ2�<�w¼��$=�e��t�Y=�g���?���<�R~<����&�f�;��;fVD=����y�3��Ǌ�����qV�5Ty=���<�<=�+�<]�"��'=�:J�4���f���#�;9��<����$��_��ѻw����3��G��S��b&=�l��2��</��<�{��L=R�P�Ӝ��˞<G�< �0�^�=���<	桻��V��o:��l� �6<a����<�"���$�<�1D=�x�cx������-=sI<��)ƻ��ż1p�<)Hw������P=�9�<��=j���$P�<�&�.9���<�	�:8ܼ��<i=�����;�a�=�6<���<��<�y�<�z=�y ��=x�0�L��(�M�`��'P1�]m�[�=��
���"=[�E=56[��#<Kw&�����~#�k��<���Z��B=���Ia�<4߁�A����S��F��6=l� =���gK��vT<7�@<�Qc=zR���"<k�$=�"��`:���VP�m\:��ӻe!=�->:a�;s��<�!��s1�"��;���<�w��F��wi�<��Ѽ�\�1[G=�PӼ?$U=���#p=w��,|�!�#=��ü�r=���^��N <�*=-���;�U�z�L=\���=�Ƽƚ�:(�;�E
=C�(<�� ��<j�b���@=l�2=B=�w�͋�;
�꼳ի<��<����A�,���ټ��<���q4�S�<|�c<)|ּs
C�u��<�j�r M�[�K�]K=��<U2�<��0<43�<�C:���!K��xYɼ��ȼ����$=Hdj�P�9=��<�<=ݔ���I���>�L=�q�
nN<�8ڼ��Z="�����7��D�T=�=Q�a�����Ӽ�~5�0�<T�˹�:2�B���$ė;AF^=�
�;�Q=�����=�+7�C�)=�F<[=B��������(#�8cy=J�~�n�y���<�A[��:�<���g8X=:]=�e=�΁:�2��ˎ��@��tp��{�A=��0�i��y�@�{�	 <{N�:�_�^�n=��Z���	;6y=����Ũ�ќ��iM=�R*=��'�|���x)�}T;�7=��T<"��<´Y��F��,=b7G=c���(=E��v���'�?��<y����s1=��ln=�=y:��~H�N�3=�[�<'8�e=d�<���<�+<Ρ�<��#=Ğn<�TQ=�Y=��|=�l={�,=)Z=|��<�q�mT���~�ˀ �>o4="���K��ķ�<��<����Pk��/�)=-��<Pc���O\�ᦫ�/J�;��2��]�d���[2=l�t��{�<^]�˧ӻ������<-�"�Dx!�$Z=	*!=�#�<�˩�P<W��xѼd7d��n]�ȫ���V꼿YY�3�<g{�<�ز<�L;=;�S=xk=��ּ]4���ݼ-e'=�N�<W�=MQ�3�&��!�:D^�*��<��<>��E�K=�褼��(�t1c���<E��<M�k���û[tE��ܪ�r�:=�e�;h�H���<�����<�<d�0=I&���<�oz���;$�=8�g=mk�y�A�e0j;�u��2�������Y=���;��<2r��UD<=�с:���<nU�'0��O =��T��ș<F�=�����;�U<��s=�n�</�M=U�X=��O�&��<��W��.<)�6����:���k���B� ��]���nB=+�-�>m��Ļp=��><N���6��<���<(�g���T=*�=�H�;��1E=sO�<#�g��y�;tPB��*S=֋)�������<�~5�y=���=�O߼�D_=�Uz��S��Ӌ=�%�<�0��1��1=U���ż�f<Э� ]��X�J�=���<�#���%���;!�;׎�<�Yj��eɼ��<��9�,a���	�O�<���A_��8ռ%
��X�$�G}=�-f<~�=��ڼ��<=�r3�E�d=!�?<S(<�R�<�OR�q��;\7=�0=L=sG=IøVSu=㧼��κ+EݼK�Z���	�<T=�H�<j��=�!)��MS��j=t�_���~���<��@�E=D���ά������e<
�t<.���3=�	y��B=�=��ü}�߸w]��y�<��\�m�:�K����;������"=7����[���O�;q�l�D> =H"<�uW<�����M�;5P:�}e�R�
=���;��Y=�[���x�1V����3��U.�O><��)=�R2<�jk<P��<���;f�]=*�8���z��;Q:l<Ȅ�^Q��Z9G�s~�<ug�;sV=�T�jx]�.;�i�{�-^(<�CC��#L=ݧq<
l"�܋�<�X�| �<�nb�P�"=@�n���<�,�<�;>\��=b���I=V�L<B;�eG0<^<κi5={u�<��
�1M�<(���s��<�=L�/<�!��˰�R�;<�7����=��U��,9���D=,�Y<�s�=$�<K�/=93;�:�2輇@ ;ts:�!��\��ӈj�ӽQ=3/����;�'=�P*��6.�K`�<�O�;��@[�<:B�6���.=<�*���H�]帺���G� �U^=���<c=v��<e�<�o�<�|2��(8�drQ�CJ;=q<�M.�+0��:����S=w�j=��=�V@=  1=�x � Df�1ɼ81g<N��E��Ugݻ�t��A)<�Q�<�n���L��@d��G�Q��u�\<��j=G�;�Z��n=$ĝ<D�=���<J��= =c� ����<쬥;��(=I���X=k��;�W=�;=��O��ԍ<��="�f<����С9�%2�<��>=��;'y�<��=k���o=���<����]n�_{4=N����k=Q�=Ӎ����<��G=C�
���H�ፏ8%*�Sgk�Dl�<��=:�V=��[�\O�;�,=Z�W=
�e=fY������<�= �#<W���
�<=k�8=a
2=��=Q���"=�E;���2=�<_�U=�O\=!+.���0��.�\=����Z<q؏=�Y�<7P=x��;'�i�x{Q�id;��.@=��	=\SS��S=ߤ4��i!<��Ǽo�:��<p�<���<f��m/�<L#,��s�(�`�/�|=�M1�x�9��	=�Sv�,�=N�{=��H�<A���^ڼ`�����<xNf=�$�;n���/����ܻ=/C=��2=2�1=J;��;��_1T�]�s=dh7��8���Y�b6�^��<�g6<�f7<X�.�q�=���8��<��<#aN�*�����< �"=�!����9	�����U��,����<��ּ�@׼�k*<�Ⱦ�%\=\/�;b�%<E㑼gC���b=�W0�8 �<��E���Q=��Żv��<]Q��j+�Jh=�¼pZ����U��<ӈ�d�&���;�ɼ������<Rv�=B62=@U�<�܄=��S���B�"t%=�F<��I�lĢ���
�o%g�\N�<y��;n)�<)$>=6ͬ<����o4X�����N�;��⼦�<.0=�$9<�<_<|�������d=���ګ�<��7<��<�7`=P-�p�M= =�g<=K�u=Y[J��Q=u=S=�qܼ���Mo%��ҿ��=�Z=������<� )=N��;UW=;�d<���0f<��S<�ri=�S=h{��1[=��?=��<��'�����?�`q�<ObN=�?��e���	=�6=��`���%�_^\=Ӂ=�eh=c�Ѽ�Y'�y+ �0�G����^�<z�O��k*;,-=*e:G��Q=�`�<��߻q�<=TƘ8;���L��=�鼽J(���(=́R<
!�/`�6{�)�&y$����<�ܼ� �{qJ<C��<I?g���;=>1���K���=���&=�/=�?�9Q�9,V��\1;��;!}<%�Y<�(���� ��M;�W��D�.GD��6��N ��!z�&&=hw�<g�s;+J���b=v'=Yte=]-R�O"����<-ŭ�ǭ�<%�N��l=��<�Rf���=:6��[=��/=l�G�HG'=O���=�˼�J8������Z:�?�8�����2�<�^=FI���#=_�=M*<!���PT=��}r>=W4�<�>=j�=������<B�=aٔ:�����c���N�l�=j�μ�� �I.�<0 )=��O�ݳ)=�Z�B�Z=o��<���G�;T��<i,�<��G��1��x^���a=~=6�X�8�
t��=���H�<��ºY.P=��Լ�	/<���ٹ@���<��D���}<���U
���R������=�Q=FZ�<�|E�?qJ�/{=�>:V=����A��<2,���y�tC=~n���o��0=��R=�}+��g�<�8�P<�5��$=y�`=�#�<�gb�T	��*=�*Y<K��=�zP=C�=/�=�i�<��Q�b�(j��� �<Oh����=f�3=49�9�M��9��/e��\=�!j<??g��w�<�,;���:��f=�K�<5����-�}	��TU=�X=>�T=�7��ٸQ��<B��<�uY=�C2=Lvr����:�0(�)��<��+��ù�s�
����<[��N�@�n=��1=H��<�+=�ԕ��	g�@kq<�;<Z����K�<7�@��[<ʠ�:l�<���<��P=ۗ)=�dO=.:e���&=2��<�o$=o=y�	�&�5�l�\=�����d=�?"=�o��{5=���= I���:1�=V���(?�	Lv�.���3I�H
�<E�<,z���`=;�9=Rh�zLX=�G��)�=��&�n7üb���X=�s�;O ��L�;�������<�'5D��k����P=-v"=Nx�<��g:������J)<�q�<��F=�����{�Qv{�AF=@�x=�`=�F�c鞼1s��g=
�=;5=UIc�/l!=R��DV`�.0�<��b�����:�M�	�<���d=����<F~<�*��!�6����<2V[�Fi���\=�-�;4�<%I=͍g���K;�T�N:jX_<�.��f#,����� <u����J�:��k�<Qz�<��<�u� <�O���V�=���<jtI=��>�͝2=ٹ�����jp[=�J�<S�6<�ߓ;(�=�l;�=���q=��<�ͼ�xl=\4�< �8=���;�U#�u9~�J�$=~��;�jr=��<��;O�!�4=�=uf�|݌��H�8�=d�<�ܼ^�F=~`!�ḷ<��m���ټ�c���<��<��2<8�5�}wM<��=Xe~=��N<r�<�@J<��6=��2==m+=�(���t=Ρ2�[���ز*=&�_<��	���<(P0��#B=DK��*d��!��=��T��<D�=4�Z=4�<����1\��4K��-=iI=w�w=O�4=|5�>��X<��9<��#=ԁ-�e&��߾$���=�:��i_=����S�d=X���P"Y��1���_�y��;��c=;Y�����<��m��[��"C�Uq=O%O=����<*:�̬T=.8����<#!/��u�<4�ü���9nk=�k�=�c=4R=[ͦ<���8L=����J=k��<-\Ƽ�&��u�XI=��=�<����<V�x<5�<��<?��<�:>="����=08�<=@��4,I�θ���� �@U��%���λ��p=��<�
����V���1�����=��<��<ǎF��7��'3��5=��=Ċ��ԉ~<���z���<!��х<�L��-)�sNú���#<igM8����d���_��7��S��ԮN=��=I
<TR=�.=I��<�˻a;=qe�<u�H=�&�����2�C\=��=����Ҵ/=5�<u�h���a=�ռem��J=�=h�j<�̼c^ʼ��=�wT=��7<��J�f6�;��	���D=�T5�ڠ=�L<�6��EO����<V��<�i;��Q=��z<u�<�� ���=������MQ;h���;u��<�u:��5��A�;��K=yIӼ���ue<H�f�07q=0G =�P�<Ta]=�<�Sgɻ�l|��ƼPׅ��ʷ�ndZ=��<��N� -==����8=fw^���<8Լ�fA�嚘��:=tTZ�����`��<��X�T��!�߼�W�<��<�wa�6:�����<�^<xψ<�'%��zO<u깻��V�!�[<�+����l<���X~=Gh��ێ�'�*�a�إO=��<����z��N�)��vs<oz�<��켡l"=|��:I��&�=P==,D:9�JB��&)�̰<��F<Xm&�ȷ�;�����3=1��;�mL<&��;H�,<W�K<hT�<Q�@=ۦ=���p�
;��W\���Ӽ�n�:*�Y=����u=��e���l=�MS�8a.�*K¼ �x�N�.�k�<�����;=Z6�<Wo/���==[�=|SH=�%�<��"�`�»c�=��׼�W��H��
S�J�R�0�;D�,=�p�<PF�e�4�:"伵���x׼�@g:��E=�z=H��ʼʏ<�U�<~m =.��<����\м�/��9(=��=��Ө =셽w�Z=��V<�	��B�ϒ�:D�=�S�/�߼s��Q��<�w=M�
�6-z<���<Z�(<ǝ<�L.�I�<WG;&��cI�}��<�q=��,=f꙽lT�Ǳ<.Sq�I=G�=�,=������1�,�i�m9��5=�ࢻA��50l���:=�<=� <�T̼&_�<��,=x�I���<���<�m�<VnB�s�t=�N@�|�(�PHӼ�?���´<�c#�l����2ܼ1ѭ����� ���B<xT����ۼ���<�_'�{(¼��
�������<�P�<)Q<�Ǽ�W��U�Ѡ:��?�<�<�DӼ�1e�_^޼5�<W�ǻs��:�����K�<���)۩�e�ż)$_=L�<�u3<���<�f <�;5��]Ҽ��+�7=�e�<�!�d��<�!�<�-<�~<|��<P(M=��w�.R8=L<��0&=�9�;1�Y=�<5�XӼ<�B<̩:��17=R��;j[��y��x�<A09=�Ó��m=�=(6���Ԓ<o�I=BX��棫��Ip��{b=��=��lD<���{(=8N=�zļW����@=�3i=�n���p��4� :mC��~X=�)��=�|���v�;c[=΀�<��，8X=��=fl@=��6����<%U�������,=V�<��e��
=o <<6��<�N^=Z�u=�+���=��<��Q=���=����<��<뚼�
;=�e��T�Q���<aV��,6�;hVD��O(=ө&�@Fu�<<M<ʍ(���a�������D=8����<�Gm�1D��0Y�^��0�Gf�A�)=��*����<R]�Os���<V�?=�薻�+$��\�6b$<�B=��<<��n�������<R� =>%�=<=/�<4��;�=��$��"=+��:�g<�`v���:�NW=5
���3=&����v=�м�m=�%̹���a,�a^\�1H�=�G�8_}<b
-=Ηx<5��<��~=�:��� ����<ZR&�dqS=4�e�����U=�=��)q��k��]�O��=Xˠ<Փa��6�;�B}<S�̚<��=��ڼ,�;^R�<�e���7=�-�����<v������=Χ���K�<��=��<�GI=��=�����q�;��T@���c=�*?��v�<�P��<�a<Mν<��E=�o�T=�*�<��3�V�d���N=��;=f�&�~T���#������mi`=�i�<?��]z�<�����Uݼ��$=��-�����5.���(A=�&�H{I�=KG<lJ�<��(<&r6=FP=�s����>����D�Q=����">=?����ʹ;B=)t��Ao=�h�;��J=�X!��md�OD�c+�H\D�f9$�	ʮ��Ƽ?�<��o�����(��c�<�4�<�@P=n]�O̘<<@���UL��Q=i�V�O��l�)<�:ü!6�rE;��<J��<�����|<�oK�P�<�>�<�X�<Gy�����VU��5�(��=�0�:�O=F琽�U]���ź��=Ԡ����<π�h��<]X�<�/��=��<��H��:m;�g��������={�<�a�<�Em=�N�<���<^�"������<�>�u6=>�<q�ּ䖟�?�$�ϙ =W{{��h��*ʮ�2j=U�8<��^�{$f=ם��:)�	�=��6��C=�bA=��X�Al�<�g=��k�pO!<���$�U��FZ=96,=�QE=f��<�>=i��<�6=��;�����?�����U�<��H<I��<��2���a<lJv<�;�0�<d(	=�4=Ƙ�<5�����!����������+���޼�O���o@=)�b;��"��J=֘C�<5�<pG���$���?C<���;I��<�`�:cs-= <V�	=��t����׭<gvһ,4���s��:=j���l_�ln=�_Z<3��g)4===Si��0�<C;<}l��F' �퓷<�M�<D�=m�t<�L0:�=O��<�t����<B�;�I9=Лټ@�4���N==;�<��<b�,=�^�B=��&����;��c�F�/�x� =eR�<��<b�l�Q� =q�ἡZ�9E��cM��Eܐ���N�y&=�޾<F�=�S��$_�[uG:(�=*! =��=�rx�ٛg��z|��̗<}d�;��L=���<3쎼�7<��V��%=��uQ�Uŭ�L\T=�	�<�փ��W�"���i�!= �����$=�������՝μ�>�;���<  �L�;A����	=aڮ�8Yb�@���X�;Hơ;�(T��lD=-�I:}b#����=<�=ud=�<��!���F����{[=��6��z�<�-<*���s�<\��=��8�)G2=�>�5`m��${���;R=kk;So���H���<��W=Ξ+<�
f�[��<�sV�	q�<sCĻ�J=Ԍ'=z�!���/�B=�y��/�ؠ<�v-=���<�@=��9����<e���X<=���<$�ü���<ar=ȏ�<N�C��l�<L߹<T&=�\<�t���V=��6<w�<2�[=V�o��Û��a<qX�[�d=��=�I�<k�V�d�H=G~�;�򻭈�.�
<l��<@�n�L���=y���i�:d�9=���漺�8<���<���;Ktؼ|�r=�pJ�t9�<�N<��)=t2����<%Ƣ<X�z<%`��Omz=�N������޼�Q.=�I�<�ü5�?=���5\*=���<Ku+�!"���U<���u<:��:.��<���;Ҽ�<2�d���M���⼫�?���8�U�9#�	=��5=�Q�:��żl�j�A�V�>�ͼ)�P;�f¼�fo�1j�����;�G_=��=�����ʻ�]<=�N=�<B{?=U�޼M:=ݧ���y�<P�I<�Q<�#�LK!=�Tl;�n�<��=��C�\s�j�<L�W=3p����<��-����<�>�<�8&<����9\������!<�(�;&়���<%ai����������;?W&=H�=<"4�<����um����=�=�K�<�=<1����P=TC=Z�<�;�-X=0 �>Y=�" ��k��d�<�g�vټ�"Ǽ,0 =�ZD�:�˼S�/<7pX��I����0=�j�<#P=��*=�3=g���M)�I�=��<Q���4��u���?�5��<B�S��e=WዼD��Ex��@=��;L�&=�	(��u�<����"/;�1�=L!�����;T�ߺm
.��T>=6���#�W=R=C�o;���;K��5ɪ<��r���.=����Qͻ��H<����[��V=l���Y�< Z�$�:�qo�<u���(�;����x=Put�ַ<b<��)�	��;@�R���=�h%����~�T�e�-���"�<ȻN<c��Cj�<�^=�뫼���<�zü 9��\=v=I=)���&]=)������<�Le=~���!=F_��^���E=��ü��h�}+,<O1<�m�6ޑ��5�<C��<j�I<[�'�'`�	s=[33�)Wa�>�+=��<x����G���==G������<��-=۬b=ˉ���ĝ<	Y�<c��<bE�����:�;f=,���ټY��5`=C(=	�p=`t�/�p<1�,��1��/1�<�=:�j=�>ۼ�.C�D� = ��类�q���d��i�<�<�J�;�N<�ȼ �ü���k����A=�0�<Rh���%Q=�;��]�<��ϻ��<�:=K"�<p��<�{��с����7`W�Y<5�⻗��<��6=��h=�_���s=Qqż���;��<���CK��kd=fbp��ꓻKq�<��9��l��¥�<Ô:�l'Ƽg���QI�3�}���7=�-= o�<�Y��bY�; ޼�)_���@<�'�j�4��и;���o�0����;��6=@s�:�a?=�=s�w�����_��<`����<�
�<�/���FF<5����o�jO��W�:=�E��8��мV��{)ӻ# x�gi5�}��<R�=�q;�a�H�_��#�&5��@4���ͼ@��<���$ul��"=�f[=� �:�_�a�R����<8�H<h�=�1���f=���0�=�: �<��=c�A=�湝׽<&��Ǎ$=���<[����ڼ���4�;#�ɻ��)<j�+=��%���<`�k���=�<#t^<���<����V=ji�<5XѼk�ۼ��0���"�(p/����l��<�ė�馇���<r���G�>��m�rƭ<I]H=�U;l3e<i�=�_�;5Sy=J�<��U<a{<��; F="�F������r�<{�����;��=��d��O�$5�t�D��zJ��/�[:C=��5<�i��n ;�g��<�uA��8:��^��k3�҃��Z�;�n=��<1KE<ՁG=�SE=	2��%�dXѼ�9l���U=}L;=c�e��+���(��CP����;���<�]<Mڼ�5F��&<��+��:�<w=�-I=�-=W׼M��<4�<'�;�ܗ�<�m���[=��=>�d=�l6=�9=~[x<���<ڶ� �&�������e=�<Ǽ�o2:�~T=G�Ѻ�Ѽ=�*<��E=���<۲=�A$=:�=pU�#�=<+�{�1=u<��d��^s����<�;���q��pK<�bx��o���~D��=���=/�-�Jr<nG��;�J�H���=��^��ڼ�B5���==?�b����]";�Xh��Y���N=SK �O3����^��|J��~��@���,�<i
\�K�n< �<�S'���;=���\�;<2ڤ���=ESh=�؁<��=:͑�9��<��]=�p�<t����<V=K>q=�s\=*�?�,�2=�"Ƽ_��;7td=r"*=�Kȼ6�=��ȻZȺ����<х�<eH�<YDB<p_�<�xP�Lm<�����=�k�'%;�0.�x�Z�5k*=�Z=��%�-֥�)2=��2�;��ϼy�7=cL���|�r��<�GM=Ui�<G����x��_^��Ck��骼�V��5a<�������H�3�0�\=��'=��<�4=I~̻��j�	=�6�;�=6���L�<��<����I�8������Oẇc	�3��<L_/=m(�MC�=�p�<GC �Ja=���<��Ƽ��
<�Y0�N�ҼѣS���z�&N�;ߨ���Ѽ;��<�$e���9=���<��"��Q����
v뻸�e<6��=\}=i~b���ڻQ�]��L�<α��*�<1L��aG< �X=��Q�a�<�����b]��U�<�
�<�O9=`��<ph��p
T;x�#=Ң��~m���v�+�����H��C�HEL�0}6;u�m=c�O�� =9%���=��<�P���$o�V�v�gz���Y=N.�<��(�?z���B=z6�;a�3�~�\����_�=]�.��\=�a=K�<*Y�pY����M�T�`���N�2�ʼ�b�<M7�<sch<2%�9�Fռ�����0?��|=������"�=�;qa�/s̼>��9X�<qfv�ۣ|<��(�h=�2=�x�<��,;ZY��|1V=��-<"5T��=���<]:U<�L��UQ�)tn<�ӭ;��Z=�KJ=�<��w2�T�&����<l�u�i�����<���::��<���<�i#=p��q�缮=��
꼷�"���;D���������T���u==�v6=@��<m�)<wP�<W�S=�$��E=��;�ы��0��If�h7�=��<��-��Y1��&@��z<�S=)0�<��(��>z=��_�g����K�Y��<��d<1s�<,���p��� �嚜<R<sH�]M�:��<:<�C��<�xq�W�=�pL��x�<�-�<��	=0�N�p=�*���Z5=�r=��<ݲL<fQ=}�	=i1^<P%	;�Ղ�����[ƃ����<yk:��u3���	=ҫ��V�~�2Fr=���;��!�#�G=�=��J=��<�a=��=��kN��#�n&�<EA=B���TN=��`;L�j=W	Ǽ��<Ei����=!:��+=ťļ��	�N�L<Um߻���@���h��JvF���E��Y=��5��z�T0=ƺf0=X�;��`�������Ɨ���wv�|TN�>v=0�:��u�����<���4�;�w&=�酻��;�JY=��K<����� =�7�<�x{��:]<0Ǒ;��ϼ���)	޻��)=�-���x�;��q=.YN<��Q�f1J=/R=������=+��<Y���=M�%
=3�3=Kb�<�/�����0u=��漺�u<�l��F�:�x�<ES���9�nR]={���C<��"=�_1=�m�uJ��P+<���<����F�E4��Q�ļsG�9^�h�\W�<�Mc��=�P��4�<w�d=洣<�ߙ<W@��(�<H���0=h�3�:�;��\=e�=*f�~`=���<��$=���P<��<=�(=��$�����k<=BF�]�?=װ=�`N�<���<��<h�<Os=����;��d<�W���i�����5���U=�;�<SX��z�����c��cd6�������ҀO����<��7=�@�Oe��m�9�[��G�]�=5'����=�x�<	><�J�����<�?<�!=��!=��9��S-=�#_�.����;�웼���BӼԱ`=W��<��n��<=��Լ��J���)��ʑ;�>=a[�<�\���kz<E!n=}�;b���;���e�d?f���1���=�lI��O3��N=���j,���<`(`=J�E=a<��&���==x�k=M* �@��S[==�5��L<;���M`�<;\Q�~Im�	��<�����o񼺯=F����)�?�7���м|( =�$�<�����N�Y]4=��<U� =j%
���d=��Z�!�g����}����j�Zu=�\~�Pi�"�<񕽼?1;.ե<�GJ="�k�Iqr=FF=ѭR��ռׇ�;e\	�S{�< ��<� <��1=%�;�����ټ�Tm�&X���D��<L=��=�\"<�����`v�R�'=��w�j�<�`W=�0<*�5���R�.�hRL<��I=�Á�iw�:\(���a�L{ؼ�pu;I��<+�:I��&=@��<�ط<2��O�ٻ]��%�J=���<��� ǅ=�=� w��RR</G��#?z�Ls��u��<L�͜���<����T0�֋x=8P�<ɼX�4�#w��ayO<J�":�� ���O������T����<!�
<�0$9��]<����d�N�=�������E�C�9V$<�1V<8l-�����~�����pN�8�<8y�����S)�;��W���Z;���<�����&+=/�V��X
��V��t\�<(%Q�c����	����t=u`���&���>��/�<]�\=�f��9,���R<���<� ���pq���<z]�;�v{<BI;��'�]��s<� =1RN=oU9=�`V�v�?���#������;cd;��A�0 ̼R�� V�<���;L\=&�2=�U%���7=��<!wM��N�<O>U�
�¼��<4#ȼ�)�<Dm�9/�k�zu�;��:��c=5|=`m�<AL"<���<�+/=��E�o��<�����r/�	��<��b��+4�O��ϧ+=�R<�����<�v�<��;�$ <��(=tx:�,b<��\k9=���2k	��.�?�<�T��=٘4<(ǘ�+�_=����,-T=�g!��[��<�`��Y�&=�<�=���=eL_�Tc�<4�� �;��ӼD�v=���<=��<������O�.�
�*�=~xB<�=�<^uk���2<�X=���<Pv�ʘ=_�=������D=�rm�\��;�<X<ؾB�����H�;���<����5/�������7��m=1�<�l=L=�*��<�L=�#S�Y�J=9�=�V>=蜻2>���=F<�29�Y�c<kG=�"��Ќ=�G�<3��<��&�X)]�J�*87�!���Z��Cm=Q=��R=�%=�&X=��%9m�=K=������<<�/�;�@@<��=ݼ�����缟_=��ȼ��g���A<,�s��r�<�0}=I�M<�@<oS(��8��O��;+���,׼�o����<8�8�46V=W�L=����8���ȟ=@�����<|�=^P%<�]=��=q9<��H=�S�" �<3����[]=:N=��;�W��[c��oM�O_$=�B�3Ec�M؎��@;����<����8��;jsۻX����<M�c#H��ґ<��iu4:I�4�	�<��;Q�-������qq=�tѼ�=�1+=�Lڼ�j?�TP*���9}�=���຺�/��<� �=]������+�ե����G=�k�;�º<�=�<_�?=�q��I�<��I&<�,=�?o��!<��Ӽ��<
�a={�)=�@S��QѼϹ��5#<x�l����<������C=�廎,N�K��<d�u<����`�<�=4=��$=���;�X�=��W�#�z���^G�Uj,�F��<Ne=�,.��*�<|�=:��<3���æ��[�����t=���M����1=��7<�W��[R=�ST���]���[��j�<7a��
=a*&<���	�=��&=T��<uc�=ɑ=D`g<��i���� �3�;�<�U6��	�<�hg="�<� |=D&���+�:N�0=2B;P�<�e='-U=3��!���!�<��=�$5=j�Q��i=x�e=��:�Bx�$}�<���<��:<�h<�=�0<�(��B=<�c�C�����R=B�=�p[�Q�5�V�鼏F�<11=� ==��`�k�W=�ј<7@�mE�;m��<�7&=u�<v�(��{�<�i�X�Y<F�<�l�<L=S�g=.�;��c<X��<�>B�.�C�<B=�L�<�ۡ�K�B���V��`�<���<��攩�y�<�'�:(��;��=wƓ�k��;�uP=�|��v������/����=2Y.<
;.�s񼳤�9IC=G�g���u(�gAD�xj��v��Ǩo�p|d=��@=�1,�6ѻ6=?��i{�U3������z�q�͢��=ᣛ=!q,�O��\PJ=��ؼks����=��+<p2G<�m*�����(@�r�z=�CA<��:��<���)�=�8;�����,����_=�򋽃�=1��<��+��)=��(��b,���:�
�<$|5��;7=�(=�z<��!=�'Y�K������<|wE=�]�Q&	=w�����6�,�X��=� Z����w_A�E|;�p@=u�@�J�ü��8�^&��.���ȼ�^�<R�/=n�޻F��<���<��<D�	<3 p=�=3�ڴ���l<��7=��;�,!�#ƻ�a*�Ȅ�<����}$��+=�\=�x�;�M�;9�<zx<������I{\=�<�K�;p�;���;�7e<��'=tㆽ!8=���];��;U��DI=�r�<Gf�<�1�<ܸ*=��v<�a�DB=�=@%�<T�fj<��=�yc��2o<'�4<ap��6��;�m=|e�<�g!��N=�L{;\��<3|��v;���)#=Hi�<��E=`�_=[�A��X��!�ݫ��O��V�U�M��|	ʻ�=��1=�=ku���ļ��܄���|=�bW;S��=�:h<��<-��<�� �(�s��V�<"Ǽ�!���e��׼f�ۼ�g=��;�<��<�f�<a��<��c=��	=�R�<8�<��0����@֝�~0={tY���Q=a�B�%��;����X=:=�c�`$�IT뼕+�*q;x9C�_;;m��x�f;��w��<y��<�+o=�,"���L�GE���ù��N� =T(Ӽ!�d��ׂ;[�:=��m���Z���k��5u��%�%a,�� f�T��wOf�H6&��2S=/�=�������F=PnW=�6=r����J����ռ�W�4&#����]d�0Rt=<�������;��1<؋?��_D=PA�;� �<�5=i��<�Y仨pN;v�O�fTG=��U�k�X�|9K�- ��ZZ=�m.=Z�&��+��;�0K���+����<	��"Ԓ;�x�TZ
����/�<��D=;B���A���Q�����L���J���4� �W�ۼ��7�`8�<�tǼ���<���:�<=�==��=��q=�K<��8=u�[���9=���<�0�<��<��U���R�|�=<�.�<�{�<�����N�#�y�d_=��>=!;�;�jQ=܇�;Lإ<���<D!l�g�����@�����þ��T8=�o
�ϼ���2���h�u�`�P<�W&���9;�a�{��'�=,�ֻH�#��8�����;��9��U;\�A=����=:�U�5��<���)K�#�q<Q�<m�@=�I<;��J9㼟�/�15:=U!U;�[>�al����)=�P��e�9c.�?�˰8=�I�<���:d��1=�cE��wN�]$:��^�rBѻ�b}=����$�`=�
���qM�+�=��z<�<9=�R�(ʆ�T��9�9��tҺ��_r=�Ǵ<v=��=:�<c�f<hm��7(=�Z��8�;��;>��<��<+b=�4�;����ۼv=�O��6E==
�h<B���K�.��e��y<S��<�Ƽ�=n�����"@���<=֡=��� �4�=��;X�r=}ǡ�X"Q���.=�K�=`m�?�v���J�SrƼ8T�~�;&����;G�5��C%=�;��}ϼ�GC���ļ�/Z�%XO���<
�����=��=���r����5�T<6�\<Y�a�e+;=��]L�R��^=�A��B�:�f�<IGQ=G-����<�M� ΄�:�u�@�=8�*��-�c�>���ͼș=?���|j<���Pv��l)=EtJ����<�ӣ<8猼HE,�X�pjG=�y<p;�u�4ZP<��<z� ���=��\�%�<㑺t �;�`��9y��a��X&=Wy�y�$=�H�-��<�7S��&<��j<G��<�N�=q��� =��r='�<���6<4Ҋ<*�#;��H��*��KN=�a��<:LQ<��M?�Z�T<���YS��=�uH=�8d=s�;ǒ<�x/=yp��<<�P��La��h"��mL�W==��~<�=����X����;c�ür6����w�������e=���<`y`=cfG��6�:,Ҹ���μ�q
=����<�B<�F1<jw%�lʉ�s���Ӟ�����<k�-=��Y=�鼛�=T9W��3�<����7򨼊5��\F='�<��<��1=�,=�=�m�|F%=��<8����Z��|�弘�Z<��=G��P�]<����@=o:=l��xz</ �Z��f�'=�k;k�/�f�Q�s�E=���<� ��=�y#;=, �
=5��<��,<���:��x�jK�n�.�m�1��� ��<g���m˕��{���i�8ĸ<�&#��n�<��=�H=c�<SB=ש�;�mk={���~V��:o�_('�܀=t�/<��K��0�<q�g�?=��w��N;=��Ƽ���=��)���i=35t;�(��(p=|���oc�<bF�<��M=��=�r�<!��<�j�<z��<�	=BP�<�A���E<�$����<�=�-%���<��A��;[����'���v=�E^=(���%˺[�+����<^CO<�><]s����<���LF=Ԏ4��$�i�<�t3�/��;��>=T�J�Xl���	�I�-�v�1<����J=)3�<�E�<��Z=��<M�=��G�5/��G�R��9<���<� ����<�����/T������ ��`%=;�_�;��<ݾ��Q��!��w!=��m5��$�.��r<�c�<Gϟ<�Mt:�����&=�.�<�y=��5�&�v<~'�<��V�e�;��M<����	_=�m.�M:���e��咻��k��95=7�"=�+�{���+-=�ό�wG^=��r��y��@=0��<O�S�qͼ<7�D���輨����\=N��<�c�;`�ü.Ї����<|&S��
��;vd!<�$��!T=��`=�i�A�<wч�M�;�߫�1�=I_:�@ܿ<��<9���/t)=}��<H|)=��_=ȅ�;��<wt��lJP�.n��i.=Qc鼺=sO�<IlX���D�b*���n9N�T�#����E�i��][=�s6�g"��8;�4� =�q.<ߢ�;�<�ZA=������<�"�<��3<�MU=�3�<yQ�<��b���<��<�3�;V�<o���7�</n�u���d?=*��<U���z���2�<�N-<��^<��<���<�򗻴r.=ꨘ��d��y2x9�@=v@:=�S�*r\=��N�j!=��Y��(F�J:<�\������,��=(=Vz��K�vv�[/��D߼�ح;;*z��'3��S�<k*.��KH��6=� �;�s�h�O<�<�j��9<GN��UM=�T=3�(��=�?i��V�<�Z����A�'ټ<.�=D�;�[0�c8/�9�b=38�<,+=������s<�)�.��<�a��o�O�';�|�a>&=R�q���m�<����0=i�N�<��<���<{�r�/�Rb�<TR>���8��{��:�]=!��<��$�N=Y<*�&�o�!��<ݼT��<�%���@J3�;��<��=fb��1k�Ƕ����<�����6�=�G<�o��P�����G=��2<@��W�B�7���#;�.�<�D��V��<*� �������)=����N=���5.ü:�U�Y�Ǽ��[<�$�{��TN9���;��=�=�0Ļ���#�L �<C;<M��<L0;�*�<�7W=�vd���@��ٌ<�V=++ży���V-�T==�!�<Rϱ�+<�2�:k:��J��,�<���s+�q(.�|š<a�Q=!�7=NŲ<�i = �<�<�ۂ<��>�]����<�ie=ο0��u�n�I<(�Z����;g=�= ��<p��< B�<b뒼��!��牽��Y��Le�,��;��6��C��ph���\�D�{=�^3=�f=KM%<���<\�P�9��y;��C=��S�"�
=f;���砼R=�/�==�X=􎼁�=6�B�HP��W�<W���<��/��7=<`���H8x<��w=����a�I,�<��h=�Z�;$ؼ� 6�I�=���x��<���<�vH��8<�#�b�t&�-�޼��:=�';<~Z�:��ջe��<8�v=:�;� =�I`�tW=�u��sA�]Ǎ<!A?���|������.�<{;��a>Ǽ��:�F��^Y=��j6#=;RH���3<���=+�Ż�'��Iݼ�,�<�׺:g�=��<Q�Eq[��<��MF=��y��f���׼	�=w�=a2�<;м_��<S�X���3�>o�63=+uF<dS= ��<Y�<��f<�����C<.���<"O�־��'=˨O�ǒ";JLl�8x.=�(e��n�ȫ0=�F��P�>xg<9~��ۼ	���.=�����Wv<�Y=���<�,:�W\=�>��ļ�v�<��ʼB�#=����mp�YP�<�=F=th�����RP9<JR�;8�\��Q;@=��2��gW=�����J�?5=�r���<y=���<��L=�ջ*�H<J@��湼�y�~Y��?��<�
K�"�	=�Q��������9nH7=�>=�?μ3O�=����D<X�<��r��C=����
=����`�}E<�˞�ܥu:�4#�����@�<�L��J�;�1�;f<��3c�����A!�:I�6�ʻ`7<�g��
�<5j�<��4=�=��	=K2����,���w<��==��T=��=�W=��0=�������ݼ5�s��T(�7�ݼ	^=h�<��:�B���<���<zQ�<v�=_�<#CG���
;�叺c{�3�E�M.�<U�=6��=�u]<�%�B�=B0�=��R=(�*=�g�;R���y*<���bY��؅<��1=��N��9�<{�޺r��<AX<���;f8={yd�V�^�����A�)y]<eJ�<Kȼb�ܼն�x2<��"=�F0<�-��z~=f<���<�4;J./�v��<�*���Y=׀@<$eG=.��:	��<3��;��<�⹻�y?<vX�<�O�<41������A=]F�(f�<d�b<�{<�څ=wg=TG�ߊ���溼Tg<#]�����2��<����h=��=���ⴻr�=��l�����<;��<~A�=�GU=�?~�}C�	���45���*=��D����<��!=�w���6=�ݩ��"�(�	=7��<9�=�_��}l=�	J�.��=s2 ��C��D;�xc���=�����gQ������j< *�<��=�܀�MK�M<=�l=���<"�:�����c�L�]=�%>=�Ug���w=r�b����;_��<��E=��X��@Ӽ[ӻ�"]=��<(�Q<V=�<��ռp4o�r��<��=�������I[�<�Mp����<�:˼���<X��;=Z&=�.���黅)�<:���\4�1�=Q;<Hx��?�+�P�#�='Dl<�����4<|i�<�NH��1Bm=��� �C��h;D�[�8b<�*<�E#=<�0=��<�lO�3�i<�b��2%J<��߂����=�	���; ���<��<�xE<�z�$F������o޺-Jc=\_5<��#�������ތ;�8u�Nul=\:�<I���I=	�ü̧�<W	=u������J=\<��'�.�$��?}��"=�(��
���i<@�*���^�<��=�M=�#q�<��<�]=C$��eW�h�Y=ӣ��Ҁ�K$;\�:�%�*�YR<]�b�7߃; ;:=��N<٨R�}�����<�A���ǜ�#�^�����9ռ,s�<���;�+w�t��<(�C�0D�=�G=]w�<[T0�)�/����<u�v==�d<;Gl=�P������Gh�NMF�'�-=P�����<�HR�Q�J��;���	 =k�ۼ+�=�<�<�N<e�J<��1���<�����<^!'<e5�<�Oe��7^�B�u�M��=<_�ȼr���l�<�.��oռ����k3=�,.<>��J�<�<I�X�<W�<��X�i+=�4��[�=M�O��
A���q���s=]�G=���sק:7ڼ��L=����Cx<���;ö�<U=����Ů��勮�Ԗ���E�1}�<�S��g1�;gg<-���0Z�1�M��<>`,��\Q=��0�0Ƽm|%���<����*='�(<O�#���<'R���$����/�]j<���d�X >=X� <�m=��R��=X������["p=�}�<��=a4��#?=�'[�u�;��L9���F=]�5���Y=��6;�Y�<6(�c���5=Ry�<��V=��;��-<�D��C=^�<��>=�C<����F ��6=9�=�P=I�T<��M=�;�����<\�.=4�����=EY>����<�G8�Ə�;4 =n��<Fa�<�g�+")�E.8;��=�D��H;4��<���<�| �~Ӥ��J�<�>�;�"K�e��:��8����"�=�W=
�0=�P�v�:�1���
=1g�<�t��ڵ��K��:ʥ[��<r��ȵ< �
��l���c�add��8H=<�; �Ȃ�;�~�s�<.��ϣ==]�M�?��<4!=�p�*���0��<?^��z<���B��;l��+����W<�������<���q�J��:;�s�H
����<��J��7=5�<=��e�?$/=I����S�ێP=��&=���AbB�T���5#�;��-=��^�!=���<�mY�۸6�q�����!��c=t��i=�m�
KM��3���l��V�8�<�"H��0��s:�<z�\��+ڼ��y=2g]��Al�{;r���5=�SD���<(�=�,�=Q�����i�E��<q&�!|���K����<�A�;\#D=Q-I��XS�|�B=�}9�ʀ�<Q�p�0S��&8��u�A��L{�� �W=�_t��=ü��I=-������<&����Q�.���ļ��=%��.%��m�<�3�<�W��M��c3=u�=��|�`м2h�<F�󼎞�<u�R=�tA���;���ne��j�dS��f»xB�7c(=��:�����d�=ԙ&�P閼�>�</��<[.�'n=5�Լ��:�KR=w�w��E�ۋ$���=�֕=���;)y�j<���<Yr��8�;�'�k��<G�����<P:�<��<������K�:������1:�o�<�{^���5��L���5=��G=yoǻ(EG<�B�<xA�;ia�R!]=꼢����w^�;k�F=%�<��	��4�6f�<e�f=�T��7����5�l=�I�W�=�iѼ_�5=0,=��=�B=8>=i�<�l�=@�<��4=^�<��&���A<s�n�8�?=߸~;��@=��&��R=�wH<��)=}D��e�����栻Ɉ �%�)����||=j�,<-�<��<W�<o�*=�=O�/=��~<n؝;�|�:^&=x��������̢P<
*
��yB=!��n�O�<�wM<K�\=�eO���b�5��=�--���<8��=����R+�ؔ�<5��s|�;�ʤ<�0�<�>`���E=��z=�q�� a(=;���b�t[�����$�D�.r߼����=��=G��<��=���ϯ��D�����=� ������=��	�8=3�^=�fp��+7�ty=��x<�ͥ�Բ-=O�*=!�N=�{�<_{�<�Z�<T�f=^�p<dK= �����<�b=Z�7�o��=�;����<�-Q=��|<s�H=Zb�;��m=gS=�96;����f=�2k��A;=� ��N�=n��������ּ<4y3=��`�&:<�5�%�5��f,���=���,,W�u�=䅒�JNI�Z�#;� G�q����K�m4��C=݅�	Re<-p�<m7�<\��=��,�O�,<=�;=N�;f~5=\�<Et=x��!�<��1=q�=JO3��p�<֣&=}�=`���Y��<�G�X�p=�B(<�#�< ���<���E�M<�?��<<�R�<��A�I��;`{=��9-f<L+==����c�(�*iC��:v���
=�<��=u��<^�伒ƼAZ=SƓ�� �<=����<5XżbKU=�C��p]�6��k�nd�;^&�VZ�����?ļL9=���;��&��@W�C��<7q�=�����O�^kV<�Z�:P���`��|��<�%�<�"�]�:���<q��G<^����j\=9�=K�<"W��-�5(8=�����vgJ=m����3=��4�O��;�I4=,�����T���#�A��
(���R�{xn�L���U�����?=KD�/�r��` =ҭ�<����jv<aXD=\�<vʼ�;��<̿�<�˼��3=��5=|�k<U��=�=۳F�n#ƻq�E���'=R��<Q#��@3�(<�.(=�x��
D=:�1=cN=��*�溫��-=��7���ϻ�̼^�[=�1u�u���
�fkB=A~�s�P=3=���<4�
=Y�=<��;�@<ɤL��� ��.8�<!�[��Y=ȝ=��#=��=�-�<��6�G��V}<F%9���3<�Dj�+[ջ��@�x�;��ʼ����<O�<X���t����H�[ �<Z�"=|�&=���k/&=�9�ғa�S�<���;��~@< �Ļ��t<�m�<���^W<QM��ݾ��ӻ����5Y��^Ƽ�0����;b,=�<Q<��<>
<m}��ghQ�V{����\:@<e<��I��˼��;�= )���.�jq<��_���d=gd)���=,�F�;-�<�.��r&=]�C��6�L �p#�]>=�9&�s��<]�}�&^=�.%<��7��o���
o��c%=8@M<�������]�Ǽ�9=��Ļ'�ļ�#<tk�������<ϗ:�D=�d�<���I�:=��X=�[���0�~��������e<e��v� =s\�:�^��^%ǼAP=��0��l��L�;w�=	��������<Qp�<C�߼i=��_�]�p��	=��<o�&�OU"<
Ǽ��)��ws��$R;G9�<�#���8=�� ;�i'����<r�Y<�O��;=^ʼ?�5����;��9����� <k��&���Ւ��5Ί=8�=D��'m=�$<W�;~q�<�����<,μ��� �f��rY��@��Hټb!�<,�=��e<�0===��<S�:;��������I��9J�r��v�<W�<f:���`�ͺ��<�9���}U=L���^�T�������^����89�W<��Q�;ި0=a��ǁ����<�ຼ�S=��<��$��U�="|��Z�=	ED�� =�&<n_�:�d�<Pd���7
=A$��ǻ+\A�����-=B^W�!Z�<�؜��N������Xw��M}�$]�p�<_�r=u�=K�V�L)k���<�tA=�a���<=ʫ��[�z'�<�̄<u��<E�4=<��ظ�9:�V=W�=�ٓ�i�)=�=���<$������^W�;p=�
��a�i=��ռ����MҼ�=��<N��⼕��L<����>u=5��Ό�<*��<vN?��:�l[f�2�I<��=t��;1:<��<�jd="�E<Q=LX=�!T=�=�L�>򧻟T�<�ɫ�C5?�?b��iZ���/�<ܪ˼+[=|��<	�H=U����SR/=�u<��P��'���"�Bʼ3�[<"�H�n,�)5�<W��<�5��&k=:ި<��=��;��&<v�ػp鼼�U�;�tM�f=�Զ���av)=��!=1|��<�q˼P��Wu�<��<��L����=Q�=t�U=V=-�S��2p��}=�U�\�2��~ܼ��<�3=�<��z���C�=�v#<Gۻ�2o��``�9�<�W^=��4=Q�Ҽ�3����\�/<Tj�����%�"�=������5 ��Tc=�O�sĜ<�+��gn<�#����<wO�<'�y���=rN�=:�<�Ó<�1[�1�#����V<g����������=� �Ԉx���V���=�W�Y���,= 3¼.1==�P=�=�C�<��~�<��l6 ��>f����<��'V<J�`���%�͠H�`�<^��e��ݱ�<�Z:���1�<M�C=BV��̯=mnR�͠<5H5�y�n��]=x㤼�9�Å?��Ի�����jd��ߑ<�va�X�Ǥ�'0�<�ђ��`��׃:���<�A=�X��p ��5f�<Y��Ln��̏n�
*;�?�=H�Ƽ9��<�,���J�aY���;�O=�㼝����H���<δ�<�wͻ**�;�zQ�e"����|Ύ��z��7C�u�Q�]S��Y�Y=��:x�B�Z
5��x[=>��)%=s����:�!�=�����'<��5=���<��<#��<A�p��{̼r��{�f;w�<�|Ǽ}U=K �<M��<�t4=�"�<�V�
o�z9&��W������v�?Լ�0a�~8�O��th�c�����<%���v3�����r�"����=�qL/<0�μG6��"�<�e=f4�U-D�n�=�	�f�<
�k=��=�,�:���<��I=Sa0�!Š;~D�<c5<=悮���=��6�[��:fw��2M��e��}������;�
t�<U�F�;��u<�π<��g�s<�r���L�ȇ�;��<
D=�`s�s=�f��Vw�8K��Ϻx;
I�=|�<MS=W/-�u�Y�j�]��B�<�?=��m=�~���L<��>�V��<�]Ҽj`�γ^=���C�=����T�<ӧ��Xh#=݌�;V=�9j= �<�"�_ :=�#H=����J�:O�%=��-=�#d<	�����%=Z}9X@��#�Quټe�U=��Ѽ'���`��Y�L=f�=C9�����@8=�p$=f��<گ����<�w�<���<�չ<_�0�mL=��B=A�<���<&
����:���<��H=�m�\�3�2�I���������`�[=�(�˵�y-��h��u��ߡ=�Y7=ӻ �y9<��Uz=$�H=A��<	[F<'Q�b={-=��h��<7�;"��<A� =ƒ�:PM�;�wB=�'3=#�6���<%��:k�$=`�Լz��<r&B��A<-\:¦�<u����-=�/���ټm����<��`:�Е<Xs=WnƻKd=�=�c3=ِE=�\��Z(=��� ��<�qv���r=��i=V��<��<�aT=5d�<R��<r�<H�<2=�<���;�BW=�����=-|<�>�<?�=2�=�H���ǝ��s=�I���S�=I�����q�O5?=���;�'�����e@=����Y7�c�=���$�R~}�!T.�����7=?d�<��e<��;�[��<��t���1�]��< w=����Y<�E�����!�����=�أ:[���o���QB=�<]  ��|=�G?��B����>I+=�_�kF�Y�o=�BU�76ͻ� t;/�<V��<�p�="/ü"��<3�_=l"Ӽ�/���5���<QK<�ۃ�<��#=�<�; ����='�#=X���,�=}g��X=���~��f!=M�=�2��F��k�;�����<]+
=���<h	=ɼ�5=W�p�($<xqI=bo�<D�+��U��W=��`�+�ݼa�/�,=��@=]�<c%<�4d���q�����A�O�����躏��<�[a=��K��ԻZ]�<a�g���z<�������<�O$;7^O�����P.=�r���f�<�l�:,E=��W<A=3g��5k.<��;�;�;5�8^���"p=X���&=cr	=��<ʡ�kRl��FG�i.�D���u�&�~��M��q]W={]=V�R<��=C0�B��pt�5�F=��@=*���0%��[=gf��q�<k�y<�=�	x<��sռ~�n�KS�=��4��@c=�DV=#��;=S ��6=��pƟ��=5�@<��<�:���|<V�S���հ���9=���us<� �=����C9�GJO�i���m�<��;8�z�[�?��s=��#b;���<��<t-G=ڵ�<����>��"2&�Y�N�fC8����< ��:��T=ϞG���<����i��M6='�<w�<
��c<�� =b�<�+���폼л?�:��3=�&<=��;��`=%hb=�Q=�z�~;��r�;%z�<���<[�<��-=��H�<mO��1=V�B��k�<[�>=g	=<x�<����tAV����ٜ�<�.�Ox���%=���$=�K5=(�=��|����<;�;����<M�]9H��Y�K��\=�Q=�	�;F�<T��<u�9J�a=�΀��8���-R���:�&b���0=��=�	=K?��ʜ����;�̌<��=���<W���#��U8=;�Ǽ0�Ӽ�C'=�~R��d��;l2��[:���[�Y��^Uo�����'�z�8��<\Й<a��<������I=�2�-缪b=��$=�?s=��A��yG�8s�<;�i< =���=�(�<��<�H����g=|��<���R�<>M��r�ݼ#��;�6=�з���<��W=�1'�j"�w�/=[����-=�ZF�\FF=|�g=iw���̻	�$<y�=��F1�T��v�<��&=�n<�VsW=$��<reh����B�F=� }=��=�m6��8���Z��X0�:�ºc��<vU��Dq���^=�"���\8=�$�X���鐼�Ѽ�1A=��������7��#=R�����=Rxx�SC=�Z�<XN=>�S<��Z=�*���=���<^�N=����w �ݗ=`Ӭ<}�<��=�0J=�<=t�9=��B=�W���*����<��4=P,�vY3=��E�=te�?�-=YQ<S�=�7+��[���׼��ٻ�4Z���C=�y�;9��K�-}=׺�<���<aλ�y�=����S��_=�t�<�6=՛/=�l4���=�=�q�==7C<$�2=hõ�G��rG"= �<A���3�l5�=�-���<nXB=_�<�W2���6�4��S=�jB����ܛc��rW�0�c�f�Լ�Q���'�E�e=�I�<;<=ѯ�#[R�g��;#�= VR���	���s�N�߼{;v<,���7D=��ʼ9JE=(��j=�Y;H�
��Le��#=�)�<"��:1E�ê{=�vB=��.�z�<&��;6��<F��<���ގ</j1=Պ�"Mu��b��&B� �<M����<*�%�=��<�:m<0ee=�&�:Q�H<B?�G�l�~�P���ݼUT<1��;���j �T
-�>=s��;H=�̂;լ�7�\�0����|��:0P=-s�=����2ظ�m��6����6����b='iA=ޢ�;�i!��=J���K=B�<���9<�B=�;��X=]Lc<����{=y�/=$�D=�O\�MҢ��Nq<M�<���<��N=[��W
�*�7=���<�uY=��"�G4B=�����zk��sk=�=�L`;��L��^K=�����������,���ێ<צ�<fwj���6����<ba+=��<>�'<|O߻FA$=s..��u{��n�;��<{ռ�w�<bm�<��O=f�]� B��,A��-�E�<Vf�#EH�� <DݻV��<R�8��S׼��9;�O���?���|=+�#�B̅�Q��G=�������⵩<�/�;��,�.>�;��;쯳�J�u=@5w�<^��qA�c:�<���b���C�6���;��n��1/�<��J�t�=�S=}��<
�t�+���~Ɏ<oܶ<Y뼘�3��鶼�>����3�҈�1=�(�}���A�;�B�;Z�^=R!�;E��l�M=��`�j�=��f=�����$=����5�-��1�=�M/;Z`<��N���W=��\�D���=�@<��i=#/(�!W=��/���=������E=c��:�`8����cp;�^�:�D�=�jP�����Ͽ>=���W�?=�r�<�>"=�y�B���j�< \)� �i=��Q=A�������G;�e��I��<#�9��T����<T(=X�	*=��W<Z��ks �+�5�z�s<��<�I���s�	=rP:=�|�<�2��<���w=�&=��n�\�?=Im|=�N�j�\�[疼_?�<*�V�~�,�;��<��s�=P�|�=��1�/�3mN=_���A�;р���7<w9^��`��{�_<�nѺ���㙍��o�OJJ<p� =����dK�E�t<�{��c�k�9���¼m�K��뼉�+<r*�hS�����|�H�;�=��1U������q=���!3L=`k=Q
�:�b��k{��m�<����P`�=m'�d�[<Σ�W�<9� =�疻n=����(=������<���N�<��i��= �<�kQ�G����9!=;tN�]5����L��p&<��=���<��S<���C(d<��c=��<��6��i;�F盼�8��-K<6k��N2=�A����8�⯼	[�<|�H�6];����N�=-N��ǫ�%dܻ-y��֥�<K:+�;���(.<�u�;7'=��J=e�x����;�L�<Kz�;J�Y<����<n�e9���ߗ���C���x=� �<&��<�<���19��	(= [v�S��ج
=^^c=/
���U;&{�ֱY=�=���<>~B=����ົ�����=��ϼ��<;�<ּt ���t=z
�x%5��\`���V�%~==��<e�=�����}i=���]��;�+=]j=�T=�d���<�%;*�Q=#e`=dC=��P�xN����<�ļBz����Fm�<x'd=N���0~<�S]�pI<���		���<��=� ���<���/e�<���;
�� �.���<�����b0=X]�}�=�K=�8�<i�;=��x<
����0g�������n<+=��M=0�'=�9��i==���;c2�<JR��U�9�C��+D��5<���;�.~�x�<M�A���;��k�@gB�U��;�|�;q�:=��%�U�=�Y=<?C����T�[�� =���<t)��`=	 K=��c��.�<(���_=��M��(�
HP=~�==�R<.��b?<�g~�o�R�.^�P�	=u��uyU�����':}����̼�:��U�<<�9=�M=F�\�n=O�<��"��tu�u��,$<��=��Թ<$��<��s�|*�b�X���!<P[�<rz��>�WO3=��;��@�S�G�S��wʼ��kQ<�Y��T=t�M��Ɔ=;_����<��(=v�#�r2輔�P=/+��j��D�q=y��B�d<��#�Y=e�
�fa!�܇<{�)�X&�Ox9=��-<|��>�q���=1�.��'�� J=k�<�=�<�9����<�Z5=+!2�(=ػN=��<��q�?��Y�����<���< l1=ƕ)�P^������Y6.=&=j�= �,�;U0=�Y��O[�I���.��$�)l�"�<����9�S滲ه='�1=��N<���<g.��+`���<����ü�E��JM:=4Ѩ����Qp';�FZ=,� �Ǒ��J�9=8X@�9d=m�C���A��[�<��d<��F���=H������������y��5[=[t!=b�м���=o��=� p:x\k=��<��ȼ��=�G�fmB��+3<��:����<� O=���<�6#�DE
=��o<�F=m�3��s���;��P<3~��<ᖼV��<�Z$���=�1<�S�=��=Մ�<�;8�h��a��@�<�3�;�/=z6]�c�9���޻��:��ͻMO�X0��7][<&L����g<i=U�e�	ê���-=3��Z\����W<�~�<F4d=��^<�&�;�^\=�c��t�<nUY�<��:�<��0=B�2=�U'��T��<�=�=�Oe<�C4����;}u[���=����P6�S��<��F=9�ݼ@W���ټz9��C><�/�q=�90�eF�����I���4>�C��)[=���<���|�X�<kϼs�(��#'�&h�;1X<���(=� :�Wb=��D=s�w=V�)���4�c۶��O8=��@�3��;��=��L=]�Ѽ�������<�㟼QK߼��=�Q꼓첼v.�<Ɛ"�����S�μޥ =��<�8�<=e�=�:=���;!%B=�e<8,f=�-���L�I�;o�<Vj&��$��d=� ޼I�i��5=�\<�v�<H��< [�;jq���f��%߻�;8�, |�L��<Eo[=�+����W=KB=���<�83=?d=�\����<#�+=kd$;���<e��ٌ�<׽����<^T���b�<��W�sݼF ��s�;{���̑<��=��;���<Zq����j�O?7<�Vt��J'�*2�������@���=�4���ǻ�Ӽ���:g�\�oJռ�^��Uɟ<)d#=��)�4�L��!�<��7<��<VC�;'�p>�<�n�<_�
=�$=�v����P�绳C��`J=�>_�nڼ�a��W3=�^�Q��	�<�l2��<�8c=R��<��5��x��f=��!U1=�m=��c<z�<nИ;�:=�H:���<�8=��漎�k=_��;�=��(޼L���!Md�k��<��=[MH��l"=�;=#����<���0G=��=�{���$���T=~2,����<�,<S'ѼC��<��μ@�6=:l# =��o=h'�YF=�e�=�|��<�<?�b=ϩA=9S�<i,��F�8���>='�[��)�<-�ڼiE�ޫ>�[F���=����,%=�I�;��&<�)��3-�X1=�\E�/�м[���G�<E�=g�Q�<�2�.��<���~	�N�%=��a=�z�;��׻�=[�=-H�<>�<Eʂ�/�P�X�N��(�<�=��=��=�E*;A@f���@=}�����s����`��c�<�C��� �<�N=z�1<0S<E/=#�/���)��50;�#=�3=�(�<:�<<�1=JJ=�ݨ����<�\h=���;]X=��^={��<>!ŻDE�<�o�<����ֿ�o��<N�<=F���Q=���9��㼇�D=k�4=� ݼ*%�<!�H�� =Q��ƌ[=H�#=��㼷���^��9u+��"��r8k=T�v�-�<��X�7���� ��s+���/����$	=��T;�[�<�Z^=�[�;�(;�Lh�����;4μ�4G�}=ת<�(�=#�R��1�<	/ƼL�&<T�<ܪ�<{ڽ<�v<��>;�i=	�=��5�u���@��b�<QQ�;�� =��i=~��;�1�<w)L<�kJ�G{A=3I�������z=�B�v=��/!<5��	bL=���-W�<��;���J�H���G�p�ȼ۹�;��<YhջiӜ��C�Z����ܩ<<Y�%�=�I<<��$��{�;�U=��R=��<�=�v��QB���"=V���Ak��a�<���<
G=�R����;ϯ#<��<=�9=����P(����?=�=�<���<����]�<Ti���;λ=�t��O��gc<��p��&�<�Ħ: [k=$oH�BD�=�|��2]�<t��<��<u!�_�W:��U��W����<�N�h/<�y={��:�4~<-��<�DJ�~
�l��;���:h��;M��<U�s���	��<���<
7����;�� =�L��4�<P��Cַ����;�/L�ԩ��fQ<�%���l�/W��=��:=T8�)w)=NY=��@����;��L��%e;Ֆ�;�����)��/�ʭ���:4=1��;P�<k@=EՍ<L�-=� �<�gɻ@�W<��J���Z<V!��'���=����:�<f�>=#!1=��4�5z���B��^W*=2�{�hh#�u=����c�V���1=S�<J�9=k}=�҅�t�H�VH��닼�S=4��<|[?=w�<���<�vm=�o��A/M=�S�(&�;c�<�~=�^��*y�<����@�8:�����&p���n̼G�K�AK=
@=�zo=f�Լ��j<���;u_¼Q�-������(���=�
I=��=��v��13=�&�<��=�u=~'��-=��c��o�����<c�ȼö<	6!���ɼ�m=4�<�2=wWc��缗A=���;�W�<pt���[�<��=���<N�z��&d���<�P�;c塺Y#�!��;�4�<�$��琾<��=V����T=��F;�T¼�u��CC=���:�}�<6I���¼<`=7�����;��h�,(<�zM<eU<��D=	�<�c���.���k=0*=~fL=t�����<m~Z����;��==��<� <s�,�֪����<{����׻�f �)T������C�9�mVD<�'<"�C������!��;�O=�-�HR��z��ض�9=�r	<�X��%=�q!=n�˺l%v�b�:=�*8�'��<M.=���;��@��ƼV� =k�=}3�<'����0�S�<b�<ب���� �-5"=���<�6�7p?=%�<@�ʼh��%O�'�U��<��G�Xm���	,��O=<
�<_�f<���<��=�P��_��kZ�A�l�}�%�Y2�З;�"42��m��7�E�[<Y��<�n��/s����<@�D�i�Z=d�1=%�<Q�]�5E�<٬C�jJ����[[�<],=��c=r�B������<i��85>u=r�<�Ϻ]�?:��e./=� ��=�)=���;۔<��伡Kj�t�<���q�<��Y:��<�!ټ�D��=h�M�z��<teN=��<ؼ�<	n=8���2�O<�=4�<#Y�<�T7=
3���=;��<आ�����<|>�b���˚%=��>�*Mg��f1<��<F�<"� �	�x�S+�<��#���`��=�v�<4��Z d=^����/<_.�;笹�Cּ�\��W��! �<}�t=��=�T����=ɓ��(!�Hz�E�=�	ؼwϕ=���<4#=��< =��+=mO��i7=C�ڼ�N�=��;e�T���Y���<d�ּ��U��!����#�j<�|�<{�Q;�
=�?M=W��<�0f=_�m=������p<?=?�o<ؾ�<�o=Os<�^1=�M_=��=��+�f��<�<_P=��=�/�+Ef�r�ؼ����/q;�����;a^�"���ȎS��|�=��<��:���<���:��=FJ�<��=�>=�Y���h=P��<�=<D=�+_���:��Q�#7<ˬD�^Oe=?�<p*��5�l�<�(���<�D^�^��<���<6/ļ �<	��<���Des=���<���O@��[��~k=��;��#=����ªG=��C=���<j�.;[�A=�i=��=����~��V=`P=AQ5��WR=�)M=���<Ж!<�=t=:��<|�
=�l<�@s=�<�Mּ��Y=��4=`�}=��=���<�����ﳼ�k=�;�<Uv�<=ʦ<�Q*��2�V��0 ����ޒ����:���U��<�ڊ�v'�^	�<Yv�;�X�]�3������6=P�<��J��6/�F���P[<�y>�*���=4�<�rؼ��ؼ��!�;��;8l;�Q=��=A�R=BB�7b��u1!=k�K=��t��b=�%�<�&�����h@;=��3=�H|�N�S�IF�	6$�۹L���=1I�T��ꗊ<~�6=f{=R=�4��|�?=4Z�;7AɼyD=Y<�W=I�u<7�����I<�:=�< ��<��{;̭5�sx��)� =�r���=n��<�=���ἜX?=�"=���<��<��q��㼝�o<9&��I*����^h�<s���=�<ȔT�{�;9R=Av�Ί6=��e=|�0=�<J��?W<ډu< �s<��C��gռh�<�e^��1=��$��>�;�=W�=;�:60���f�Wz�<�?�<�!��t��z�E���a��5��M漤䢼��i<x�=�頼��n<�aN��>=�$= .�=]49=a���<]��7ۼ��� K�<��4=Rq=�P;@(Y��P"��n��)��XJ��
=T�@=�JX<^-=@=� m=��%����<,\��I�m��H�'�R����m
Y=��λ��O��$�<���;�UR��Jt�'�<�:����dAD���B=�����1�<�\=��x��Q=8�}=}X���eλ_x�BfڻGj==�i6=E�*=����hG�_H�<i��zҤ;�d�=�r<jrB���_�8�:����;]ؼv19�)��������(���=��4<�22=	���k�t�;=lM;B�ļ��;�G�:c��9�=�⠼��1=N	c�E��p�4�w@B<(7J=7�!���k�V��	i~�Y��!ڸ<1{=`MW<��K:i,=G�:�=�a"=R	8�*D��� =�|����7���f�s��<P�r�1�/��K�"m���=г��	���5�������<�Y]�g=W(K��M�<�X�<�LB��Y�d�:=�K�����<.��-�<}�ܺ��{=��[<�k�<}R<��:��u��W�<v�f�K�U=ڣ=����z<-=�:�H�bUX=H�U;9��<׽-=�7 �݉���?N�ǌ!=�v�&�1�B�<�Fe=�뢼���vo6=��7=�?=jq��r7����<�pr=�"_�3�P=꧆<�/��L;�Q]��/=��9���;�%�X=+����		�[��=8¼=�!=�G�<0]=�s�;��k���H��Z,�׵+�y��<z��w.�~�=�VY��+Z=1�<��!=�H<��0=���;��߼K^D�<�=Ҭ,:#ZF�ga=�@������;A��Kf;��;��L����<:r�Y������<C*=ԕ�<N�S������#GF�[إ<��w���I�0��<��t��pj<��u;�d<�"�;9�h<��J�D��<��;u�f���&�9�#
�<B�Ǽ�=! K�lqd�t�Z�'�=��<k�����$���;=�=Z��*=To�w�8v;)=}p]=O�o=�#v=#)��.�I��]K�_�;^Qﻋq�<�%E=���ߟ*=�?=Ɔ�A�a�^�6��μ���<W{y�s��<�jf=+�e�2�ͼq��KB���c=���w�-=x��7�9�����9����!=1.��x�5�Q���9��<R'z�}��+�t��bs;i�	=[7;;���<��<E��<:ͻ�dC=H�û�t=���N��s��'<t�<.-=L�`<Ƭh���,=v��<f;<8�l��n�<�]�;yT==w'�I�Ҽ�l��e#��e�8���<�넼������ּ��<t���k�<��<Hiۼ�y�;
�>< �p;��=��	�<�1w=&��<&�<f5=���=PIZ=F�<G�<%9�;4���P?��-ۋ<��<ja���#_=O�c�`�2:Wⴼ�l�;�|�<�X�;-����]�����2c���4=˘.<���<[7�����U�8=��e=�<q�f�O=�H��-�o��������<~#�<a�>�s�0��-S;S��;Q=�'-�rG`�BmD���<�u=L��;"E�v1=�;=�3h;��A�S7�<'��<��<��;���2�K�P�=�ڶ�1'�<�:Jp���r<Zi�l�<h�=U�>=��<���<oͅ�(b��](�_�ݼ�<�l����y��G�P�<�d��4W<d�<�v��������:���<H?=~��:��:7X󼬭p�|�G;��
�Ԭ.=��4�3=ɵ<	�`=}��<�kP=�h�;��M=�?<��Ѽ�f=�'=��<�F��eټ/�)��{<5��;	*�:�sr����[����μ���<d=־�<bŞ���[<�jּգa�J��<��z=��� 	=T�7�	��<�®<E<F!:=i';Dc���<,]y=�e��W���<��6�y�4����(Ȁ<�k#�)BV=)�<0Ӽ��m�u�=P��¿�6?��k#=��S�c�<��/����<~�1=]�4<�G���&��&+�]�a���F���<�Tl=HMr�����=3uB��*��I=�Df���s�|^
���=1�i��Ǵ�.�G����ӽ<��=H���ӻ<.5<�lռ1F=�<���;�N�<=m(=�:	=*��<`
�<T��<��F=�l��y=�������X����ȼ��<��U��[��b�y�X0=�;!<�uV=(g�S=��Dx=v!�D��G �:�t:!(�<-`=�o�3�N;��9��
�<\�-=?����FG=�{M=�+<�>�3�;`׊<8�N=v��<u��?P���J=�e:=v�</� �<s0\�>`�<�k��i��l �PgB=z<�V�N=��j�Y�2=�/,���?���<��=�������<���w�<�ǭ��L�<5�=��=�<'��x)��Q7��9={b�<x�d�G֒�+P�<�&*�Bec�77����&�/��<T�=�ϼ�4��\G�6;��ʻ�;��te�1���5����;�D;�kf��OмZׄ<�?=���<b�+��8P����3�)=s{3=$m�<�Q�<��<�9r�["
�5Bk��6h��g �-=�^!5���y=�Ļ�g�C���[o=&1�;ĭ�O�
��@=�G���<�����<e����}�I�;�zP�5N"<~ c=�H�C�(��==Y��;���1yk�S	����]=;��P�<��[=���=@��a_�˺V=��F=epB�ܟ6�������
r�U��<.�<�j�ռs�W�Ŗ<E�Vp�����:�o��[�<�'�<xW��+&�<=�����*����;18��o���G��,�����<`�t=Z�	���;'�1=�Ϻ��Q�A5B�C��~n���ˈ<UO=�O�o�P�'=99μ�S�^�<�S>=(�~=�=�{<J^��`��<�m4��[����;����In�9_R�#v<}F���x#�Nk;d�P=�4���(�l=��l=�Օ<�꠼-��<�o&=QD=u]*=x�=�X�<�B=�6����<�U�<�ՠ<D]�<�%�fe���<_�C;T��<���<x;g=�,K�V�<�~���t�Sma��GW���?�ܾ(=�U� ��Q=w=��[I:<vn���� �R� ;���>����==��	�Ejۼs_ ��%=F&5��� =���<Ww���
=V��M�M=�Wc�����>f<1,(=G�,��B�;ZY9��A=Jɶ<�֍��0X=�]�*�=;Q�=5��<.�<]o3�<�<�@!<j��;�����<wx�<  ��r@�S��=H͇�{Q�<V���Ԏ�⦅��ZB�}@�<��O=o������<�d�<}u���yN;�z��ZP�<�t�;���;^&��:�9=�0E=�#˼�o<��r��n��k�(��n�;͆껗Z?=&���_ރ<=.=�E=�gW=P^l=Vz����=b{V�=b�<"�f=]���hK�Vi����.�>)C=R�>�
U���@��F;Vw=Wl�k����h0=ky+=\�D<��L��u_�!~<�#�<맏<�O��p2=X����/=��;����<�#�;�Z�<�f�ۼ�c����:�<x�K����<P<;���+��Ղ�	F��M@�<�o��,M���I�(��<�8Ҽ�
�<�],��4=��u���<d<�E�U1%=��=sH�<�Ut<����ڳ<T���:=n�����*�o�B��Լ8p��wM��c)�Ϭ�;O�C;o�i���������0l���=U�E:��G���:?�c=r[=��=?�N<�ֻ!�����њ��������ټ:�U=͕��t�r=p���#=��=��;��ϼ*�,��YS�cЮ<8Y��와<H=q��!kf=l	�6��FI�x� ��B<��k���<�^�[>Q��3E�<4g=�Ҹ�H��<,�)=��@=B�H�1OK<�. ='�����R/�,Vt<N��=���9u�-��"�<��� �K�gc <�BE<Ob���5-<(}W�8�<�K�<���Ą=qT+�{3��A��#��ݟ@�78ҼW�#�Ӂ��c��X/(=�����5=��<�6>=��W=ϴȼ�<$���N=/���)�<��/<Ն%�o�׼��&=t�7�'ɮ<�\[���(��6�<����'��=�?$�<@hT�v��;�#�΋6=n��<��i=�<�<���<�W4�oiM=��%�����e�<T���{�*<�5=��V��+�J%��;� ����ʺW&)=s���;�&�Q���<�����.=�uX=$%�<�5�����  s<�=��¼z�$�������=�ȍ�|� ��Q=e^� �R={+N=�Ӑ<[M�<NE<�FF�f1 =����<���<l���<>j=�B�B���]�v<^��<�{4����;[�U=���,8��@��`�Y=��R=kY=Px�<��%;k-O=9l)��K�<Y�=]U��Q�:=�;5=��=�U�n��EY=YPS��F���:#=�^�<);=�GD�wFM=V�D=�L��q�)=H|�Gk<�i<ɤ0=�<5
=��=?��۪�<M�<���l�E�ë;�~\�<Y'�:���º���<>=���<��=q�K=�v�:��W<ܬd=��Ƽ��=J$�<�4��.h/;!.����2=�	���z=o����=���;=�=M�B����<���;P;�����<�d�<�!=�=��;=��d�޼��!��{K�Ƒ���(=�u%�ķn=��=�����&�7�>�nҟ������<)�=���X=���;����2�;��H��;M=4SO�M��<Qk�<F�=��N�R=�*:=���<�<��A��<̀U�
D�<�#�;�Bp�:��<�3=�Q=��<i�3���`=��=!�<�y>=��@<��k^=�R�<�.ѻ�p�>P]�B�<�X'<ɢ�|�B���I��֒<U��l�<d,�?�F�;���J�y�2<A��;��|<�$���lX=�0�<���m�=yv=TF�G�d�H�J=#�;��ü��߻��<8�0����ٰ��m.ټ�� �^��;�%�s-X=�mC�~��=f��<�1E� �;�}���H=d���O=&����k<A�=�"m=]�&���G�N ��ݷw=���D�ѹ���<̈́(�=�;}T�<��<�V�<_�c�"���B�C�μA@�E���#<���<��9]�<k�Q=Q��<�.g�^�C��i =+Q���̆<{�<��x=g^�k�&�&%��򝼵-"�n�<k�;�0�j^�fWQ�͊缪Ķ;T7S�D��Y��F�E=}Ƅ=N�<G�'=ʶ�娐��fV<��ƻ^��<*v���'<��a��h:<�5���l/��컥n�MW=�&�<�s/=�#^�*%;i|�<�_��(i���<��t=<m=p�ż�f=D�k����TS=��'���ü�;�;�3�<�μ0��h���>�<` ����;p��T��<*b�;�~;�c�rV�<�
.���=�<�S��H=��	��z=�ݡ<�S�<xK=R"=Dsp=w� =l/3�b�@=�V��\Qm��'=vJ!�g(�<��ܼ�7�;J��<�¨<�I��/����<=D?��<��1�K���m=��ռx�X=��K<`v�S�/<��ڼJ��;ె<u���]K<欍<Y�=����W{<
F4=�5=-Q��4 ���i�"b{�w�=j4�<����,�B!μKR���;�� �	m<<(*<��<{�v<�<��{�rݞ;�9N=w����_>=��V�_;�еJ��e���`=⻬��>����}H����.<�G_=��E�n=�ՠ��Q��kּ���<m� ���b=@=1��<<
�<�-ݼ����/m��5|��zU9= �ub�<^׺/�2/=08=6x=�\4�,e�;�)��}i��
4�s���@�=8X�&����u={�N=�&޼�I�<RMY<X�<BŊ��0�oR=��3�{��;��'<�f#��X�;;�<
�'=����=�3�#��<PQ��2�*�=_��?��j��;����|�������b�U=/m1<�X�,=#=��=3�^�Y�<9=߷F����<{tл�y�`����������<Hڅ;SB=#2�_�=�S�f<`=C�
=�9=3ʱ�G.�<��9��$V��� ;�}��t~=w�;�ր��C��v]<F�s�@����:��'6
���K=/Ѽo<R<��r�a4<�����<"�S=�r�<���d#�S�?<hN���_=�"���3���LG=r���VW=_
¼P�E;Qـ=��&<��}����8����<~<�Z=�G��w=����n_����X=՚�<3z=���{Ty=�Js����8	=T�<��g�"�p��Q��-����<�O�<�U,�9�R�<��<��щ=l�*=�t��,�<�t�:��=U�<&j�<� �<�1,��>�*e:=TÝ9^t輁�:=�E���g�<�yD�v?=��Ƽ�p�<�`�<(#�;��'=>컙K�;l�r�b<&P
<@��<Ղ>=c�+<��
��tw��ӌ<x���� ���4=�<x��e�o��A�%��_�<rgw�)�����<�D�=��<��=`S��+@=�:m=��ڻ�=O<y�
�i��;1 g��<�<�ּ��=^6�<��D�S�]<�<��;?�!�*�%�G���<`���0<K�|��1Q��H�;�P1<z�:<�� =UӞ��Q��m�<��=���<P���{ �� 꼝c��@���(=o��<R�f���|=_=���6=�`�:v��+S;l�< �Z=�`E=�{�����.E�<�t/��$E�q,*���<hخ�;��<(��;��=�7'=܁s=�Y����<��<BT=���:�>=��ܴ\����i�&<�#�H�I;j7A;��:�#=�&A=�[=CT���8=l�W=Ӭ=s�μ5�����了�A��}�<�'n�&���������%=�n&� ���~����<�û]f�eW�)�*��ּut1�~ 꼰���.�<���<ў�;�����T<>�)=�H=��^�< o�9�Q=�m>=��o!���:=}<y3��ȼO�M�ĩۼ��j�M<9`l=�2��?=<.��EK�Jc��Q�;��-=�:ü?�<_�P�
���^Z����<3F����=�P�<J8�6�Z=+��<VN3=�ֆ<�fҼK�*<bq�J��e�=#����m��Ż��^�Z�l<򈙺!�4=�VT<W�=U�;����;�w=3�>���O�����@�����A�k:����Rߪ��Ny=�>(�L�<U",��?�<�2J<����'���;��_x�<�x�@�<G�)=F<�<��"=�+=9ZG�k�08<�B5��7=b"��fp�<��;��<��=/Ki=(�;��F�"Y��碘����^������\=�'?=����'-l�"�!<�u���j�;��!���K�z2��O�;�Pn=����ż��&=pI<�8C�091�, 
�	��<� Ƽ��79��k��ă�W�<��+=�W ;�u�;l��<��]�BPZ���ϼ�׾��݇�Czu=���<6�"���<9[=�,����E����< �V�m<H���95�=��Q=W=O��t溼n@����y�iv}=iU�;��'<6A� 	���5�<h�={<eZ��BP����<��X�<9ּV��<�]`<Q�V�H�n<�����;�6��b=y���^��)�<�q��x�G��*Z�24]<"�N=�'�Z��< �����2��@!=�[�=ZZ�=����P=�?���P�<F�H����<Vǻ?ѻFGH���<�u���I�<.���nb=Ue6=I�<�	=�ɕ�`����U=O� �J�M��S4�XIV�d�:9R�K}�;O���g�t�IV=�z�;V�c��IO=#��<�K� LG=i0�<��r���,=i~F=M�=h���c��h���A�s�=�yI�gk@�><��8����zb=ا�<G�#=�5o�g��<��=�B�]�A=or�ga<�=&94=�%�<fZ�;�O�<�tI���s��=ݞ���p;��:�2�<��7�S��<�@v��H�<"�:;��
=N�[�0��v^���"=�xa:}��I����i���>�M�����U�'�b�j�,!�n���;��v�<�ü�����4�7���1�qJ���<�cs<��O�՝����g<D�O=)G=��H=��e�d<�=�\L<��<���<j�
=�pK���5=�N����</�=���<g1����!<�=	��v�;;�-��|�<�S�4�g��<��J��k=dW��|<��<(��<]�/=�J�y����
C;o=@=�!��*�;����Ҽf߯<�<�A�<a_�<��=`G��=�<���߼�P����_=��|4M�u�"�z���!=
i�<�g=�;V�#�����&���缝�F=�v0���;Ϋ�<��&=�a*=�8�%��箭<�f)��p=`F�l]5�ԣ	=�-S=�h*�#qi������F=�ڼv�:�y��~�;G�,=�bC�D4��c<{<��<�^<|Jt�ܮL=�r��6.R=�\b=��	eF�"ɿ<����eϼ�X=]IY:~�9==�]=�^=���;k����;��D4���X�4�2<P�G��s=߮�<�<�y��m_ӼL={�ֻZ�J���>���==���f.=K=�<�3=��'�mU=�yK�mR'��������� ���)e<�Yn=_�y��2(=�U��0W��B:�����8^<�#@<1�=��$=�Τ<aiʼ���<�8���N=^7�i�+<�����	����G<�0s�/�<6+P<�w��FP <k�<�E=� ��4h=#�=�ȱ�L^=�v<��=�M!=�D �q0<���<A�=��L=+����z�A�W<�t=Mm����<P'%=��I=��F=g|���5=��>=��'�N�'<���Ib=��U�s=���<�<:���g�x�r���ǰ
=b�2���?=�)�;:���L_2�����HF<25��P/�Z��<Cf=��Z<�]=�R�<{��i2=��v�m�e�A��<m��7S}����;,�(=0&2=�=8���>��;� Ի��=�2:�#�Ӽ��λ�ֻ�{M��{Z=(D@<I��,L<�t�<,l/�޽<Ѫ'=0�R�K�;=�"=(X�==��<1���>E��E��x#��6y��0$�$[�Ǐ����<6��q�c<wč<̶�;���<�K˼|��=8�C��D��7��,����<Ãm�#��<�8�|���c�kfL��u*�C���K=��ռ~=��=���<�͸���5�N��<�U?<VaƼ�<��=�l6;\Oؼ~��Z=%i�<�IO�����tš�γ�<���1#=)9�3
e=�=]�c/�Z�<��<� ���D�����ּ�哼W���r�I�.�����w���.�;:R=�D�MF�.��<��V���ּ2<����y=�k7<Ji�<G��=g�ܺ���<��<=�X=�?�<���lw�Kv<\�w��t=�ת�y��;V��$���_U=�k�<��\= 0*=�@X��=���=hwk���
=�=e~�<��E=M���B=���<�h�<xc�^h�<������<Wc�<�]��&)=��<� �<s&����:��x�z�N����,j��6=O3�;į4��=�. =q�%��[=��������3=I���-��D=U�{;�=�<,#�6��<���I{<����]=�f�P����==�5=��x<][���!�gr=f���ȗ<�&�:}U=K�w=eG�<i�I�+7ϼcJ�;q�4���;�'�=��E�@�=j�~J=�N'<���<�/�� =�%.�V�X��]��<g��m��Q=�KM=!)�n��<�=<l��<U޳;�N���Q<V���s=���<�>=�=�;]8:���u<t��<��Ż�c=��#=n-"<����%n��Eg��;��=Ҽ�=d<���;�>==r`q�P�X<�~�;��?=2[�<�"���H�</V���g8=��<2V"=Z�(��X��P��<5��8��<B�0;%u=y�<�<�o=�U<_��WV=z�R�E�=j�<!��<���<�q������<��#=�t�����i!=3x=1l�<�-���\��=%2��2;�m=�;���<�4�Ȅ�<LG,=�f]�>��<_�:kS<�-Ⱥ|[:��!=j <��O�����ށ��r:у1�`Y�%c2�������r��Px<9Qt=D�.<�<�.]=;> ���
=��<=�wۻx�+=qJ�;���;��=�<Ƽ6c�O�+�B��8�I=���<�]ڼ~�y=�-/��bs=�+'=�׻���<�&��}:���Z��ݻ�k=dVC��4���/;x�$=���*1�.%�B�K����ڼ�*W�&�O=L,=���@0=��m=��+=��<U��X1��?"�;m><]� =a�!�>�u�<<��=Q=1~�0�M�	p�<��M=Y��<��o=��<sW� GU=���<����s�[<ǵ|�Q=�?���}<B�_=�iݹTv�ǂ=ݰ�<ʸH�h�=Mù�5/W�a����v��+=�=���B�л�0��O�C��{]�<7��l�0�E8�i�f=���<�]!��u��Ј=H+=p,�c��ƺ;��}~��6��p�<��<󷼼�?=�MX=[��<�����N=��@=C~�<�5����<���94���k=����Pc,<�K�ViO�JM�=�5=3OG��<�B��@Ȣ��=��R=2O��B��O�X=�ͼ&����=�(�;�?P��?<��=�5k]9�?�(}=���<7��<�<?������S��nP�<}�ݼH_2=�0� q=���3�]�s=\U�<��D�6q����< �=�糼&�p�]B�6��|�����;g�ڼ_'м}u�<7P���C]�h9�<���<���[<�;&��;�
���׼ǘ7�;<�<�y�;�p���<_����<'r3=;�X��e򹇀���Q=�wtP�)�
=��!=����&<fr�G3�<b(�:�0�<�O��6V=��~=N��;&j=�� �p�%�!67������:=o9���:�h��	�:�S=�_�<[g�<�=n t<�}�wk2<EP_��Q�<Y7$=>N�{�f��<T�<�R�;i�8<�*�<z�`��:	<	]S��&`��BJ����<��*�qT.�>8}��ˇ<���<�|�<��'��$�:H�<�ZJ�/���3[�Q�����ַ�dZ�� �\=��ׁE�`�m�A��ڙ�C��C�O<�6̻���;E�;/��<����Ʊ<�Q0=�U=q����0�g�I=K�	=�7���ƚ<r�
�|?:��;�'�<�;#j�m��G1�<K�=>����n����M��<�Ǽ7����׻"�	;7=G����۵<��Ӽ�x=�<=���<Vj���T=߭+=��<NN�JᄼwJ����"����u0I��ۼ��Ѽ�<���;��μz*D�Ի7�g�e�2�!�[�<�E㼉�����<��,���K=1�ͼ���(���)<]�̼��^<��0�Ǡ�={�]�i��AD=�;��z��m8:�4�|���*=�;<�U`<Si�;ŎW� �P=ǜ��q��wb��#y�x�����I�Z.J�Q>=��r=9����~=��7<~F�<1
]=(]{����F�=BP*�e�J�z��� <��\=�*=�4=�o<YQ3��q���:
H=r�=:��<��ǻ;�s<�A���3m=@=\�19���J���j�r��\N=1�=�B=�S��O�U��噼iu=^2<�am<�`=�7o��R�"����20=� <
=��sQ������&1�ؕ��6���v�<BÓ�&�U=�{B=�@>���k�ǽ��� B�t�9�x<j��D��<���ck&�A��<˃�<��<i�<O\b��_�<�{=5m�<p�Q��y<�_����'���K<9�S;�)N��`
�t�=y�uJ9k4E��ͼ���<�PP����D��<x��<����냽����U�<B�:H�-=b�J=����[�üD.�BJF�.�=�D�"S=�g����;���=� ���<�.���A=�����ü4�м�5/=��w=�^=��U��É����I���kI-=�a`��*ün.�<�/��Z�����fl=�V$=�<-N��������<|eC�k���|�༑���e��<:�9��E=҂�H�<�����;�!=��=o�"�1Γ<�k�0v�<�
T=RB0=ɫL�"��< ��<�����0����\�;e_=�;�<Q>��/��0���Q;!�M���	=M��_R�ݳ'���=�t_=@bN�u|F=�1��x`=���<��@=ϰv=}����iZ=Bo�<]t<+��1�?�p�k���?=
��f��`�&{&���<�A�6��<y:�������g���'=����		<|�h=������<�B�n1<� =Fz=h?���)<�cI<���;��4d��&)=E�a=:(o�����j!��fN=z��#��<;r,;����Eo�����w�Z=�-�7�<�;�;�⸼m�;H�q=#i\����;�b�<&戽���)=6@w=��黉�e=ua;���9�T�>p����h=��<�J3�*=l�n��	�p�;G�)=h�X=L��=���5��]4J�_=��<�Y!��;���=>�.<� 8�9о�_L;===��;��X�(�q����>��<ח,��==G�=��+�.uF=*��;���1o����<�O�<��^��9=q�����&[=�f=�6I=V0=��-����"�.�Xོ�,��ҼFI�<�x<��<l+�<d��;��	���,���k:=}��� ��D�;��ʻ�;<S�K;��	=��z�<�Z!=���<�P=��M=�O<RU���,��<��w7=KP5�Z�+���tL��t�=ɲ=vFV��=�پ�/�;��M��F�R�����<*K�a̹��_D=��<�5���8=�P=���<�n�{z����=g����'=�40��U\�>�E���Z=[<KJt�`��e�����<-=��8�2^ۺ�_m;f�=���<t�<D=�8z<*�=a�e��@,����;.q�<�M���>� ��;���<�>=V�S=uZ`= �<�2=<��@<��/�<v�<'4���Io����lf�bK=�~�Gg߼7�N;-=n�V��Ǧ;��=��������=3OW=*:;n4�<�T������h� /�<-��<p0��2�<໼�
�;"�;���q�<W�3;[N�&�м��.=��}<�kA�=��<m~>�ք���f=�dU=pC7<�g=�(�::Dż$Q��#(3��}߼Q�6��_=��j;7?<�a9=:}����#�:�.�a9M<w�=J�=1zͼ��+�T\�;0�VR8�@i��`=�:��1e<_ M�y仼0�4�_�=bP@��=��F<b���[�� �<]���;+;@/�;�\�.�ļ��y��1�=j��6J=�.n=�8ἂn<�E�<�D� �o�N��n=^���%�Y	]��u���&<9��4=y,>=�f<�Yx�mӼ�G�<�-F<�)c<�4=��=��:K�)����<�����<]�N�,oJ�
;c=scH=���<�^�<�D��^�;F�:=.<��={���Z�{�x�.�,=���ϏJ=��;ܨ!��`�<J6y�k�Q��d�KhP<���<���;�
%<H�x,	<X?�˻[=F�b��<�~��$hQ=�`�<��7�fG��{=��^���;�皼�U=��=u5�<�#M��J�<�!/=��D��a<���=6�x &=�d�<�i�0��;,VE�K@B��t�<����ޅ��k��s�=����hk`<��r�� :=�j�<y�Y=Yn�|�K=��^�a�<��ļi?��'<�R���J���<�l�<-C=0\���\�Kآ�*���s=�M�<ے�%�=�ȑ��9 ��v���R=h5��&=�#�=���}=>/�<��./ϻ-������<�pN��9o���@<;��<�������Z��dx=��Ǽu���/V�iQ��� `żi�<���<2�;a��<~\%;��2=ȑ��U�
���<-��	<���[l�����K�|d=�^�Hױ<�f=�.=4=U�<ko�<.;=�5%<ފ�<iP>�d��հ��ǽ����=j�5=�`�EY��<�t��O�K<G�C;� =*D�=Wj~:ݡ=�R���?����<� ���<��v��md��?��>�"�(�z�����a�ռ ���c�ż�l4=DF��=6=H��P=��j=)H�<7}c�u�`<�
=�۴<�м)��;�S=^;<�����<6�式�7<�L���k�� �\K��P��"\=�}c��&�A�7���<��M=E����:���=4�<�=��T��>=fB=B�W�<H��8�>��?Q=�}���C
�R�n�`"p�TEJ=O�*�W�=[X
����}
⼋�=}Ӭ��== ���]7�r�$=�~�Iڞ<A~	<�=�(R��{dD=�^=9�<�0���V
�*�;� ˼�����<=�:Z���ػ< �Ļ�[8=�Y�;�q=p�<�t��:��I=� %9��e<�&=r���#=�P�Pg<`0�<"3<.��<t2��p���]=�N�<�aZ==ܗۻ]Z=В��+8�:\粻B~$��z�<9Qf=TX<!=Y��ԗf��@M=��n�A�@=_�f=]�n/��`V���żK+��T$�^C�<�~v�����c��;���"�;4|���=>5@=�D-�����8<%56�b��<���=b�<}pW=B�</�U��,�{=Ic����9����f�껃,�=�����3�澤��M�����;�;�<�|�۬9�j���M�/=D�� 
n="�<� ����q�=)��l��@L����k�i<i=��F=K�u����<�_��9����A=�Ɂ����<b9^�|�=�j��|b�|��������˼��}����Q!m������<
�\=�<�}�<�T�<׸e���L�Gb<
�#=���;ؿ?=�X��&bм��1�u��W4�<�fC���ú���<VE�W���W���)��ED��;���T�h��9,	J��TP�TF=���	8���IX�E��:�Zb<WȤ���<z	c��=���:�f<���:<�_�=�;=)Lݼ����Yj=;�:��(�a�N=�1<�
n��%(���.=E�f=�!]��?==�P�<��s��.����Z�9���zg=�ǼP0���:�%������I�ُ<�'=�f5=�`�<��t=�P.W:�$Q=�.i<��c�<H|���d�9J=�Zt;�@+��?�<����~ء<��=�R=��M��U�<� Z�cU<�P�X>6�;�<�>�<�O:����]=HO%=���<��=d:�<��߼#�;��K=/9�����<�] =t�=��M��-��1s=<��:��M=���=D�6����5�����Y<+J
<�=qѼ�"*�s;*��=��<�b=մ�<&a�<�����n=م��nv�<e�Ͼ�Ĺڼ^9c<-�9��ȋ��/<�+==dJ=`&��� =��H=cH�<'t�<�f�;ni��3��^<TuB�V2$=l�ǻ{��/�<��:���=qҬ;��/�JO��^x|=�GG=\k=���s�<L^q�&�A�C+�;�cټY�G=��?=M+��9�oaf<�e<+3=��+�=��R�lgc����<���;)u"��G���.D=�[=
I8=��<�[L��)Y�����S=��F��=��<�x@���'�i�ܼ�Q��o����^��t�;���<6=4��ǟ����CQ�9|�=�f��u�=z��p=��l�����Fh,��{$�,�U����M}�<�+=���<��o=�2���(=��;$��<�ۼZa����(<�~F��xU=�E��2=̕������_$�T�ۼw��;{�A��O=��<���*<C�|<�0�[	=ڋ�<�.�<�<����/� �ܻ��8=��=�G�1�W<0� �� ��r=����WI=�5	='�	��<;:7=��x�/�e=����O��u=|�<H�3�S�]�S��<�9
�Q�<y=�5q=8����'Լ��*�*�л0��;�M�Y�
<�i@<��M�L��<p�=m�z<� ��)[���F���<T�'=��<����.����&�x
:�8l��=�]�F�ueg��/=�5��]��r=cX�<tF	�F���J6��W����U=Y
[;M� �t�<#s�+�6��Ju=�*= �a��-=:��;�^=İ�=Ka[=aƊ�H�+�w�n��Q�;��V��9��A����<���<&%W�������<c�Q��$}<
�/�B�M�,��n <��g��T����/�%��<����`;�/=$�H���H� =��B=�{k�?��;[C�<R����F1=�a ��?B�,�N�f �<�ET=^�-=NO.<1�켇V����ҼS�&=�b���<܈5��\o=��:�h=Q�=��L�';��<g�S����<�@b=�+_<,��<�(�cy==x`=��*<�/(�fJY:�,�Ή�<�r5=D&��X�; m��C=�<��K��	�h�=5A��N8z���/�>&�1o𻬽�<S�=��c;=Ҭ<Z?g�e��<gj-�w�Ҽa#=x�a<�*;ǲ?�-K=��ܼ>sP��g=��?��)=���O�[��&�;��������=|K�;�f�<5�*��a`��3V�e��pb=Q{c=���5g�F���{?;�� ��e0�u����V=�r��~-S�̕,�������l"P=Gr��(�+�?.�<��=��/=~���u^;�U�<F*�<~B�=�Q���n=���<��3=�;���e'�FG4=\�y��b�M��׆<M��=�D==C�<�`=]_'<��⼊��<eFT�Sѻ�M������<�H��b�
�fy�>=�	n��,�<=�	=����.A<��p���<�=k�����R�#w1�"�ϼ�T�<o��4Ǽ���ى���V=k�;Y�&Z<��<�#)���=��<8�M��%a;�-�=a\��u�U�YgV���a��?�����ub��=��c�!9��e��2�I��;6�����.}M<���<ϫܼӛ!=0��;�=m�E2��P��<C��<�C����뼸�=�_��=�9ļ'�>�T�!=�|4=R;*< �*�;��/mX��E=�m��r�N=*�<��<��r=��H��<N)��U��֍�n��<Wټ�� =_Ny�h &=�PC�(A=���4��<�|G=�=q����"R;V��I���<�;I�;Q9����;�-=��Ї5����<g%�:c���K����;��=�4�<����S^=\����F�<�f{���~�;=� "��KM����������<��D����5�=���<��j�����a�=qji;����k��}�ʺ3ZS�����&I9�7�&=x'z�}Hc��f<�"=��;�1=y<ר������=�� $	�(@:�o��;kF=[N�sc�͒�<�[.=��[=im�<D�=%�j^��h�<�ټ�jt�[��</�=E�ٻ��4�±�<����~��<A�:�-���=G�d<��;�,�#5K�EsM�K�L=�<2���U�'�O�&=��\=Ar�}�<�ļ�8�2�<�}�<� <��^���Y=�XҺ�h��/��N�=��M=f�;�E7=[��<%��;�jD=�C��&� =��¼�QϼUjT<V�μ�#<��t=bȜ<j>d�C��7c'�K��=�<��G��Y_�#u���S���(=r�z���]���<[���m�<E�f<6q��5�N=��������7�� =��A�k�0��M9���B��|��MK5=��5�,|=b����~7=�a�j��=^���xB�<�Ҩ��\�;ד<��n�t��;���N��<o�,;�n;�=GC.���Y<��"���i;q$=��(<;~���<�朼}.=�=��F<#9F<@+㻚IH=G�H=?M1=���ѭa����<�c�:�/Q�@�H=[`<���<�ɼW��;�@����,� a��D�sYɼ����< ����<2��<m�+���b=;�O�^o@�[�<�=r�2���J=?/�<;W<��Y=�98=�\��5�k���v=��t�V�-=�v�;P0�O^�a�=@\�<��5�i��;�Th<\����:P=�bs=P�=��<<�Ѽ��S=B=$'[<b�/<[�l=*s�<Un=r��TS=���������>=���;�,�<O��Z�<�ӑ��ϸ<Kd����<��U�vW=�� �� ��n=6?H�7���b=H=�#!�(���B���<�)]���[�qXB�S�<g�d=?�u�"�:=����0��V_���!<��&��j*��_z�n�g<�Z�;Jb.=bZ��!:��o��П�*E+�Ր%=���;f^"��qE��|��Y!=�<="���M=��Xψ=�@"=",=�;:;���k9~=�,�?Mp�����o�<��(�}l������7=ٽ��n^�D���Y��<�P=
�J=��Ǽ�B=��ռ���<?�<�M��y�k�; E~�V�Y��J�<�J�z @��7=4�#��c|�*0�$�-=5*��E����<��+�@j*=5b#���ʼiK<<1���@N=��<`��t����A=iP󺌨=�"�;΋D�� �<��n�v����:�����T�~<���<@���+�༓�/��#�<�K:FC=ۏ^�<G=)�a�^���OZ=ۡ<��h����;���t����p��֔C�X�;X��<��=��I=�k׼�]v�"Ҽ{ޕ9e����9:=�J�<s������z���z2=��z�\�)���LV=���=�ק�f�W<$��;z��qD.��Z'��J�2wQ=��<Y�<r��M�d=*'=�,��s棼�sG=�an�.߭�>�6�:��h��DV$��u�<q�x��M3=34(=U�<�1=1�R�ҁS=�D��e���5=|߼<�f=��<J)<߿�<�/=�: ���-=��߼[��(D2�"f�0����]�<p�#E<ֺ�<�%���R(�3c=BS(�P{�����<c^�,��:8X<�+L<�?��@<J�D<�׍��Tn<l*���*���%=1|F;A�,��v¼���<���;Qi�Z�}��<�?=29=��B=�-񻈘�<W�A���C=�2���+=d2�+��;1F��=@��]����B��XN��QO��5�cm-��:=��c���'=�)J��(�;��E��:4�ۼ���t�K�	�"�L=U�=�i�̾�L�Y��<�G�߻(�[�6=$A��'m�o�<K�r=�Z���@<j�S=�(=�F���*=� <���<x�ܗ>�,�ɼ��`;�=i��W��ʏ<�Q�1R��U*H=p�=�r��;(�W�/>�����<GM�<�X��Bk��J#==�5��<� =j*ȼ�r�;NA\=���<���<AX�<t�	��އ���;��t�O���$� �j:��u=�p�}5<�����<B�;��N��=>�<��;��<�@�Q�<A��6�<��-=+uм�R�`�S<��F��)�< �;��<<��=�-�<e<=)�=�:7��/=��&=�
��652�Q�B=U���<x�^�<�Լd c=l=��/��;�N=�40��.=|D2<2�s�"�<�,$;�$��^H�P0��E;�|ͼ͆��7�,=?�^=^�T� a���#`��L=�r=8A=�˅��5&=�9==��<-:=��I=�|p�+F_=QŁ=On���<r..=�Zy��τ=\Y�;���РV=��O��պ�T��;sy��+�h=�r�<��,Z�W�<����w�Kp���<g�9�A�|��<�mg=5)";��d15=��c���?�pƼ��<=˻<������f:�z^=�e���N�)�H�S^{��aH<Q�?�A=�5�;�����%���&3=��+�TX=�h��j�¢i<�JüP@7;�Tr=^��؎Ǽ8wV����2%�<Ce�<��"=��F=Y;���'�(��<O�=M��L���A=m�c��5y��3�<h�A=A�º�y$�l3�<���<eN��}=/=v�м��<&�`=�K�8M�1=�=H�=nay�to�<}��<�ۓ<�0���"<�q�����|�=VѼ�3�<K<=��<*����a�����м��H=�t�<�0���D�_�'��s �U�*�)�ͼ/#=j\q�;HM=�N��jj;���n��c^�07��P�<ï<wހ���=?ʉ<��P�$/켹�����:��ܼ��;$�<��D=�@���qȼ�� �<�����Ҽvm/=k,�;�}�<r�׼�^~�qDo<��ļWz<3[��|��K��;��3="\&=٪��[@<���<�9�f�<�uR=Y�+��4߼���yx=�T&��Y5�^-�؀=)tü���=���;#b)=��޺���<��������t3<���[J�<�/ ��4������ =O�4����<��^�۱6d	���|M�v\=��<����r�����=f�w��޼������;TR-�U�?=��ԼR}�;��$��������;�Wq:������?v���７F<o\�;��==��ȼ�vd�k?��.g�q�����NN'�t(<V�A(�˥2<���-s��^&=r1D���*=���Ɲ)���s=F<$��%�<��C=�@,��
k<j7N=��"�~:=��=b�ϼ� (<���1��2=]�����:���˗=�C=<���]<B�6����2<� '�i#c;C�
���0=�׀=>��<�Mo�z����Y=4cK���鼒�N�i�E=Q_n=�l?���I�C�<�d=��a�k�J��
�%S��W��;B�h=/��<X�<���Ǽ�<ʪ=� �<���vP="�<��R;�h�<#t��x�i=�w��;-0=qu;��<� �<S'&<�)=Gl=�y|=�_a�kF�=�Q�1��<��<y�%=� =�F8���ܼ�q;3�)=�=��c��#:i�=��Q=�d���S��ʜ�N�=��� <��<ix��B2=w9=��]=Gp$</j�+f=�G<'��<�!G��.L���<Y-�B�"��A�<�=�Լ]	�;��==��oHx=�e	���*��@<�X=�옼z�<� ��7<�s�:�=}�庞�lϦ<ۮ�<H�5��g�=��G��n6�� 0=�J=:�}�(��ՋM�y�.�K=J�M���<��Ǽ�Kt�kx�<WNj=�> =a��<u*=T���=�R4�,�5�w�<�Gb����w�==_j�^��[�;�<\S�<%��<ڼ��U��fU����X7=� =�e�9�B���<5��!��T�=�<�<xH�E=�mԼqa�ɤ�<���<*SW���ϼ߈/=�=�إ<=c��˻scF<4'=j�Z���4=|����%1����	|<U�2��.=��[;fZ =f|<p�c�]�;F��;�.<�_������[1�<S>��z��䬼�8�<ջ�v���}�f���*�މ�<(�=�4�S�]=A�O���=P�X��������]�<t�;=��<�!(���<?�	�,���l�@=5Q��=ճ�;p9<qLp<��u�='QS�;t=��1�i�����U%�<�����<_�h�|�V=Q�<F<��c<pH�<C���&_�;K�<��;=ִ^:I�#=v:��*	�ע��������?��[=R�\;�{#��5��������:�M=wq�����:��<C�j=o2�.�(�H�`�n�0<�S���r�ǘ=�� �,q��fۼ�%ۼ
(����D,�=��<4��<9;���<�X�;�2���j=61��Z���iOP=ଔ��>=Dg�ל�:_�=7�,=����!�r<��x=��<�i.���(= G`��8*<%���(7��'����}�=O�3=���;s6�<���߼!3=.6��hP6<�U�<�������%�<[f��ӡ<��G�Qt=t]o=Sˮ��o�<�� 5; 8��mK��̆=i�+���=��8�&g<�̲����<
=����_��H,=���{���e�4<�d���ܼ�}�<������Y������D��<JQ= P�;���x�P;������9�&ZW�Ӳ4�6g*=��G=�&=�����ƥ����;�ؾ<�XR�,˼/�����l<G;���h(=�)��3?�V�N=;{Ǽq���0���U�"�S�����!=��'=	Q���7�
%�<�M4���<r�����=O�_=T�Q�d�%D��mw'=����~<�<�C�.���6 �;n�cx=^[���/�:@�<��y<f2���Y;-�<���az��K#=�6�<�M�<�v=�]=��<*B���[��k!=\j��Q��<k*�<1<u�<��_=���<B�Q��h��@Ǽ�;��s�@/%:T����<��j�g���d;b/=�7}=N�f= ��<{��;�"��jTx=���<�-�j�����j=��=�P<���!_��N(j=�P�h�+��z&��Є��Pp��3%���/�X9e������<WwA;���F"_=�%�<O,�<c僼���=*�
��� ���B����<"�M��*==*?X<�ͼ�O�<{T}��$��8���H=CE�p?�<�|�:��=��ou.=z-2={����=�@=w݁<Vc�z�=���:���k;�lܼ~=�p%=5���K<�I�~�u=�k˼��;�F,=4K=A��<
ux=`wo=�!=Up;=�'x��&k=^�D�:7 =��<Q"��:=�Z��<�n����A��[[��J����!�9�V�쐦<X���xZ�K;ټ�B=���:�?���L=��	�@+.���h�0/z<�f<,+[�|�λy-����Q���=�x�<f�=h�&�\M��g�<�<�<7�<� �<�4���9�G������8_�<�4��9���<�[== �i�("�<a�;��<��ۆ��{��Ab:.���K��:=��c<٠��w�;;��Q=�F?�Bi��5���B��l�����Z˕�?��<��F<��2��
=|�y�t�]=�}O�#Ȕ�A'%=��������xw��(,���sE<Zoļo�o=꡴���k�5�;=��<�|�<�%G=ť�n����R�<]�<��	� 9�Ue�=��<��+����;��C<��;@�#��gл<Y�kz����K&��Q�<r����H��=���<��X=�����<�!�;��=9x=�P<���;N`=Bk��ي�j��<�WW<�;��%=&��=�+=��e���<o2��rHS=�h^=���1�̼d8?;�>'=��<�����<�
p<��<����*��߫�<�V�<��<�m����<�QG�7ﭼ�4������I�Hc'�rx2�D<7=7�=�G\=��t�м�.K=Md<⢼v�=0�<D�=�$��	�9���%m���a�5�=�n�=��u"a<[`R=�~ =���<�;I��Z�ᆻI=�����O<V�󙌼,v�����)+����L�����<e��A�=K�w=UE+=���wĐ�����A�N8�0+;�ֻ�r�<\���Z��#��\ǻ_oٻ_�4t2�# �2�{��Я<p�~<��������ɼ�i/;"����/=�!�6ߌ=VH��Q�<M�<Z��M�^= �"=O#e=&\�n�ܰ�=~VS�]�w�����лƖ<��=T�i�`����w��-��=ED
;Ȑ8=�q;��\�k��<v�F��s<D�<�Q�<��:=��D�3=��<ZNQ�����cG< I�<K�)=˰�=m�Q=���gJ=6���S� =}I0���Ļ;�/��^�<?��<9�<̭=��ļt��<�󼧏d�o[N=e��<r��=p�8<�����@"<�X�-*������=h�>=V�i<P�$�3���ɼ�-��=:n=5��<�%����(�=�rj����=��Uw=>��T��<	WF����Db>=ZMF=��=9��<�+�<�s4<s�<�Ր���`��(�;M�F=)����?=@&�<S<�<�л�;�(7=0��;�T�
�=8�ҼO�߼Edx<ڝ�.��<:���7=[�2��r<�#�7�"= ��<�i�D��;�$=�H�^<��0�N��<c�F=!��<U�b��^�<hrM�4��m�Һi�;�9=�+���7�:���;�?w=�;:�\ E���'=���<P�����
�<�y�<kK��v�Ѽ%�I=XE,�o����W+��[�<L��<��
�UL8��$�<AG�;nn=$n<gE?<1��K�����;�������H�)�̼{�<�S+=�ϼS�)���<��A��=���<P��P�4=�b)=+�x�H5K���
���=gE��Ɔ<�'=�0=���<k�-=�<e>8�y�8��6R=���<y������x?;����ȪI��Yd=��"=d�<���<N�;�;EE!�^�=�Vk��?�<���<cTV<(^<��F�m�_�_�S����<|J}<7V�<<�'=������I��;.�����u2<�=��v;���<���<��O�92=���k�=�a��� =xR���=;s
=�/��&;;2tҼ�ż��Z�ȉ&�0E4�9��:\B=u�p=���;<Z�86F=ڞ�<��=�Ƿ�d��;@c�<m3���M=�T��물��Q=����O����0��(�=1�x=��.=s]G=���lڼIbo�^%C=LNt��R�)�[<zn3�1�;�B<��<����)�<�:~<4��</�n�(�<�=q��<��]�����=y��%�����?:�n�7U%�@L:'�==�#.=��=L��<��s=��K�Z����`��cS;���;4�K���=4Vv�l��8�SP=��k�r^�<��I�럖=���<�8=��=���=鼖�ؼn�=�u���1�<� 2����Lp�<��ͼ�>��4Y���=�m_=|�0d�;w�+�$=��G<L��&Q<�I�q��<Ԡ�<ua�<8u=��<��$=b��-;���<�%6=FЪ<L�r��+Q=6�q��;}�ټ��)������>�:�	h<�RY��r"=�1N=���=���<�Ű<+�;(�i='�������P=r$.��?�K�=�X�=�1��	a��t�?��)�PEJ=��"�[]=��}��}��!}R��%=p{g�0+j�� �]օ��}�����;�6ۼ��N<À��h�;�P�<����	��e?�$�=�:0��'��|�6=�e}=er=c{��1x�<�p�<i�2=��b���/�X]r��h9=�N�<�<9�w���!�q=c�^�'�;�h2�Z?�7%�9:C���j=�8���)4=&�ü	�f<�?��i'�WL=�B��!ۼ�雹Vu�<�>;W,��0��/�<b�=f�(�ۯռ�N��D�6�4����<��:=e�[�&ޅ=���<~|�<t�#�"�V=d�=0���	�<�]S=DA=�l:t�e=o=>�=&�#=R滵Z<P�y�ݼ� �;��!���!=xZ���:�;��<q� �g���My�3�-<v#V=i?<Dp�<C:q=�缚�@�*��;�����U�ֻ�SU��s=śm=���;F�M�I�=�^H'=.,�<�=z�:�)޼bs�<2J�<D�K��l�<����K=šn���
�;=f4=�l˼����z?=o��<�^=���<�k6�Yo������<,�j�\=w����fP=#�<Խ�Y�-��J"<��߼���:��Q=����	[�Z#=��9���$=9��#J%��S�<3g���f��<+��;�H��:�;�h=�:E�fX=C�#<�����ښk=�O���3=S�e�"Eּ��;�Z=�Ĉ��ﶼM��<��]=9���t�;r����=���P�7����<:,�<i�<���;V�7<��C�������</ؼ�3��';�<}3=�[�a�p=	F@=�l2;�1O�]�C;���o� =v��<A_<�*,��fM����=ӱؼqZ=�ulC=�Ǫ9̝=>m���w��,_���ϼȿ�:g�B�v�߽=�<dG��{ ���<x :f';��<�&2���e<E�<䓘�c�f=uQ<*^�<}��<���3�&��8�����Y=#�<��h�z<�]�<�SB<}��:�ak=��<R}����=���;0ʧ�xH�<I�(=�#D�uړ<#|�<��;�^J<uK���Å�g�=��뻯aj<RG�%�s<2)=��.� 1=�Ԉ�z��<>���1S!=�)=U��	l�EH���e��EM=�nü�>=��)=�1&�;�H��n���׻���KA:=�I?=�N�a͢<���<�ܕ���==�1=�h���&��Q�T��E;=ԂU=��<���<�"�;v��;�v��Vȇ=�5*=��0;�Zu�8�g<�=�����	�;0*L=Lm>��p7��d�<i����U<��5<�K���$�ÎT���>�BbK<%>S�0�g��6�3��X��=��7=>z,=NV�<f�7����>�<d�u�rj#=&!�L�`<�=��ռ�;<��@=�/����g<U�>�{�S=L�l�R�2���μ�{=-�켹�E=ȥ�<5j=�x9�x��;"D=1��w9�<H��<�hQ<"E���}k=��E�m;B����&�*=��)�q�]���N=����|n=�q¼�*=�߼�Q��ѭ�K�<6�v=r �:Юf�}
�N�=��<#o7�n�;���!>�<�5��0T� �$=1�i<��0�Ng7=4]���o�戏�pZ�<Ҷ>=�W�&�=��<,�x�F�T=1��<!)=Uj7��t��n;���;E�C;��l=�?G�=�g�D�dq=�J?=�+	�r%r=��	�0�7=�ӗ;tʹ�܂ �0:l�Ē�;X=KP<�؝� t=5\����0�S�u?y���^=P}>����^A��Ta�2_=GV6�EH�<M��<��<�j<������<�pD�bߔ;kwM=`���X�����;���<�����4+��;=>�<G��"�O=E]P<�M<�ou=|����d�d{<��<�/z�B~�<Q��h/<L~�<�E�+�+���<��E=��G<7\��)/�#s���O�9�=t=k6���[=���<���<�`���w=��<߰v��
�smx�K8�;�-=KJ<���<�q�<��ɻ�=����r==�*���;Y T=��\<J	S=��Z=��9=�0�;k_ȼ!Fz�tg ��;y�!Z$��I�3=ʕX=?{<�
����m�V��!=`>���<�ԟ�V�<Zʦ�O��<��=\��<
|��
v	��8��èѼ99j<��e���ϼs����^r<��^����\e<UX��k�漏�0=�c=���;�)���i��m�<V�"�DA<�=�\f� :�$�c=��6�	|������'{;U��9F�/�!�Ts{:�]k=Iʠ:
�:m6���?���i��
C�K�=o	*=2���R<XY�:��L;$�<�c����<�bH=�P��[�m���!��F!��ꟻ�}�d�=pX=�H2��><*��<�gE;��s=��>=v�Ѽ}�5$Y=�Ǽ(I�<X��<�8k=�FؼJ=h�=�o\�|�Y��L@�Ĕ�<6M< �@�t�<�@���/��}��U=��̼<jD��T�<=�Ƽ8k*=���t1���׆U���:�a��s�$&�<%����^����<�6_:>�Ǽ���Ja*�D:j=��=�=���I9Ҽ���Owf=6�.;���<y�2��J'=� =�L=����U�<+��ޯ�<A ^�4�x�`J�<�� ��(=j��<�z�n2`=T��;�=Yd=9*=�i�;K�?��g#=缶;��/�,��;�h@���<��=��=?ؼ�=�n3�1軻۠[��$�K�u=��F�<�=�=u�=>��ǘ=6�M��5^���M��{º�޼x�ϼ�I�Dq�;V���F|�<c�o��<���Yq��YX(���D={�B=j�������i=��1=��U=eR��b=;4'=avl�}�`<�W>�2�c=E��M�9<���\
�3a@�m�D��|	��N=��,�����v��s׼OE=J��<B? ;�t�<��n�8�D���3�z'=�;��!�.=�QP=��R�VQ<=���<o��;�K�<ZC=�1���l�<��=|��<�v�<�*㼀O$=�B]�w�;t&�`g9V��<�j<�g�m��;Q�=�!�;(β<ɾ�<r��<qu[=�#G�V^S<`�8=K=}@^��v�<�m:�%&��4Y�]Op�ҝ�y� �bۼ�f2��A�0D4�N�A��uH=��#=���i�T<��6=X�(=�Użܨ�<r|<��Z<[�?�?~:=�s<��Y��)=N���M<`��&�'=tQ
�D�q=L�=��\����<u�	=*�~;��<D觼AP=��A�dKI�ܷs�_�=��:�����>���׼��<=��<�=���;�g='�=�����u�$R=�����(=\�3<�i�<F�W=����<��ջS;=C>�K�ټ�s%�8�=��<1t�<r`��I�<.@�̃��AC�K`�<R�H=����{2��φ�<
�
��~�<��=d�M=��D� �����?=&e�{�n���Q������9�����p ;-=�X�<�QR��5=���:�o_==y�n<B�D�g���qɺ��Y�VG���N��"�=��M�+uo��ט<_�<��<gp.��t2��q�<;ݍ�>-=p�<��2�&��>?�<!��;EW���y��&=��7=����WL=~Ƴ�D�r<��3��?<�{?�Bq<=�c�;����0�W]�c��:�
�>�t<~��<_E;�	$��฼������h�q���O=��<=hɏ<t�?�?���"'�����V=���<2}�;�Q���S=��<���X=S�g���)�"�c=;����2�yjH=3.|���<ܯ�<#�'����,�2��(ļ�_�;��=�F=���9���0�=�[�<��A=v!<��G=���<�E�<�UI<�~뼯�=1�O�d*��}K=���<�\�n�<�Fb=8��<c��<��������k���:W���A�dZ4=�J��%��b�1��;�@ �PW��;�S��|�������;����,<���~����<	�<�� =�2=})f�?�=xD%�7x =�(�<���<�C= .&=m`��9 �ePἃ�5��S=I�R��n��1���:J�0��_4�=&���@eּ��)�^�a�1��<���@��U%=}�:=�9�hm�<z8C��4y�t���k<Y���w�<*QT��B��3�T=��<�Hb�,.�����\=��iz�<%�;���7�[=b���;w�м4�<,,i�`�<��<=�3Y�J��<�w=z���<�<��/��g�;��<�.��Q�A��@�<=NZ=�	?�y7=_�_�!%�;ͧy<Y�-�'��<"�»Mj���=X��Bz=�@���t���<�T=ujg�O�Q=�	�<`��ui3=���<d̆�3�<V�S<V�q=J�=�{��WX<��O<9!����!�<=}��j<<R�o��G�<��/�t"׼�<��<�=��<<n���C<=�mA�NY?=�QJ�w�=OV�;o�+	�.jI='c;Kü�=j<n�k=�S�P���P����;K{=�>��o� =�,l����<�m��fy�{L�׳�<��=��=2d�ɷ\=ob�<#�$��@J���;yDu���m;2�$=�.=%H*=�1�;�c��%c+������5;3_=�Q;�؉<��W�<�׼3=�T=���!X�<�^�^s=(�==˻
=�H�T���U=a����N=�XA<zE=��=i���4�<b�=O��<�b=��Y<�Ct<���8}��H���<�E�<�->=6g�;ٓ�<��7��zM� ��H��<1I��rӼ<9���6�<e+=�<�=�
���ػ�����&=5��g �4����e�=�'��Hڼ�<=��n�3=W�-�B=��=[���%=�.���\й~�<u	�����<�)=$k!=�����?��#ּ;U/�<7 k<b�xe��)=˜�(ӿ���L<���<��=i%��D�<!�(�������.���8�6o=�O���	o�hX��{:V�d�;ܜ�<�<�W~<��D=g� �Dr�;�h�<��N�>��<Aז<���<����#�[��ּ���F=�f;D������=�8�<��=~��<Y���i�����<�(l=�V5=9�0=9�`=l�zbP��f=��=��b=���<�T?���_��ۀ��<]��9NЪ<��?�4�"=tL[<�sU=����/�=P���Z�4�_=G��1�<���09m<!�ȼ�i�KȾ<`��<�-=��5�ID߼.�<s_=�;>�,�}��5�`�C����������˼�I"������ǻ��2=��,�e�<�W`�
:יѼ��)���;�Vp=�Ƙ<����}�#��An�K�*��4;��<m��m?M�h\=��r<e�<*p��:+�;�'=�+D<ؗ?�	9�;�9����<�N�=.=�i�<��;=o
���p�����QMO=o�=�#S=;#��������!I=֟=�C�3�	�K �<�/=��1=��?=Ps.=�H�<됃<KP�?�S���=�I;�P�=�-<��=�j�;��;�}=g��<�$K�%K�<Z���bL=t��;	�k�(�+� ��g=�A)�\���P�V=�S=�鶼��<:Z�=4C����,�w�"�������7=_ae���A=��H�v�(��ּ������r��� �C��s8<�#=ӳ
��2�� G;I�=��y=�����hW=�-��H��;��!=����L�% u�s�缗/�;uε��\)��F�$"�=D@.�۴�����&У���E=�A�<WRb=�$�<m3�������kg�<w���F4��ۙ<-��TR=���[
{�\��H�X���=y�<��|��<$�8���F����=��<���;m�<-���LZ�<�����<x�|=чȻ� t<���<,?��~�P=�?;�l��1���zO�^v�<n���X�<d�'��5�<;�=:-D=GL�<e�N�>'��V��Z����4��3��ڐ[�q��sh�< (�;�-=̊A=@�=�]2�c�F=y���<�'�:(&�<B�����\=�GT=��W=#���l��;�L���G�u}=?�j��$�<8f���G�Y?�aZּyX�U=<��7������%���R=	�i���;I���y<;�¼��R�m���H����<��8=pM�����<W[=,C=}_\��1��$7�>�3==t ͼ��=C߄;�;F�R�O��BK<�f����W�D�
<hx�=��W!==�<��,��� �9��4<ExQ=�R2� ��;��w��};���g��T=x|8�D����<�[T=Z�6�-��'�<�K��h<��*=6�м��+=ܧֻ��o=��q=��;��h�EA�<ꧼ�sO<��\=QA=�zN���<
�G���<�5w<V`0�$ϳ;��<ia�L1y�����B�� ��P�0=Ā��.7L=��f=U��;<e=�Y��>�`��CI�w(��B=<�<h�r�6�V�>�^�V7z���7�ϧ4=y/�0��<Q���=�1<7wӼ�H����<y.�<>M�<�X0�[nJ�{����8=I_=��=n9n�ü��� �,���"��ImC=��;��T�X���
:*:��Y�����:���U�˻�_����:=&�ݻhk <��'��� ��$^��PZ<�f=��;F�==,V�<q�<R�R�G:F�����en��T!=W8���;�V��ּ�(��m�<t�q��@;=5���S<<֒��ǯ��wȼ.�b=�<����<#��u�<F�`�\*��=��}���m99=6�8=�2��NR=s�=gM��uP<��	����+=�j9�u$,=4@�]G�<.J��&�(�!����f���}<�
�ݓ�<CZ�<S��;�7������;�iE��3�1¼����="�<����t=��u��lu=�l�������<o�����<��`�i��D�+��=b5h=�0H�(�"=�/=�҅�H_��_-R���1���
�D���I=H��<�#��%�<N�=}b�;���<QP �ч�<��Ӽ=��<�ڋ���<Vt\���Q������7<�=ĲǼ0��:�C����`.8=��<�87=ߨ�;� ����y���׻�>q=�����&={.1�b�{�<| ��<&:�#ƺ��;��߼@�ż�G�9S=�H{=H�S=�Qs=�,�<W�<�s����<�<1��x��Iҥ<Fܝ�(>��Ćv�́�<рl��j�<���苼� �ʢ���Ӡ<U��s*輠�.=[�;f�=n׹<ҟ��!�<k1=�:e=N^��A|<��Z<9L�����s�<�=D�2=�{C=�V[��)L���N�<�QZ�_�#��&=�Vq�:�P=��u<c� =�p=�$�;M�=%=��x=~�;��oA���<��i=��&�xD�<&��<�Ā�Iۼdف<�.��W�;6�t=$�0=*�=�p#;/�d=��4��,3�U�$�W3'���<��=�������=df�E�p����>�v<jL�<L�f=_�=+V��]�����<�k��-�<�.8=9,�;���� ��:m�N�nx3=���c�<��N=���<�:�<h'f=���<5E��"`=��a���p��0�<�B�A+���<�ͼ��5<�)��B=�p=��� #���s�-�[=�RD;l�4<ZN[=��ټ���<����4�^#�� �;U:���&;�Q޼���<-�N�6m[=P>�<����o_=���<���<�<#if��P����<�p�<B{o=��6=������S=��a�r�d�����<�p�+*�<��K��?=��P=W��<�&*<"\�;Ⱥ��y=�%�<�t�6#�pS����d=�=�0��<qμ!�=3��v=7I��Y4��4O9��;���;!T<����;#���Mۼ�so�jj7�/��샵����C�=�
F��2�<�o0=W�=�c"�6񻂶Q�M�=�������;�nB�e��ze<<3�ɼm�T��f�<פ���^d=K��&=�<����J�e0;=s����5=�����<��ڼ��.�^�5=�4X���b�^�żN�$��#�8k=���<�n3���w�a�\=�q��[�J�R=pr<Joh����:<�&#�����E�)�4=�o�<��4���X=\� <c=����{$�zL���:1Ʊ�x��<�1ܻj+�;�;=���l�5�r�<���<]�<vk�;����<�ge<#<�N���D</) ��7=S�<�g����c�Y~�<�����<�����&=F8=��1(�<���<T�[�$����ѼHWc���:�� =�^��O犻%�(�3kG�8�üPo<Sp��H^=W`=x���1=�*d�|z�;e����^���=�B�;N$ �V�%=���<��H��D�	����_=�����$�;�F�SiW<ǧ�;_EǸ��<�b�=��V�W��<�$=���<rd;����9�;�֊��ü��X=��N��Y<
�,��%�'���1QN=��<F�$���Ѽ��<T帼� �-"<�Jq<e=�w�<E'=dJ��I�=��<n�<�7D��<��h=m�<B �SI�<c����B=}҅;cӻ�,�x�<��<��<�/�<�ݻ����XY��Ag=� -=5�G�wqU=��<J��<�f���g������9�,̂<� <�Ѽ<�Q=�rg=qb6���3< *�aIW�2?M�~��6��5�1=z�0=.Ɂ�Є1=7c�Q�=Jf6=w����%=�jm���5-Y=�뜼��5�x�<�ɺ�N<=�e#=��W=f���'��i�(�6��#=U��<�+/�؇�K�����:���<� #�}uH�ٲ]<��=%�5=��<���G�U=���<��伤���7u=+�=N!=��"��;��y=���3��:(
？Ow��� =T\����(<pO�<��Q<��,<�
�b����~�G�<�K��x<�z;�p��^=�5��E��:9G=ޥ<iC�����;��W���2��6�;V=�F�Z�T�6��;oU�$��9��= L����kȁ<���X�<�vP=Whʻ����/^<�P�<2 ϼ,���&�c��%V+<�܀<n'=�~C=]�?��߼q�O��,��<��{��,!�eXF�����9N�T
�;�>[=@E�,�<�_<�6=�;P=�\W=Y�#�}��;�
<@#�����;Ht�UƼ)�f�y0=��&�dd�<��<�@���U=P�A<m�0<I�׽Z=��)��������(T�����p���� �D=�\̼ �м�Z�=�-�<9X�'�p<^�D=��=i��<5�=<�oV��y�;m+��g�<��=���"C<=��;��<w<�vY=��<r�!���`=T�D=����#=2�g=1�����<qt�8Z���>:=��f=��a=�+��%K���=��Q=g*H=�a�c�y<%�	�:��8>ˮ����XS=�T���=oI!��P=�=�;� �=)=�R���,��:G�eI����kSa=;p{��*<�=C=1[�<��<'�߼�����W<�2G��;
;x����U���r�N=.��<�����<֬�:~MM��4)=�g�<�q�\�<�G:=��<e��<+k�8�I��;w0=U�U=�)
���Q=V�[���A=X�������,=�A�;�=�<��9l�[;p����
= *e=2�q= eԻ�gH�\�s��޻�G�o��i5<ׁ�pXr<�>,<+�<=t�=LK�:�y���*;��H�ג��|<�U�����F1�¢�^]=��_��Q��f<C��<��>=�(T=�E=@-�9e5=���F���"�ܮ�<ߵ}=j���RP|=�=1�=�=�o,=+�E;{�<�L��߀;@�i�x"=*}=�p��/�]��3޻\r����c=�Q<Kb=M�9���<�5�;_�=��>=6�!��{=Д(=f�<$�@�^=X�����^-<�S��@�H�`导��-<�j/=:�����;����E?��c� =p��<��6�ğ��\:g�D�<LI[�V<�ٺ+�d�q�����;�7��n<=��I=�sJ=JS���	�A,1=�Z�<~�S�Rc�t2=���v=�=wQ��Zk-=�X�����D=�:�<Q�Y<�����P=7W=��㼽�}<�rt��S=U �<d�	��bC=m�<�p=��ȼ��-<���xl���x<R��;~l<6�)=�\D=��<�!0<:�#�چ~=U�`=l=]=��<�)�
�S�kXG=��=xS��\[ =��`�Ԇܻw�`=1��;lO.�]���!�=�4\�\�żO�M�|?C�Y/+<�;�j��g���=�Z��<�b�O��<�e���򕼐3�����yT=z��<����m=�l�<Ğ)�V�L=+�<�t���QH=�O��C��b�<��H=���4�<���<xX=}l-�ev%=F7���<�ԻJ�}�఼x�=����?м`v�;	ju;�^ȼB-9�щ �9���B=ڭ\����^Y�<'(�<d�$�j�<Y��<}�p=Lt$��&=�"s<Hd=�w^� ==��g=���:�c�l��8�:�t��L���d��Y�C=�0ڼ�5}<Kw*=x�J<ӽb��܊;o�9=o9e<�ǻ''1�ld�J�!<�^F��ֹ<[K8:�0����<����=�=ힼ�H����E=2��R1u:�m���R���e���N���?=�/��G�<�R=5��;6�<��X=>a��'��KSH=Ň.��Bx����}��<-_=�[=9�<e;n�M= �%�a�a=���<�]=X^��>���W�-����ɦ�M��;zU$�~q	�h:c�~���<u�<��g�hk==��"=�=����<	�(=w����M;�K�5�l����<�=��4=�f��d<�4Q=b�9=��;���N�`�"�@5=+��)��������>���_�fV����i[_�� �ԚƼo#�;!=���>��<��L=Z��<wrA��9d�]�ռ�P� ܼN?ϼR��<^G��'����:
 <�	�z�ݼ������;��?+=y�<&�E��f���C=�q=(���2�ސ	���;3������<�����2}���m�;A/J=m;^=M�����;�wT=�&@�oc=:<#=`�T= (����=���`bD����<����M����O��t���<yg��[������ܼ���:1����?���i�<;��m'�ڏ6��6�)=y�C(c;W�� �(���8��J=&qj��<>x�����1�=D<�g�e&
<,aA=��<.L[�}���"�<�Qd= ��<�?�t�F�w�ͼ�$�<�f)��J=ۭ1�`�Z=��^�\Y
���=�֢:�*I�U��F!�:�jɼ2c��C0���D�<�n��~��㧑�D��&����"N=���<~�=�<�C�9�=���=񲳺Հ=�8�\��w&�Fd����<��ͼ&yW=s�y����}m=����_=����ɛ<Vb�;ٌN=`�F��C}:�>E��	r<�<=�P2=�/<�h��e��<C���O�/'�<Z�D�d�,�i�	�$yf�,- ��ێ<xh�<���˭D=?-l<��=�;�'��7�<M��;O	H=�8N<ăH=��=���P�@�I���<���ʊ{�;�L��I�<���<R~Ҽ]4c=�>���/=�a=������a��F=%�Ƽ�*���S����K��KU��޶<�z�<�sw=�XY=��6=��V��ߵ�B3��<�ޤ<S:N��%ʼ&�z=����Y<�i漧�i�o=}��%�X>=S
5�QL���-=
��6��0l��(=}Q+=�C�<8r�;���4��<ԉ����<x�< vD=�i�<K���O'�9�70�?{ڼ=sN��-?�8 ��(8@=�K=ZoF��P^��ļ�L�7�G=� ;��u�;Fw=~��d�,�ꋊ��;��=S"��	F����9��#= ;��˵f;���� ���_�[M=��F=Ay���<�MƼ�XϹ��<��H��==��<9O�;�$=����\XP=�|0=.}�<r\�;��<){,���f<gP���e=F?,<KU3��F��L=<L�k��H����%��;Ŗ��F��:5�ͻ44z���=N��Ͱ=�/!E=/���f\�4l%=�x=�F<d)#=6�U��e�:4�؎ټ�4p=���<e�U=�^�;��q<W�{�<r:L=�q�C��=u��;�s<�-�?��t��˻�<� ��uD=NJ�<h�9=mጽ0��6��+�:uH=�	%�#\�<��<4�=ZU�<3�Z=�U�}�<�����[Ȼ$7�:'6^��W�Ly�;rVt<��=)H=�J<=���<��-�ݑ ���i��'�<8J�H>ۼr�=w_F;t�6��f���o/�Q@E=1����=ZQR�m��<x����n3=�����<���o&<'I:=�KI�BOC=�GüuU�;Ɉ#=PRb���s=����-\=PΒ;z�:�ѝ������vJ<�Լ�K=�{/���U=$7���Ǽ��i*��쓼�ɐ<�&'���<"�N��Լz1����/=I15=�G;sg�=��<x�̼���y���Z~�<uj�<,�M<qpV���U=�5̻iW=A���"��n�3�1y��	k��]�<��D���:��aټL��<>�f�<�ad���:%@=��]�qw���M=N���&���0@�a=��<�I��P1��}�<w�=�$�<7K=�xT=X\R=˘.=�$��of<Hx&=ϟ�<z�#�o�M��BƼsM���5���W�(d=���&��w.=�2(��E�;�m�<�2]�"=qԱ<��;.�3�%?=0n�� �=r��;c�/<r�x�+��^�3<y&]��˨<��I���S=i�/y/��>�<B�*<.N�</=��i�N��=���;�F��ʼ��]=]�;��<Oא<��<mj�;�d=���<�6`<o��b�R=+�����#)3�3�μ��F�~<��ż�P;ex6<�����O�...��Bd����;�t@��FI:�ag�KY=k@=���W`#=�L7=z/#�ڼ)j��e�=����_;C3=�w�</,�<����D,�"ԕ���	��n���9\�'���{<�^���������n=����<���<ѵ =��&��>�=1g�;5��7=[���ϵ��K�(= ���t
"=�=_���rg�9�=<$��<G3�B�I�� <�s��zn��]A�<�6=��
=��=V#�;��:j�z�q�0�W<�!~<�[R�_�����;�3=,.@��P=�p��|=�1�<�b=7˚:�������=��z�Eg���h�(M��=�]<h�/=�<<dx�ɇD=�4��==��
=+抽P-J��:<}�<��񼪰Y<]��<W=	�m���<�N�<X�޼dN���熏<R�<ݿ�3#�<b?�9[7�;.D�<���;�p==���k� =?�,��y	��S�<�% =.�E=[��<d�=��r=�E�3���M��1g�4�
<��G<�Dt=�������<��ż�g=AY�<wne����CR<9��<��f=E6+��)G=�'����<hߊ�o�q����<��<�#���-y���N���<>Ӟ��#,���ͼ��q:��Լ+x�����g�y�=<��<d�<��<���
���ϼ�:i�=-�.;𙀽 R<ӟ(���N<�S�d�+�?�^�@���1=fD==9��{V����<X��<��A=��-=�����~�<SP���<)�����<ad7�H�%^"=����?�=�~	=��R�C=����ah	��W|��ȁ��I���Vμ�<z�^�jv=�7��<@���NK=��*=H�E�\���nOB���<F/)��`V���<�B��+e�QNZ=�AQ=�<�-ּs�)�e��וp=h�$����<.l�<�4�9a��/�<�=`�<ު��S�G�N!8=	|g�y�=��!ͼ�RD�8&=aĻ�b<��+p<�3:<��\=�d��D�ڼ;�1��wx��B$=�����
=X�[=5K��5l����S��R/~���=D���B��f��]�����<��7�>�n�8�;}��<�P=Ω����;t����4<�<{
��ms�"��;�E��G=�>�<YC�<�I����<��E=A17<�fC=�UB=`O��[��׿��"=�U�<XE�;);R=�J�<��;̏p��T�!Z�;qT�uA��8.�o�#<R�=5�R=:G]<��Ѽ�MZ�����X���=�I#=hL�<��<*�ϼ=2h��+����<9�׼��c��Th��ն;�l��B߼G�ú������V�;Ch�=��=;9κ+� �	�;��7=�ؼ: Ѽ�Ȟ���x���=g�d=	1=��8�<CY �F}=D���d�<�2���-=1`�s��KW��}���$=��߼�ZD���6=�cI�w3r�%=s�#�8$/��W=h!�<7�\�������<jю�t������;�����5��،<#nZ<�1�<��W=�$;�'��O=;�����=eA������ټ{`һ�:����=�z<�X�B!�lA={�#<fO@=�� ��M=�`d=�2�9d�r������][�r?>��u;>M9��*%�O�%��%)=�;�#�Z�ۼuļG�_��́<�J���1=ሁ��Լ�n���+=���<����b�<�R=-�R�%��Ŗ��@A=�]�*�H��G�:�#��!|����<9�8�߄�Z�s�����=�&�<��<�2���;��y=����NS�0��<2x3=
����z��i-=�hT��x�<�=_��;��=y��<�.����<�ӕ�C�{=J�/�c�C�1`$=��¼\��d�����<"y�����<%c=�f�=������;��ۭ��"N�9e=��D���z�5+�:a����:�1v��.���^�q&<��|���	<[���r<��Y=������O^<O�
;��t�� ߼]_Լ���<B��<]=2�#������C=�X=�mp;�4?�����>�"<�K�<��<=���<
��(�;�w�<mN�;Ĭ=�Ը<�"��͓�$g<��O�^���$=Gy@=��D��Z��$/��Y=��
=ri���6���=��=N�<`4I�jR���'J<�5� ��g��<^#`���ϼ8��<& �:5��:k���ūa<����)t<%E<�a(�<��=�1�����Tn��ټ:@���D<~�n<Mn�m��;  ���
�l�<�Ċ<��R�>�����=d/:-/`=#��풀���<�j;t@/���������ܻ�d�;2�r��='='S=��\=�]��s=��]<�V�<f����F1<�� ���<G�*=`C=��=�u<vC+�2.<����GBa<r�Z=ҝF���B<�ZZ=yy��/}K=���;�1{��3U�X���F;;���<�ڼ3�<f��=�\<� >��wl=d=��<@�m=�n�h�<��=CW/��K=���<�[<�w=�<�[�<�ż���<������Z<0���ֻ4"r<oN{<�[�<�|^�yyk�?�ƼXR��y�<��I;Ĳk=�gr= �f�=B�*���+=�f�!�"�K�7��p��]�<b�s3���j�|q=
����� =�q�<�+=�id�їл��:ā=f�b�Om=�$F�)=�0�<�Q6;��޸;7�-=��;�$3=�f���ӻj�=�}�<Y$�<ynʻA�E�!�+���;����M=�p=NS���j=�:��-��������K��o\�Yq=��<l=�q��0j=~�=(�ż�|U<�ti=��<�ɘ<,s�<_�=��M=���<+�t��d�S�f=�j==�}��B�j��<sbX=��<����:F4=�*�</���\��$7�;���<g,Q=y/�6�V=��;���<i�ȼzeQ= ҂�\��v��Z�<����#�� ��<��=N�ڼ��s6�<�)�a�<8�<��<x�<b-�󄜼jՐ������/<,e*�Č���-���4K��%a���\����<q�c��H=�Ӽ�
<+��Bj�ٙڼdX��OTK�*>%=$�=��!�+(�;IA��=z�=G,�1	 =ve=�_<[�<ȀH���D=1��:>��<�$���м���<@b=F�.=AKf=QV
<�_軀
i=l*��p����9=V��K�<_C=F(&=�a��Ü��;���<�@�ག;����뼕?�;W%k<�q;܇�<H����a;���;<؝;%�Ƽ!m���ǻXW=e�Y<����`
��-Y=�#���T=ю����=V;�;�Sk��U�<q���@=k�ڼU[:=*ۅ=j0�<� �6�B��D��~�;=�������^=$=�z<��ܻn���<�<��=�]��.�<�Qb=��&=�ݼÚ4�W���=�X�<Nٹ@�p=�[��n#=�2=[�1���-<C�2�,v�<+�6�M�<�06��7�<�	ɼ۽�<�N�<|-ۻ3�|��=�<=E<�u��*�<���3�Y<��=�M=Fbg=2�������a<���;�����5�q,2=S)�<�=���� �c�^�]=c����<Swa��CQ=q�h=����H=g�</=�r���Y<QDB��yڼP�I=t���F��< ��<�W��YԻ�(���"=Z ʻe�+�q]_����<$���:=x3s<��p��&=M%L��&<�o�������ra=f��<��7<�S=Q�5�����<��<�g�<�`��C�}'`���D==����]=�x��Va=*=�hp}��o�v�n=�3,= I= �W��EI=R�u=k8�<�ߪ;(%�uzH���U�:��<ܞ=�4�:�v=@0<�@�<=1��;�l[���<�5�.|���]���ļ�d��	[=�^m�d㐼	g<<M��3�ظ<����V=C�^;�o=�b����<�C�y?=^6���༂|U���=8�?;�-����<�z���ps=�Ɏ<Dy�<5�#�z>=��
�`Ot�X<�j29�f�={7�;��Z���|=�4�<<3=Iw�<��@=/=���[��}���=>La�%:m����+n�;�*��iU�
�A�-k�;��A�4V&�}t<������-D<nj��=�=q��;E:=�h9��2���;���<���<L�-=�;мZ=�4V�!�����l=��B=ie,��L�;@T<�GR=�	=}!�oу=W�<�8<n�3=�s=�Y,�ݼ��>ȼ����M7�[�\=�;W�y�h�@�f�۽s<�Y̼��!���Z�{�<�1</A=ހ�<�[%;U��;"�l��Dy�)�`<E�*=�E�<s��<�#J��=��#�B=Ӛ;=c��St<�Y+=��9���{��J����Y=�"9<�;}�뼟c����A�o�ݼ.��v�r=X`L=��G=a4r<�(��¼�U3=P�7=3�����M=���J)=��;�X<�x�o�X=9���ck�g=�.���<� ��v!��p<�n�<�EI���'=!��*5K=~c7=��=�S�g42=�^���D���*<�V=�1�)̻<�����3�l��;�Œ�V=M�R=�N���.�:�s�~=��o���:�5X�x�=0�'<�Y2=�b<LI=�4>��yڼ.�i<Abn�q �Z><�&d=��=��=��d  �� 4��3u����;�
)=�{ =���<���;*��;z�f=��f�M=�vU=]D=j��|�=�q�<S���鬻�_�ZK\<�H��������<�M��!7<ɉ��4�=��<A�M=O8q���T#&�C�	=�|K=����Nx8=CQK=�`�<��C�jp"���?��3P�;�:��R1<�oj���;�A�<��U=l����y=hk�<��/�u�P<��;�J<�?�<���;P�.�Ї=G΍�LK��ܬ,�Տ=x�@�E;��;�^D=�
���.=�=Լo1�����;��<U3f���1��]<�0ػ�ぼaV=�=u��N\=1�%�DZr=��=�1=��ݼ
�_����}�</��;z�< !0;
��BK3�Ӕ�<B���g�<x��*Y���6=�3$-<@���z����(#=3�%=��<k�<�a=@����"��I�.��<z0�H[=)�5; �|�7� =A�=����ʼ��.�\<�"�<;^߼d�5�<�_=o,ּv�<>g=E�<�<���N}T=s�#=��,<�����5=��u<�T�i�S�&����/�����ݖ<���xZ3�&�o��=I^мs<��;��;�T<;�"=�H��64���_=Ya=hn�����6�^��)Q<�9�;.d��ڟ
<wDC=�5A��/�=���;�=:�P=>�����E�ܼ(O�<�Z7=C�P=I�S<���<�N;E����2U���x�BR�<-�<��(;&�i�s"=��ԼR��< S��ͼR'<����{,;��<X�=��<E3S=�?Q=��	��Sn=e�=z�9��߹��T�<�@	=[�0���,�8��<�=��e��φ�8b-�S�N=���<����K�݋';�/;�Wr��b�<::G<���F��=-8���<�@/=�>9=E�$�1�G�p�\=�"=�����*=��:�q��E�)=��2=A|;�j�<߼�={6-=8b=Y�N=Q�<!����E=���=�S�� =El�����<f�{�*�!=΢¼{6���<�^L=�aC=ᖘ�������׼)}���kw�v�8=�4�:ͼ���Լ�]x���=
+=�:=��g=�>����<�;�<2St�bK/���i�w񼤏�;��;y�<Tm��4v�<����g�<6�F<Ck��Q������:S\�5냼v�v=V�~�Gy���_=]��;oI�袸<��o���O�ʼM4�>�=\�8<^�7=c3��6���u5�_��:�l�=��U��Hr�I�e�5V=e��:��ȼM��<^��13�Я;�5������:�4�<H6����a=��	���<��<
��<�%<��v=H�E=0�T<˨�<��T�I�1��=���Ww%�E��_�<�d&<�5�<�e�<�Ǽ>�<:ˁ=	ʅ��iX<F�j�5��[�<�J���7=���A�P=,�s;�b��	�<x*!�cMw<s�<~�2=��3Q�KР:<&<=1g
�z,��=T_[�7	N�}��<MF9��L��ɼ��r�XJ	=G"$��w
�y� =e6�<9ޚ�_(n�c,!�� �^34��U�<�0Z=��8���6=]�R=��	>1=�6�f����=��
<��q��������<ػ�$�M��:5��q����;7=�O=ԷO�Έ�<�� �c
�<^�=?b=T�=#��<c����>�<]��a]=�F�;� � ����;OM[��).���m�<���<P�;�����V=Gb=�?k<��y���V��F��b#�^'���<o�/=�ܴ�5�;��<��;�}<�Pb�S+�<jNɼJ�Ӽf=^=�(=�a6<ΠK=�t=��h�h�_��r��=��a<�Ԁ�W��<a�"���^=�<P^�;1U=�1=�
��m�K��=��μq�=��!=D��<u��<Y=��i�"h�<��!<�D����;V.<��¼xg���HR=�L��o.3<�1-����</�󼵁�cM,=VT�<�Oi��`R��#�<Y'���C=5�:<g�f=�"Q=2T�<S�I=�x=ȉ����.<jA[��r<�.g�����'���y=rTL��~�<gB�<J��<�D�XO�;}u�H!�<�=�&=P����-���`8=��k��<�4�<��=��6=`��,�A=����e!=�DD=�{\=c�=�3=�M�1�?�Fż�<�G<i0.��t<��<�Z= �=���-W�f�k�,a�<�s�<O�<4"=Mn�;��=��[�xӃ�]�<<�/=�[���]�\�<��켈[X�펮� �j=i�8=֩�;�6E<]fͻ������0�����7{;T��<C�<aX��-=EO)�!�z��g��3��ƫ<F�!=4�"�Q�q�����\g�����%��<�<�AC=�|;�/Լb"p�v�<���xd��azq�d.ļ���<�Gv=�8�Ji�<R��<��;�k��,��:=,&����Z=,�e��M=�0���K���;D���%���*=j֣�g=���;m�N<���<ÿ���@=�8q��*��.D�+����j��򹹾�m���=���<a�м�\V=�:'����<�^���<l]}=��N� C��84�;�彼��<�]�VuV=ť=Sf��=�|O=L�<&~
=q�;-��m%/=��ż)��W���Sd=��Q=��(��љ�SP�<�n=�����<������Z=�)=uaû�X�mY�<`������W���I���=_o�xz���Y~;��y=�	4���#=e���>���u���w�X�=Y䪼�����#�0:�<�8����x<d�;<%w=�~[�<�-=uMH=��x=F�]=��<�Q��/�[���<T��<MS/��r�<�����<��`�@�O��;�ˡ<����5 =�+�3]=��cjR�)�c=[(a�؍�<��<���;\C�<����̀r����2kY�&� ����(0����<1��<}�B�������4<q�%<�f ��٣��G#�?�Q1=��h�ǅr=KT���s�:��;:Q5��l&=XD!��� <uI7�VT_�����<б<Ɍ��؀=�E���M�:��(�����;T=Z�һ�K��Ò�<Q%e=������Yr<�ߩ���h��i�=6�k�`%J�ǫ�T�B=�n=����[E�ˌ'��Mغ�N����r</=����g�N=��@=��=\����;j�:��o�<�U_<��e���W=V<���<Tjc��4`�)z����H�=z�?��q#�570��1!�D�E=�X ��b#=�������>��wL��䘼����������=+LW=���:D��=��a=x&+�<�J��J����d�<U�7=	cD���r<�\<r�x<�vS=�X�<g���Y{=ln�<�y������E�F�S�������ҡ2=1�<c(.=�o7= �*�2|軸?�<��<KeW<V���.j=|���FC=#	��n��~����q��<��Y=�2���<c,���;���`0�<�"��z;�Y��G.=��<�Q3;��ϻsM�;C�N��+�;�=�}=�2`=53g=�<H�=ތh��#"<d�!;O"�B�<���<x��<�2X=wƂ�S$N��Q:=3��:�T�<��=�������;}�����<���<8��;�&
��*}�d�;��o���Ԓ<�]�?��Z\_=}k�I�M<�<��S=Tn
�0�Ν��P�n�=F�-�W[�=:=Ram�UK8�� =�����)���<����T�*�9=����0p��|=d�D=�I;;K���Q5�<� =6�#=�g���fڼA�(=��<�v(�(8<�\�<�0Q��sI���<��_�n����=��ۼ �=!!f�� �=a�/=��H��>=�m�,r�:vt4=��w��G=}�Q���
�?��C2����<_�û��?�46=�t�<��d�kiw���K=�����:=�J=�r[�0s�-��<�%_=�lF��p��� B=�S==��@��<*:=q����^���<1u(=�]�<N6��<&��� �?�(�E'���<7�$������r$=�7I�%��<Ȧ|�W�<}f�<�Ia=gjH<ƾ���1g=�a=�<~��;Q:<�e�ui����<�h<��E<�< �?=���;�2�<- �hº<'�Ξ��3�������=Eͩ<��<�޺�D�<�F<ؿ<�j,��޼!�����8�:�]N�<��l�?(Y��f�[6޼B�D���<؛4=ϔƼ���N��<��"=}>�W�м���<>a�`a�O�C�<E���^=V�<���=�=���kL��U�<�ّ�[��<wy<�S=����W=�D�;AC��\77�(�ڼ��C���;c��:^��<���Z=yjK<hd�p�����=4ƫ�bMt=a�y�<�w���,��<�e���K�VC�J�1<eL\��N�C�$=|�=m��<*3<��"��h�_L=��m=�B��T�5=�W=���<�)�9�>���=5�0���+��eU�jP<�!=Qi=;��<G�"�ǒ�<����'�6i��XG<f�_;4�����_��vK;X�(�H�<��6=\)<8�V=P�<�͙�ۼ�GW=�H=�v�<g��<&T���(���?��‼D饻��%=b�s��y6=J�;��=ۆ)�wa�:� <�28r��<�^;���;Ϙt<�b���:;ѥۼor��2�=֤������F���=�� =�r���ͼ/= d9�r=���x�f�=p]�<���<��=�?�<�q=�
Ѽ��6;/b-�����ɭ<�l1=KF<��I�b&"�D4�n�� ���=_�=w٫��C(���<ڶD=�)
<��\�%��
�<�XZ�@����ǻ�CG=~\���<�V;�9B=葨< ߼�F0=�D�<���:`;[��<���<f_�<�|9�m;՘Q<�}3��&O=/���DP�ɑ-��@c�,�żl4�<�$*�MS=s�}��5��dR=nz��3HO=��<���<�-M��~E�.yc=�5Z=�<=[�d;"��<R(A=�������u=jQ=�2��C���2���o=��<{9�<���z�<��w7�=W�=%��>0ּ��Y�ӑ!=��ȼ�~�<��,<:��:��{9�����m��\���%Q=�(�#�=���<tM+=�r��R0_��.M=_e��̀<�0<��ۼ�>�G%X=�/�G�`=q���E=_p5=,�<7뷂<`��<���<��=�m�(=��F=dX4=�d
�0��=��#=�-��;�е�2���a�<����L���D��8 �K��)3��0��M��)c��kٻ�nM<�A;]�-=@$ܼ;k=��<F3Ѽ�O=�T��P�<;}�Tj�K~�>�m�ԅ�=͜��i��<�y �܎/=+��<A�crF=��(�3ͼ�DA���(=	4=?¿<Qƈ��6g�Uf�g���;9b; ��2w+��ET=S�,=���<���</�A��*߼�/��4�<
[�� ���;��=9�߼T��;�`��w	�7�<��ڼO&�~��<�Y=��r�G;�;#�<�޼�\�G><�<���G��P+=5�.<��5�'��;����%h�K�1�_};��8������<p����2<Fv=Q�/=���<Ʉ��@?��8�3�}=�+=�T;/�<�$��<v!X�	�<='�/=�,t<��;��2�H�K�բi�9�\��"=�%=i��4� �?���ϧ9���E���z<h�����<X+�<��<[�\��<�.=�dǻ�Gʼ�2^={������ʼ<�=��+=5M5=r����E��`���y<@�=p�;ξ��:e��;�h�ێ��ق:=8�@=��!��%l����;:�(�N�#=����>U=ٺ��</�_<�%�� =�>��Z=;W=��=z��<�
=S ~<ZL������y�e<!<`}T=U�4�h�r�'�B�w�=�J� ֺ	:�;�Od=2�2��=�k@��:=�B���,����<A��<�@�`�V;Z6=jM�f�)� �<+ԡ;-f׺��A=�<F�ʼ�1$=B��;�aμ�t���u�]�:��'r<A�$��`�'B=�X��j�=|������r��!N����<��nS�=ʥ=%[$�j=�q(�Wf���`�; ��T�Ƽ�8��Q���o*�@�<$�h=��멨<�ު��:���M=���<m J��^���V���1�)4�ѡ<��P=��6<c���=&=&��!ۆ���S�8=I��=9s3�hr���(��P=�M�x�I�4�f=L�����D:Ec`�
4�<I�<7��:�1Y�ZS=H�}=m�v=�%�$��<�NB=K=�����&=m�L�(�>=S���P<PY#=4[�<q��&/P=T��8ҼG�>=#j�=��B=�:=-�μ7���/=�+�W� ��<+o�;d�*=�����A�����ϣ�<A���]��f����ň:7��<�:Ǽ���<K�.��S�����	�!=���;��<��-��L:���<�*��w����;��0��3.<vs��Q-�?-�<����*e���x<u��<��=��K=|P=�W��up�Ζ���<+� �bV��sK�'/@�&/�<�q���<�Ho����;4��<PG=�a;=�t=�Ż<ۛǻ;�Ƙ��L�7��c =|���q<�g=�[������b���=6��<\�e�`=�ɼd?=�]k=�?+=~�2�qc"=�˱��r<��0=U��<��F���������g��?N���V_=�>��y<=��м����C���#���<��$=�q�ƴu���M�u ~��@=`��#_f�>ij=A���#�=�"(��</�8��<��z<0���;��rs���y��+H�� _=�㶼�@(��Sg<���A�l=J
=F�K��	<��=��:
�4�E�<\=��:=}n�{�<y+��(=���:�4=j�<t�
��9=_ߣ�ew&���9ě�U �����( =����z</V2��oO=AC�*eS=�u7<�l�<b�ż���<��Q=�{�@S#=�C�:�*K��:�m`@��ul�i��<���<5Xo=���LO}�#���W@ <i>=�L�<��&�G�T����*��ӡ��t�T=�<��4=uf�<��<��m���C=SOI��k�<��/�#
=_hk<T~��R�8==$`�i��V�;�t������ ��� ="b)��J߼�d<!�c����q#���-�}�Ǽ��(�jr�:�\M=�ʾ<�?.�%^�<2̏<m�<�μ�U��r2=�
L=ju�b��<�P�B�=Ek�<l�L=�!<MG�:W�,k(<b�I�w�=�Vλ�]�!a�p�=�8T������RH�O0���/�?x�<���]�<�b����<���;wU=����'��X<��=��S=�Q=p9=`EJ��U|��	=ô)��I=�����tg=3>=VP��ށ9�:��[��� ���y�K�^=L������~����5�6�=]��<ys��*�t�<{���x1�m�{��qt=�1�;N9�<�s=�Ե��NE=��iJ���G<��k�l<�X���Ǽ��>�86=�n	=5rg<�i����'< �d<)�9K �:b�;VV=�Y=֖����;�!�T2�<3<����BѼ�Ue='�\��~U=��I=qn���	=�٭=3����Z�3����[���������<caN��Cu�a�=H=x�����ռ��@�'q=�e:���Ȕ ����=�!�CE�<�?�<�<a�;=�.=������}_=;Ƽ��R��D$=���G����<��Z�#�+�{�	�fG=�|=+p2�D �<�� =C�;��Ϧ��9D=��.)
=��=��:���<��<=�v3��`=I:��aUw=p*X��v�<���������s=��7<ق+<~Y�����%94�>l=PxE��<�+�<���i��<i$=�ѿ���5<}�7=]�:����E=��L�U�<�<N����<fU���)=3���Q	<��=��F�%�<���ʼ9D��|�<��'wM��G=}	g=70	<��;P9�)��<�J=;�<;��F=ߘ���O=r��<���Ƞ���<>(�Jżʾ����<m[~=^q�V��<B6<�++���%�aؽ���<��<���s�;`A;mp����:�G��1x<�K��䘼F�q=e��<w�p��ɹ�K�M�`��]��H.==9=�
K<a�v��M��C	=u��<�V=B�Q<�mg�_�`���޼�F��
�=���v�_��!ݼ8�,=E���,���~��y�<�}A�d-w��dF���<(�J�o�"=�
=�%=����������<my���Á<Y`���q.=,=�}=�ʔ����or<=�I�:�����ӈ����^�(A���2�R���X��j</Ɲ��*�<�<'^�<�ŕ<9>(<i��<-�=�(��2^��;��o���0��~1��I<}@�<R��<%�S.ʼ��:,�̻];tC ���WB��@�<�ٺOO�ajo=��L�N�=/�c��H@�:`<<��=�/�<�=�>=�x<�>=����|?]=����$�p��Bh�r����	̼��O�@��<J�ɼ���1^?��k�<<���Ҋ���Z=�q���3�y; <�g��=BA��@,׼�09���\��bz<����	��gj�H���#����w�<n��9.&=�&d�܇��3ı��iH�+��9�=�3{��6�<�~���"=N�M=��=�f�[iP�E]��0i��X��^D<�D\=��<"�6=P�{=�\.�������<�����C�H
?=�{y<�@�l��=R�@/<�'B=�.�����&g�o ��>��V�=���%�:2>S�`0�=Aʐ�d <�pq������;s���j� a�=<��<�6Y=���<�⇼y�=Y$ؼ�[)�J��mμ�`-����b�U��S<E���:=�������<�>�\�����;D	�<��@=�U�S2��!����<E���^��E=��X���]=E�=��;�����2O!�P�<�������<�s�<�$6�б�<��<�9;�<��d�)-=��u�a�������h���D�9>=n�7<ݘY�'.�r(<��<<<�<m�4��b�<��<8�<k�=���C���L<��>=v��9o�j����;Յ���=��=�N����L��=K�P�@=��3=�b�Np�x\T�$�6=y�6����̯�<ɐ� +�����7����1�G��τ�D�=�<=P�M=Z�O=4�G=+N;ا�<C�~�� �=��{<d#t<4�=�����<��=4U��D<��C;�G�<�G��`=�R0=$EA��e�< F����:>_-=S=�_{=�S���=1�t��
u��C<��<�*�_Km���x=���  ��RP<a���7�#<��c=If9;GA#=ݜ�<ǂ�澂<�jd;u=���;���i�=Z�<��kC;йl<>~.<NW'=���<�6;�_�������<�D��f�V�8<⳻ny�~��<�2�5���6�7p�;P����=E)X���ػ�<��%=��6�<A�<�������#a�dC�q�=�����;���<�̷�מ�Fė<���<�=�j�<�d��~1����;���<��=h�λ��<yTA=��<��@=<�����%I<�1=̊^=:7=�q�<s�缟�$;��<�v�<���<4)=uJ7�`w]����<�<�s��˫\<�
2�j�q�0��b���L��^����<͑6��M=󅼂n�<Ű=k�L="�2���<�9=����Zu����=�)=G�м�{<I����G�<,�=�6P��H��w/<��!���p=����#v�{���,X�<6	�<ǌ��ړ��=t�=�'{<LiC<wpF=���þ�:�2=�p�<P��<���<i_�<�<�+/�p�=Ҟ�<�	K�4�s=[�H�fo�<b�3=�=w\r<c�7�DL��p�������u�<b_=Sձ�0�A=� J=�U��k��+���덼�釽�y�nQ��K��5#�
8L< ^u�,��<kK�V��<!6��D'��c�'=:.�<⅃�)��<�P8=�<=��`�/�n=H�=���#���t�H���o֥���<��<nꏼ�D�<Ǘ�<`T@=}�s=up���#=#�;����vjM�s�����>lüc1�;�f;���<��	=Y�z!=p��<���/K=�$�<q\��n��k��;�(�)ѫ<$�<�8E��/n=&� �O<�i=��y��Q�Z�>;�P]=�,�uќ;�w��F�< ��<��<*I<n��<�����:=�-��=�������
�r�m��<~X =�w��T�=�e<5�<=w�4�;D�<v�=$��λǻ�7bL�0�|�ţ⼮z*���qU)=��m�v��;�<�;>�	�&4=��u�q3=��,�H0�lQ�t�i�YTT=�|��<��9=��;��;����:���[�m��=,��<�*;�nL�!�=�+����'=ꃄ�B���uF=�kw�j��<���4*C;m?,�`�<rj�;O���-zS=�x޼��.��Q�	=�D� �S��v2:Aat��/1=_�<ؼ�<�<o<h�c��ؼ/�����
�󜣼tl<�^��;}�A<��B�D�<  ������2��<"ټc�<��<&��<\+���D�۬#�}w!��׼|����>��ň�i۔�p�k;j.�;��<��?������ǋ�J��pl�W=���1�<"ռ�+;���L;�R��1�<�<L�z��<y�=�jGB���Z=�7G�R"x��E*<��3��eX<=�lC��煼P�&��g;�ZC�yEü�n��0.���6�֮O�GB:��I��)=R W����<�~I�?�=����;O�w���a��dܻF��|bC=jk=�w�;�V�؀�k��<ߠ<����<d�;=(r����#����w�=$�A�� <��"�!f�;�Y8�eR#���E�0�~;K�ּ,މ�":��)?=���{W|=C�N=�a�<�h&�D�d=j�K�,2�F�7=3�˼�}1�p�j��-<���:��,=9V�%�=.DƼ̲����X=�0f<�Q���m=��<�<���߻�4�C=	�b�;x�m2�<J�<-U���7����<Ľ����� ��;<�f=��H= ����7�Q�R=��Ӽ�h��:�;5+���_���t��O=�^=�$G����<��<����C=�A������<�!	=�
�<)sp����yɣ�0=�o�<�E�D�:�J�<b�����0��^<q��<,5�<)=o��^3=odc=�=��p�̓=}!���K=K�M�",��K=0�7����m�<R�z=�v=�6�;�K<WyB=;���$��<-x:�C�� _=Ҥ�к#� �=��<J�l=Z���D�Ļ�>��V�)��[�Ɇ;W���2mv�a�<;�<r1�G�?�����M���Y�
��k<72ܻ�Av����<��<݀Q=q.<� ��ZR=���Ā=!�A=p/�<�p���=t���M)� 6=��}=��=���<\�`��Kj=@�m<�7�OL��a�NO�;1�[�Ԭ =Y�	=������/~.����<(����	=-��<�=�,=ϙn�ѫ��JX�
]��&�<v�Լ��˼g�<��\=���b<ѬY���F��x8�37i=�t=��<��b��%;=�[r�Ɣ�;�~=���F�'��E=����n=b�?<=��!���V���0=D�&��S�,=5��Z�^;߲¼�l&;�5��~�<�F<�--=+#P<��!�{<j��<���->?��K���<Ί=)	.=ե<��<^@������<yZ49�?$==�E=XZ�����=]m��ͬ�R=9Z�<��n�a�E�9}�;֥���z�<�i?�g�0=�k�<�QP=�q;=4���P�;�=Gw�<�b���H=�<�����������[<)��z�D=�O�� �P!S=��&="�N=�	&=f0���Wм�jV=���d�=V�=LlL<^��</�+����<[��	`���i=�2 ����wȐ��ma�I�6=u�|�	�4=��ͼ>�X��;H��<U�K=�E �J�d��<	�=�
.<��<��k���7=�=C��o7��U���g=<b=-7k<��$;.�<=MK!<J#Լaͺ���b��+�<�F=��̼�'=i�
<��<֠,<��I���'�i��bv�:_g<��.=�"M���!<�3�q!�<��m�e1�v�5�^�[=<S<Dw�X����<T�<<^
<���8�=������:~�<�#W�o�ڻ>��<6���1�<��F�ĭ<�K�6�4=B6=�3�����fʼA�y�K��;�N�<
�.=�_4�)��-}=)���P1=g�5=��`�H��(bS=�9(���q=�q=��~��k��5Ơ�K���uP�r���P�Y�cj=�};�K��N��]=i8)���Ǽ��i<�j�� �<	�O=���<�����V&<̀K=�A��S�8��!=��1������<2�%���=����2�<�&=/rS��7;<��ἳ�g�T$��Ӌl=&�%�dY=�i)���I���<��L���9�Ob��H���(=�|��"l9|������<�K~=k����=蘼(�������M=��K=���<Ю&=��'=��!���p��s�<Y�=��1��@<����=z�b�<�Q���=0�=�S���;��{X=iTu=��
="�[����<:� ���=�\��<���8_��=�$�92��G\�c�D�^i9=�d�J�9�/Id��%=�z<��n�a�<S0=.R=��<D�!��<�ٴ<�v�;=!��[�;��\��R=(��<��s������<P(�-�O=D�3=�3>=�1��8�K�i;&�6���5=e[=I4�t!o�ܭq<'X:����)e=F�^=49�9�@ܼ_Z�=o;@=�5#=������<d' �c��<rռ��.;|Y`�|{�~3�o�v=o�����'2s;<M=wj<�ټ��D�O�<=-V$=0 *���˼3# =мq;)�(��wV��I���U�Th���@n=�Nf��"2=���T[h<��;@Q�d2=�m�.*=�Rv�$�y<��Ļ:�Z=�A<]p^=5$R=���;Ub���<o<=��2�A��׼g%���(�~���ke<gm&=��<UW=�=�m;�ǅ=��<ܵf�`~�:�ӂ�\��9�F��+e=����վ�W����6;=:=�<'aq���^=�.<�< ^5<�g��9=���<�����0�@�h�~��<o�A;��=c&/=h�D�	9/�~Pm=�ỷ��;=�λ-pA��	�qg^�$��<8L��.1=�<������/=�^�<�����[<��<�h��RN�@͝<66=URм�J�<�[��<���9�l<�YY9=���<I0�]��Y��� ��;��A��gɼ��{='�4�DV =+Pi�$gK=J�����cּ_��<�J<����a�<2	=sٳ;}P��U�ȼ��M=���<��V<�Hu��Ʌ=#\�<�r�;Mo=�}<�a�;���<3��<���6�<|A�;M�@��yS=ތX�]K�<r�ϻ��_�)��<��j��K?�<`v,�oӻԎ�<쎩<&��T��K�5���D=7] <��=2 <�Eb� �!�l�=D�<ھ"�&	���+<&�9���=�>�;LY���E�%8м7�V<O.�<x5=YZ�eA=���<,o����<{�)�����;��;N=K;LӶ<R�ۼ6�e"=%�M=9�ܼ�f���8�<h�=T�;�7�<@����t=�����M�ct(=�b�;X�=��K=��м��5=M=J�A��4<�)=��Q< ��<f��<`��;S'K���E�x	����`����<��7sO��"=+5^��=�O�e�"�\u9��jǼ.��<�#�<��LI�<�k���&<f��;��=6R.���h =�/:�n����@=W��4�{=_��$r�����;n��菼D�C���0���K���=}�W	t�{I=��;7E^=���=�ۼH1W=��ȼk���2=.f�秩��=�B�#K����g=p�rFn��|r<R��<�a��l�˻nc�=�Ξ<+�w�6�$��k���~�9�8=��G=Z��!�~;r�:�<��;��Ѻ�X�@�=",�<��	=��<9�D�u�u����<:jҼ<����<��x=�k�=� ;�l<�}p=����:ѻtg<��a=�<pi��Q�����ռl,=k�9=I�b�ђ.=�w@��+=�N��K��/=a =~�V=a=�}�%ͼ�w��u�<\�M���[=�?"=c l<{�'��n�<��T<��E<�;3=A����6=���<[��hP����ټ%�Y�)�=41� ���B�w=�L"����;�S ��������-�'=u'"=*S#�(�<c|r��ܼ��;��C=��=��><�ݼ0�\��7�;|<-�Ij9;��;��∼_�0=�*�J�G<�ǁ;Xü��(�z�@<>��S�<�L)���"=��鼇N4�H��^�C=U^`=>�?*9�[�<�6�<�G���4���u*��O=��8�������غW�=���/'��G�<�&����L�
�<����=A=(5=�W��:��P�wr[��!�<��/�N(s�;6�<���<���{b���;��]��м��5�lq=Lkۻ������eI_<s�Y��3�<��H���f�N��<�D��)�
'��C
�݋����v<�2�<�i<#඼��=+��XK?<Fz��J��<�����2�:�<e=laǻ?Y��.K����\�=;Uv�]�|=`����N��6=��F�==n�\=)\˻w=�fZ��:��Ӎ&=挆<��W<:�=�x��?�!�&P컲i���j;g���<���<�V<�ʄ<�.<v�I����;��[cC=��W���)���3�S)&�̵�<;�׼2_/=J��<�*�:�Z�zY�<8{��ce=|��ŉ�8켣�L=켇���?�f��<r`]��/��$'�:�ּ�o���F=��9<֩D; 6d���q<��F��@ ;�߼�Hf��L������+=L_=�m�<��%��f�</il=�G�%Ԍ��AL=��B<��P=a�����v=j��;�����;=7Hû2�=�!��O#��zA=̵<�>�SA<�������z=��k=b
@=z�=s::<H������k{*<O�;�)S���ڼ��h<�H���j=7�8�۲F���<�B��Z�B6=̝2�`�4=,ׄ<��<�d�<k1=��e���<O��<i��e�<	>���ļN��rԢ�-ú�'l��>Z�K\&<�<J���<��ؼ��6��~��
�2�e�D=���<���P|q��=��t<�1���A=�c={`���^>�\��:�f=a�8���K<[F �v�"��<�m��	9�<0���W�!=�Ԉ;�����:�vhj<��7<7�L�	K��82��)�=4�.�&���o��<oȲ���<=t��:�`����I�KX=�w5=�o���s,=�x���<����/(b�u�a=��f�'���Y=d�=�h�<||�<�A�<Q �WrD�Yr��8=U��<�4w=�=V�-:��<.=%�u����<�86=�-'=(t�;Cz��U�ի��;.輼E=��i=���<��<���A�}=�����=��!=��w���;���<��'=YVs<�u��ޖ��Ş8=��B={V��y4=�v=�C<hg9=�`�<�9�<h�Je<��=QN=��<��F��;=�Q&��l��{�������M<��?%�M����Ȅ<r��<n�軻�l��a=b�V��3��9�%X�$�������}	< <��`���N=�ؼ��p��	=�%"=��<vC;��sɼ���<�O��D[=l��W�<�i�:�\=�r"=���<)��<Gm�iV�<�@\=\;7=�D���<�Y�<�:5��gL<���<~]<a�/����<�D�<�5���<��<-����M�e=���<EA�<-�,��2ļm�H=:>�<�X=*臽A����V�<BU=(~��;���-=>�Q�,�$=��~���Y�`5G����:�<,�¼�7��{+=Н�<t��<��I�q�M��\=�&=�,�<w�$��nI�u�G<��¼r�u=�`#�lռ{o�A�;.�b=s����k�<��=f���[3��͟ =�ng<f��!���J�N=�+ <yD��T7=�%H=y��<��my�;�+�<�!�_)p�����P�����=��<���<�!@��h��χ
���y�jX#�-[$=:`=�(�=�b
=v�&�%I��7�&��Ax����<���<D`���k�:ЉO<#OI=9��<!��0�0#d=�{@�yZ���H=�R��<�o=��E���E��f*=H����;�C6=�}�5V)�+a�<K&0� .9=�S<D�~�-�u<�鄻`O��¦�������;gO�=�I��a�ܣU�@�:��d��r�2��:Mn$��B�0<E�%�(�b=w09�Q}S=�r�=v��EP�<�������[��<��<���:�&��J���-<�d=T9G���<xSƼe:A�-#���=�R�}|m��M��أ�:̼q�Ӽ럖���z=�ƼW��R>�a1=�<=mvL=ƶL<�W<B2���M?��\�<)o�L�=��?=�3!�ſ ����a�@� z�<{���{7�x>�<�\g�A�E�T�t|����E��2=P��]�<,)3=��V=��)<Ұ~;�%<���<���?�<���:֓����6=U3<�P�q���;���<!S=�m�>�V�����o�� �	�M5��h����b=EB3=[l<JvO�3*��<3�<��r=����9�.�W=;��;�?�1�I=Q�;K��;8�==��4=���<H|,�p�\�B9���:-9���M���:�|8��T���l�|����}�<�^=��#�*�x�&=h!H�sb�;7	�<i��=mh&=F��<�M~�Ӣ=����/=�#=�C)�n;/=�=�;�D��=�!�
֕���޺YK�<�=<z�:w����<bT=P�<���o�I=8Ҋ<�(%�h<=�0�y|=�Q=z�J�y<b;���<d��<	��<��E��r*��hֻũN=��d�N$=�6�<��l~D�������;f��$�<�C;
��V,��)��1L=�(.=n�;=�~l���J��P�<^����j<$s�<V}v�C!=Y�|<$�b<�&�<6�`<�O����;�K�c�+���N=Dć<꾼�0f����������t�<
��<�\�^����3�M���A���z�)gs�]R»��D����F!���%9=?�a����:%2�=�1\=����E��(�4<L�^���<?<��<{�*�M��<�%��e'=5�5<;�ڼ|uU=N�;���I�;�؏<V��;�ħ<���<.����J\��~��<�lS��~�<��{<�+X��WY=B�`=��g��#=~�ʼ�JT�tI���	4=��q=��=&�-�'_�:vH���9�m�8�`-�<\��.Ɵ<�--���=�$	<�=�UB�0�� <��=F~�1G�=�q�+�)�� =�˰<�,�	�F;#wG==��%�=���� =2~��`�<��Y<�U=u!»�R*�F�N�11=%x=�%��m*=})d<�
@<.cż�0=%֖���<P	V��`�e��<����/V��_
<�i_<Y��Fad�-t<Ϝ�<i�"=����&��<��JN<��;=���?�ج�r�:�)*�7��<H�<1��<X{<x6�Q�?=��&��;=c#��y.M��݂<Ky<�PD��tH�v�!�C]�<��+�5v2<֘��*=[������/'=���}�*�R�U=85z�@m2=�lS��C���� �� l�j\�Ʒ\���<'�R=�d!��܆;��R�+|<���vh��E2��=0<=Oá��Pq<�1=s ���<v����輥==�E6�P=�C��I:�<� �M+�<��-�� A�_-p�gN�;7�;3�[��P�K�s=Z�>���<��
�=O<lµ���ܼE;j�J�M�g�=�>&=�$���/�=d�Ҽ���<8��+,������^����"=1�;`�<���޼��Y�&��=�*����p��
E=��*���N=�|,�=�[���˼���q�ͼ�D�<>������>��`<$b�?zP��a:=If	��s���G�:��i�;.�< Om��=X��<)r�|oݼ���;�I?<��]<	�M���p��[1=�N�f�v��wd=m�=�ZrƼv;��u�׀��|=�����ƅ�?�輿>6���<�a�U�T�>�;~�A<�;=&=�6^=)�Y=��ۼ�J���=;��<����Z<�������:�r���r�6c=�p)=�k6��.��$�[��tS������8&<ª㼢=�� ���B=.�<(	����=�y^i;ǘ�;�	���=3qϻ6~�=��<���<�s`<�G=\nd<��T=��<FF=,ʑ; �3���=��5�>�t����5I=�#�=��=�s=��v�I#��(��=�҇��x����G���3;8��<�}n=F�?<��F=���<<�:b[s<�f���< ���D��@٥<&΢;`�
=;_���8t��S}����;��������z�;�[=ω]=A�!<�x=��=��=�3=w��b�V=�'=ݳ~�&��<f��=J=�ϙ��hx<U��NI=Ƃͻ��?��O��O3�фJ���
=Kt�`�)=6G <;$�q�t��_D�V3P:��'=�MV��c�;3��<��t;�z:=It�q��;9�ւ;.��<�8ԼЉs=n-=f�I��h�����t=�:=�`ݼ������;ĻV=��t=2�9�I#<��,=٘@����g����q�Ƕ[<�X�����;Rf>�\��n���� �UR�<�|���~��~c=�7�<�\�:��h�������ջ��ɼC�ͼ��̼;�����P���̼�����|��*�+��"����==s��<pz=�O]<?8��p&=�bD�\׻	=;9�~r�(cʼƪG�ި����;�k<��l���<��;5��=ǟ�<!�F��=�ļ�WK��� ������<{�,=������;u�:=��J=�;)K(=�*&=��3=<'K<� =��B;18��#�=ӂ=�=�Tm�\�M=k����=)m���.=N�"r����=��<��'=���<
�=�P�żx��*=�E���3�W==u���[a6��;K=�9�<�A���ռ��L�~�,�V|0<*ԍ;�,�;Y:�1-���ɼ��(=%ᔽ�ٲ<�(^;�1�0b=9�U=n�i=��m=��<\����<��ٺ�a�N�=Ӄ<9�J=m?q<kd���Ө�f�<�B;)9��4�����c<�K�su����r��(����D����&=�l�;@�L=��}�]���b�?:��</�7�N>�S=@#��=��Ҽ.�A=�������z�Q<N[%;�����:=}�<=)�?��u�<f༬��<�?��=��A"�O�׼����<�Yຈ|u=)`I�@9�NG�<e4G�?�:I"%=���=�Q_<�C,� �I;v�6=��4<�>1��Q=+��9�=�8=I5��|-=�x���c=\)=�u=��6=�ȼłu���=����;�I[�_͉�<�;�Q��.Ҽ���<��ҭ�<y�=R����=��U=�74�k�j�CQ�(|=qg=T�=͙��� �YU�<2rF=��;@�;=�ͪ<��T=]	�;ŔN����q�=I��Y�^;7r*:���<W�<]8�^k=��m�t�A�|��<bE��B�/8�<��<�i޼$U=Nz��lü���;~X�<������<q4@�պm=��=K"K�[�.�`+�Ӥ�<��{�aZϼ��,��X�v�W���h�y�����v��梼%�%�9�x=�<6=�������g�贽;4�2��uN=в׻WV׼�G<F74�Ă�<��k<Ķ�<���<Ʋ�<pN�<`�;��e�u4=l�p�#�4;�g�;���L�R=�z=��<B�<2G�<��h=�n%=�O�6=���<��h�=�t�<��<�$=��P��^λ�6�<�񃽦����V<Y���5�W=�z�<'n�D��;��X��������m�S��l�S<y��!�,<AC<�p=7�ռ����~�e�����A�<rq�;�`��f=��e��4���)<�K�U�����<�ϼ~9:�:xἧ�:���N:w�>=Ě�2	=n��<2��h�ü��B=jU�<@�a=��"=P�V��BC<���;ʨ-=�i�<8�c�[�<˚ =�`ݼ�N��ΑD=s�p=�RT�o�	�� �=}+����<>9�( ~<�;�k:=�|?=���xlѼ/���cN<&��9hS<P:=B�b<u>���Լ��V��Kʼ �����<�J=�4=��(<M��<Oӿ<�`�FM�<��=�F=�_���!=çl=R�O����<j=<=�sʼڛe=xa�QVy���N�PO�Pƭ<S�$-<l������/�-=������z���X�;ʆE��X��w/;�y*='�#��jV=�u�1J�%�=]�=�b=I����"=
�Z��KF�Jb!=�M���%=�R�E<�����%=��=����P_=�	�;��;<h���hc�<��=��_��j4�r"<C#�AS;�
JǼ�J�;� =��5=����L���=s(f�(�(���f=��<����Fn��&��B�A�^�h<��:��9<�P���<%F��7v�:���<�D� ��=��<���;Ѵ�Z�?��m�=��=��<<��<��P�V+	��ck=26�<�K�;)=Q���7=��Z=f}/=���� =<�=��-�n�w;I2����9X7��I=��+��?�n�u=z1�9g�P�����ZӼ-�Ƽ��)��)��t2=4=������<�/=[k�v�N=4
z=�>=��P<{�Ѽ�.���������<,?�%�<����;� $�<�P=R �8�E<U��=�u�����<�}�Z�<c��;�"f<�H=*�H�h�ƨC� ,<#_�<5�x�$�S��Y?�J�����P�<*+6��;��< �s=�qq<[w`�\���*���uf=-[�+�N<^/�<���<P��f�3<�k��q��˕�tF�ޘżx�a��(������r,�E�P=�����y<e�-=w⦼��ٺ�k�� ��<�T�<;),=T_�<��%��h�v�漘�U�'Da��v��?��j=��&��ڽ<���`���2����a;���;Fv=DѨ����������<��p��H=@i<�L<��5t���L!��K=��o��\\�l�^�G�(=FF@=zM�;��b=�"@=R
_���7={����@���H�$��<JV���m/:�<�7��#=�-=Z��;�F<��X���=^�����ü��L��.��oL=gGZ=P3i=s��4�<h�p��և<��<ޤ�<�
�<tee=N2�]�>�֊%=�߭�%(���R�<��=�6���vW�3�a=b?b=��ּAs�<��?=�[�<:
<�w�l�C;��a<j�f��x=9�H=3ͼ��긬�*��D=�$=��R=��¼�=���1[�<�6=ۗ@<�<=���<��	=L�ź��}�p��j� �<��=g���1��<��<lw�<��-��!����:��:<�˼�|<u���k49=��=�c9���k=ڿH���`��	�p[/��uH=+�뼜D�<���?�
���$���E=�:��,���4�1��@I�<�[.=�F=7�鼢�6�cR=���u0S=3�j=E����V=�<�}�k�0=�V��3�h �<E��<pk�<��g=��q=4�ڼJ�Ǽ<Y[=��;��#=�:	=/�0�������&=������<y��6<s�>�d��<�<c=P�ջt�<3<=���<F�����)���<��`ҡ<n��<�3��?�}=��<����L=�H�<zn�<Z�R���N�U0�0�<��=�q����w��sI��D�n&=�'��
�1��Si<�ӊ���H�����D�;<�a�D�<h_�<�BR=~�������@=���o<V]{�ǨE=vz���`��_���;ɼ���<25.=9��CX==�n��7<.^>�xo�<��#=�<��Z=%S�^s[��һ�����L��a�;")���=DI�<6���TH�N�*����<�Eļ6=�<s=���kYռ�@5=)�H�@���X�<�=ɷ�<6�Z=�]=����n=3=�O����b�<���<EsO��ѵ<0�e�]s*<T.�<(물l�<��,���G��2��d	��s�<^����"=�0;̭+�m(�:��=?�J=�2�<�����+=ľA=�,ʼ�!=v�߼��<�4�v��K�<��2���"����3@��v�мz��<��2���P=R�'��f&�Y|j<<��ڞ�=������ݼr��<A@R=#?@���<-eQ��#e=[�|=<]W���=��qX�7������)�#�<(�J�f#;�:�=9�5��x����<=w��b8���7��i:��~/=��R��N���Ԇ<����9 �?�M=#~ =��-�8��4]�Y/���7<"�=� y���
=�-�<�i�<A= �W=�XӼ.p�~������"f�:���<���9<����y�%*0�`2=�O)<S�O=�dg=��~��`�߽��jDq<c#�R鎼�e�<��Z
��B�<�= �=S��;�R�;��̼�C��r-<k�9<��<��/�ڤi=���;�|��`-��=�MK=�����43=hQܻ�_<+��༰�E���<{�B<��=�fK;,��<���;��=$b,=�Q��[�6=�%�Zy�<�<S���G�U=Z�"Jc=�	�ɞI�+B9<`?����%=�+�<_��;[�<��X�QV�<��=�Lh=*!�<��`<�ǡ:E�a=o�F��&P�v4���_�u����\B=5qܻ6S�����Jq���ć<H������n(���*;�P=�Eq=�;H=��ؼ����6 =_�'�P2ջSD[=�J߼p5x���qU+=T�|��FR=�+4<	J�<�����5=�X�;��׼%ͼ;A�<��a�Gy.�Nؼ��=h꿼Fk,=��!=b�[=	�<�jr�ֻ*�Pv:=����C��!&=Td�<�~T��a�_˼�a�<�$4��0��!�<���=|ҙ<��;<�C�q�i<�7�<֨K�ٽ&���>;���^�;=�+=q*<�<v��й,����<iRb���;��}=���ɛ[<(����\��8��GԻ����K�W1�<�rJ���G=W�=��=Ŝ��7T����;�-�˼%�<<���	?0�(��;�f!<�J�<����i	<N @=�N�p������O�<��f�é=K9�<O����
�pn/=z���%-=�E=[�o���<wW��U�;h��<螙<�xW=�'=��V��ZE�j�<�H�<�v����;_nt<�7J=�=��9�=A��;�0Ѽjw��g̍�7���>T�9�мc�O<��D=�sM�InH=��)�f��<�	J=�E�<=ƭ�=O��k�<����S=%
����zi�; �?�U��;�/���)�����;��y<s�;�<M5�t������u%<��<G�k���=h����=#���0��<�5�<�i=��H<IvT=��G=h��yԠ<6�D�C��J5=p��%t�L4^��qh=�c�P�$=�r:=�+i=�M�<�N=�p�<����\����<y_=8=����;�$=Q�j��{ż�dʼ?�<=&~|��ɼ�q��Q��<��[=^\_���8<<��<�L;��< �j=b��<�kS����;���<���Τ���W=4��MZ=\����<�hO=MV �|g����<�s=�s2=J�=u�<9<�X�<�g"=0E%���J�?^��Kk��'��0��T[��|@��^8d=&
���D���m��Ｈ�[�ei=��<4Z�Ȑ�<x�i=a��=��<I�=��~Җ�o�=юJ=ҟP;���a�Z��)��p����� =N��<��<@���GA��=c�<�T<�&���F�<Xe-=������`��]c=�x]=�=����a�i�gW&=�[6��0�<�#h��N�;h`����	��6m=b��<�j��H�<�~F�*F��k�I�J%����D���=<�׼�'��N�Y=ag=��¼}F]�3C8<��h�+�-���^��I���<S��&%=�}��N��<P��վ�;�6ջ���k�<����b�}8��=~́<]F�ְD<��Yм8#S�L���1t;WV$� �<��<;"�;}� ='=�#�o}7=Z�¼�����O��0M��\g�,OY�:3�x̘�����<����~?=��~���H=���<'R�;ζ���;�0�L�*���Q=>�=�{�<׃���R&=��v=��<=U���.z,<��*��@㼿���cL;��c�<`D��]O=R�4��ҏ<��;=�ac���=�w[���}=��=��?���Ǽ��,<�Ƅ=��<>=���<����)M�;'�<��h�x׾��8�<@2S=�R=���ܿ��u��Z�<a~G=��c���=}~Ǽ��0=7� �J�X=�6<3=������T��<�E=Y/�ts���94�L�̻�E=�h����X=�t3�\�+&=���<��<o���w7�]�>��x"���=�'t(��3�<1�=<�h��[�=�����SZ��r=��	��<qJ�=�E�p=�(=��_=e=U=�l���L=�����$N[�R0�_(Y=�u��)���O������d=l�;p��<�º������<�o����Iʻ��<�@�<^��<���;q(c=�<R�.=Cj���y�:��&���<����	��� �����<���<���������o�C0�<�)�<��R���&<7��<��v=��.<��#�~�a=��d�!������@<���� =���<��E��]�<=�Z =&�ӼIߺ0�J�Ǣ��;⮼+ �����T;���� �Լ�2b�15=���<��弄D��,?���Rzc��3=�G�ڳ=BFl��Py=��;U����ͼ��Z={ ����Ǽ��)�� ��
(=ѭ�<�%<"5¼=�jn�)�=v�=�P��*�I;����$C<�7 =:�Ի^� =ʛ�<?��<��i�(\ؼ�n�;h!><�_F;H�b��>=��L=��=H�������@=|��V��D������DF=��
� /V;��==-��1���<B��<�]ʼN��<? �;��F=�6��e
� ���<����[��F�<�'=e��<K�-�[[
=�9<����O��<�V��=4�0Bg=���P�U���7=�yO=���<�� ��ļ��c�K=d<?v�>`=m�+=�����;ػO��ӝ�:��v@�<#g�t_<�{X=?Z�����G	���G���M��mb=��a���$�_�/�,k<~$={<�����H���<..;H��<c�<@N`;# =I6&= �:|1���<tGi<c�����;y�������nS�?�<�xs=e�=0��<5�=Fq =d]�9{�� t
=�/{<9��<��O��0:+�/|�<�N�*�;BjQ;@�^=���<&��<A�\<��N=E�=Z��E�D��͝<���;��=�I�n_�c��B�<�"<�>D=�W5���O=Y��<:�.=xzW=���9�"<���<�<�!"6����</�<H�=���<�Mr�Z��O}�Z�C=�F=��<�+=/-=��<��P�A�Ƽ}oӼW��;��0���v= ��<�Aڼ@¼̰�<�HP=���[[;<��;��b<g%�9�弿9��v=!�*<�Jj<<S�<{c=�[����=j���
X����ۼX�q<�-=5����<�3��9U���4=[T=W����m�;�+H��?�K��1 �΅���Gp��.%��,;�C=_S�glK=���N6K�RC=��<��a�dd�e�<9�
���A=m7��&\:�]s�����?���<�Cc=
��=���<`�<Z��ȓ�퇦�����i�<+�!=t�+=�<e�@<;�� =�&�<=Z$=�:���2<V�=�| ��^a���o=5�)=^!�����RF.<(���pP=�_�<��=\�b=�w<<d�0���u<�0-=e�E�����j�4�L���2=�`μ@<=-5;Р3���#���E�8�C=�=gt���.�o�)�C�<&+v;�����e	=*���V;fO�q�^����<�6���<�L=0rS=��t�>�@=H�n�-r=��=B�=G���I��VI�r�;�-<N�?;N�}����<\;<�y=�켱3��2]�<�m�;׆���د<����I��^'=Q5���+�<F��$�`;�.ǻ/AV����;o��<�8.<@�ȿ<��D��#�<�j�[��PI�)C3=��_��5=S�=���W�M���0+�ϯ�T�Y=
�t�Ux���;����4y.=��f=�#/<?C���
9��6��c���<=�TI<y��<���=�q1� uj�}�>�Ό�f��;��D��5�<�)l=�dH=�y��^>=�21�K�<�ϗ�M|O���Q�#��<��ռ^h.� x��gZ=�0@=Ψ�;.r=je�ڟ�b��%�q=6?=�Q=�;�A<��ͼ_Xk=դ��H���ؼܻͥ��&�M�r����A(;�=�WV<Q^�<�
=�$%=�[�<(��<֯J�x�:�8��_�T�C�=Qr2<�w\�M���P��C�`�!L ��pe�C1�<)�#�8l��WK�[흼#>��kVb=[=P�K����<���*��;�=M�<jۇ��:+=R3%;AV��)^��e��m=�o��p>���u;�hY<���P�\=�l=�lC��'!��=׻-�=�6M=`�==��:s��9������� ���<G^��0�q���W=�� ���'�J�	�����Xv<=�@��1G�:����6=�v[6�
U�:軑<<;�v�e�g�8=�D����<����Br<ⴀ=�'{=gw<<QI=鰙=�b;n=u�#�Ƌ5=xv<�#����d� �D¸�g�=���	�6���R��<�=��b��&��Щ<:3=�9;��<��O����;u�!��UR=�����<Э��<��;x!�D��!=2����X$��̼ן��� ���Y=G��<�8�$=E�m��o=h\ۼ�'���I���;�mV�����Y��jFݼAD���=��Y��q=Ƀ�<NBV<衉��~�A�[�&�@���K�͚=��N;��ϼ��x=���/L�E,��q�;��C�ê <XAK=;�<�3=	<=c��R�<*�V=�2��I�G=�҄���E=T$K��0�<%�]=_u|=%W1=dq�<���<6�N=P����A�_^�DjQ�{�ռ�o!=�T�<V�g��!�;s��M��b��K*�Z�;=*m;�ea=}\<d=�
�P��<<H0=��=8l�<JR<��;c7F=�Fx��Qh�ؼ�;�&I=����'=�Y����ٻB��<��k<�s���K��Ŗ;��0=�Y��C��<J�>��;�h�+=�Ĵ<��:<%Թ<��޺�/�<d�S=��^=�E6�?�Ӽy�u����=��#=QP*9N�ݼ�<�+
x����� Ҽ�'���#�<!�p�_ҏ<o��=b���m9=ƇɼM=t����Ƽj��7�A� �d���;=;b<�ea=�Q�2H�;���<�+��tR�=��4=�%i����V�;���H�;<��;��:=V�Z= �<��;<C^���IW����U�D=����β<���<�j(=0N	=(�<��;�ovW<�K�<U�_�d�ɜR=t"D�ϼ(��j
=Sr���=y�ƻ�r3���ռ;D7��g<�	�x�B��F =A	��E�"0,=�0��%=&�tI�mb�;�X����Ҵ��~<>�}�р�92�<�,���i�:�\��xք=���<ԝ'=��^�w@I���!���<C�(=Ka0=��<���<�^=��=�4=��=}���-R��o%��7	��3��H�j>_��2@;����9�^E���~�8�c=a�=YG=����b=>�B=T�w8�L	=z�[�T�.=����H3����M���0=0DL=��F=���� w=u��<~�<V=V����o=���a�<cI���Fȼ�b<��/=]�Ƽ(�[<slK�B�x<@o���&�����<%�Լ L@=N�;�;N�l)O;}�<c�V=| )��8)�-��;Y�<t�� �C�B�=E�<��ʼ�p�-.��S�}f=�#�5�,�?�Q<DH=<�Y(=ڻ"��=�9$=^��; �D=y˒<�/=�!ݼ�M
���G�f5�<#L�<�t����X<��{�N:���n�hV��%|t=�����A`= E�CN=���<�)
=9��pѯ�KV=�^�<�˼�o:��E��+߼�!E�d�<R �<�&Z=9d=��;5e����<i_�{�<lp^=e����C=���^=<��<��J����;\D�g޿���=��=kD�}�<DE�?Ը�"*���9���E<�6��C<��<<}We��r,=�+)��X����<�&#<&Λ<�`���(=m�]:by$���L=MJT�]�S��H>�0?N=�����b;_�]��u�<��f<v�A�m�=��ļs�5=:��1���;���M=�W�<j}=i�;=�X?=�"��H��<Fn5�����<�;m�N=|�;�li<R%="�x�A=Z1<i,<�M=�n�4�`���x=�X��ܼ��<�i=D�<�{(��9���ɺ�*��GW)=;��g�8<C�:��^=��=�<OD=��ۺ
�<�~�9[0��z��7���vY<�j����<<��¥�9��X=i�A<� *=�ݹ<e'=r��,27=�F�����$NF����<�W���u=�s�;�t��r�e�.I$=4�<3�*���S�DzM�?[׼#��;��=��;|�u<�.=����%A���q=büO�ݼ��� ��l=;-�<�[�m�[�sݙ����<���:��=�PԼ?𻻎�漁=�<��}=����;��꼵
&=�"̻S?缆k����@<[�ؼ%�=��e=,����3�����	B�<�)�<��=5��<i�<]!=�4�<�& =B4D=ǋ=�����"�m �S�C�Ep�8��<î�<C=Ƿ=E!<�`=��|/���<�W=-�m�TC9��Iڼ�"=_�$=}�~<o3[=���I�N����<�޼��f�#�<G�;u�D=F�!�I�м\�.�Ay�<�;+ۼG��<�v�<����sg���2=-k<�"=�W����S;�=�,<,"�<��$��i=��/����<X�x�`E8=��}S5=�!�<���<p�;���鼼����/�@䲼�'=t=���<�]=�t)�-�&�n�,�$�<����x�L���;<�� ��=0�=�O���<���<���p�;��=W���ٹd���;��k=c9�a%&=_/<�0�<- ��M;�_hL��`3=%B��c���->=,��Vܼe�=+��<���<Ʊ\=���+<[�S�F��<��<��g��}��"s�[�ƼS=p�^=w�>=%4�:v��� =#���'=ރ���S�;��H�3�"|ȼT=q;f�='�;PV4��=�b	=�[�<���<p�=�Be�#%�<,�<�y=Ȏ�<��_�]���=	����(��=����H��g	�<��"��1�<��1�}+��m��< T�O�J�g48�{�ku<MF]=�$�<.&�������=��<8�=]�@�s9�~�ƻW6��3�"�#qd�A�:v��|K2=$��r=/�;=�u�<��\=���<?R��(��<���;3+��+U�<���<�F$=2��<�"=��<�L;�/�<��<l�=�c�<��<�4	��}��J�aF=ld�3��X�J�,�<F:A��-`�$�
=��=���D\ݼ�
�����ݼ�B�w��@&5=�滼���;�23���%�dfv=~ػ��=�Q��C=C���$,�;��<�]=Y*�W7U<���*-�$<=N��
��<�ř9
:=w�0=ǃ~��u����9=�<ځ��s�5�x�j�;R�e�=��V�4F�<_�f=`r�<�c+�dĄ���+=o�	=�����6���1<��|�$���k�l�M������44��LM=«�=Z�$����@Rd=czk<G�Z<9Ż�=�Zؼ��N;���5�)�<������7�<%W9�	�����<!;<�/T:��_=��L��a3��,>�����U<W�k<V��<|N?����YW;(j<m�Z=�\�<���<��O�?*=�Ny���d=��)�P��B�<�X4�8"-=�X<�X5�w��h���<ǇY=Se�<�p���v����zu�a/�<�q��8��#<E�w�%�:�B�<{%@=O�<�qO��֔��57�bf�<��F�/�9=DV��s&��Q�;�q=c�ٺNY=���q�_�PMj=%n!=��F=�Ǽ�(�<$�%=�=�X�����E�#=�I�<S���#m�D8�<B���#=+%A=�ru��T��T��~�<;~��!C�QLE=N�<��<v��:�<�+��1�<�
�<Tu̼+=Kd�<��q��ڼЅt����<��*���=�U<|�9<	y���n�J(M=��@�F
t�ub<N\�$�(�Z�m�rB%=�yA�!����<����G�;9�]=�	�<\[��3�<e�T��;��)&��?I�T�g9�u�<@�T=��{<1G	=�W1=��U�О ��j����<f��<�h����&���?��=��=j��I4��4�<�h�Q�E;����|����DA�-��<�`=��E�ִK�EUI�|P=�7�;�V������2Ѽ��!�f��<vR��7�<�v �(D=NO�(L=3!�����<��~=�(��������'<�X���%�8=O#9=��F��}&�.�����=���p��<�����Si=�LG���(�_�\��V�s�<Γ.<Q������<�$��T=��=���Xm;c@N���L<sr�h�e=+�*�	�<n���K�����l�u=��h�A��<��U=�	M�H��<�r�<j��ǳ��C�D=5�<� �<n=9���v=��P=��b=xdC�Ȁ	�:�<n ����ϻ��O��/�<��<{��<b�h���=��<�.(=�����E9�\=�՜<��]��P~�x=�߼��Z;�Y=�5��U+=aNA<��y���J��H)<��s�a�==��<6������<l+-=!�E=�u�m���
�k�"6 �u��S�Ѽ'	t==T�<�R;m��;Q�E��?=���l�`=d3`=�M������_V�3��<ωƼ%"W���=O��<����cV��[��vʾ;ZV<�I�<J���:}F;�+%���<�3�2	a�����ˬ�=����'=��8=o\=�=
�W=p0 �9��3��$�DF�Zή;3}��0=d,�<��u�Y��=��<��+�-�j�Y��<��A�]��=/[J=S��;�m=GS1���=�	=��==�<K_%��a'=O�@=���T�Q���G�ټpjR�8��<�;��,,��f������2ڸ��G=%�=�=��ĝ=�+#=e"�<�8>=U�	���=�3k�C���x�=��=R�S<Av���Rz��j�<���L��������μ\��<�l���;�H=U�V=_�A���U�
��L��}
���E�����0��:^TD=���<B1%�#F+�zk��<;K��O�=�߼U����ȼ�j�<����N�<~�<�J)���=�O�<!�K�i��<K�ʼ}*M����;c׼��b=�;[S'<>��<�� ;��g�<�>#=�Ǽk��_[;V@=Rs���ٻE�y=^[�<[Ƶ�ޡܼ�:-=k��N�I��j�<�Z�<�'��",=kg��%k�<bp�<�JW:rzc=�OռE�Լ?�x=��������>�1�n�H����&=�<�<�>���}�:����E�BtM���;����B-�Q�2= �w=���<�J��=b�aV�<=��<��W�N�J=�y��N'<�F���/=yP<��7=�=f=Y�$���r=0�=������<I�{�\m����p#=ۗ#<y�X��"c<�=���<�Z$�~?�<I�*��A¼�ځ<<#�Q;��O���>�K&>�EA�<���y�,='�:��!<p��<T��`mG;n�B��켆bw�pYG��0=���<���<�n3�<�Ȼ;7��|r�T�ɹ;���!.��&��d�;:�j=횵<=�<,7�<_� �9㈻H�G=�J;������������'=���sr<|!=��_ۼ��=b�@�q=�֏�<rBƼ2��1<���<.G{9[��xƼ��5��;�2~<?5=��9;�x_=S��DG=Y8�)߁<�*=ˢ����O��,���;=�GI=�ҏ�J":=r1�=��<���;�JU=F�3=bNV�Q�^l��Ѽ���8��<�B[��Y��t�;�ED=��$=Ir�;��;�Q�Žd;�J��ޔ�T�g%��0h���1=���\�<VG���~=V2�=|W�;���R�'�<3t=ӄ�����O 5=`�Y;RTм��k=ƀ�;�)�<��P=��_�w'=X�;?��<)ǁ�.����,=�
�<1�;�㈼�A=Xx�;ͷ�<��0����;�ϊ���^���<�l�-=��=��<��η�c6=�$꼓"ۼD��<��7=���<B�����<H�<9j�R�.��g/�"�E=<�Z<���<)ϡ<n��<�>�~eM<�G�B�#=1'9=�!�v!@�d>=�,<�q=�e�<�Z��D�_2��I�.;��K��eF=F�)=�Gj�b1��d\�ҭ�}��<��o��M��P������ΚP���ͼy�o=t�<��O=�<D��D=Gq�=������[����<�YJ;�v-;�;����<SQ=]TZ=��6=�t��v>=ʼ�f-��p��FgE��$�U<��7����Z�=�z	��� ;d@K��J!��s;�����	=���<9ἴ�л�sn����=~eG=]V��3�	�6=�;<��=�)�;[�;��9=�b�8 /��ف<���P'�<�o��k-=�=�lܼ�m�<���.�޻:#K��t�Tc��C�@=r��X��<0JQ=�\�;�iK=�u�:�`=��[�N�`���0=s�$=P��<��k=@�E=��(���@<�����;��;:ܾ����<wV�=�=<3��;�;:�=�
7��k��Y:<�;��E�<��&=ɳL�)�t<Ʉ��I<C��q�=��6= �=8��t�<th=��F=��`��:���{�N�	���4=��1=r�;Ҟ=��5ͼSD=�9����U�I�<��[=Y��<S�;��Q�B$�;��<��s�-=k��<9S�;�x���mx=��/�)oż�G=�sŹ�2�^�4�ǃ��@�$=v=~M9�K����2�����r	��a�<7(V<�3�}w=��=�%�����S���M;-0�<nT=;+�<�S ��N�}ڼ���;TkC=�~���@=zGR<���<� =�!=�@�;5�<D����<Ǻ�;��7=5�~=`o���4���k=zmͼ�e�;��Լ�(񻕏��ֽY��T��#���NP� �K�	�=;L>�;�`ļĦ�L�!}�<ނ;��bX=���;X4�����h%=5�(�|�<k�3= ���]�?���]���|�J�=����<%)=io=�l<��T=�=��=)��<~F��Y=�;��<�c=� ����6�L���@�Y��<����E�4�<;��<�Ѝ<���J=e^�>� �>W���<G$���b��RC=L�t<^`=t0߻�E�f�=���]]-<ۂ��+�<P��y�a=r�a���=,M8�ۄ^=R�=Lܡ�lX�sx�cق��&<}��,��f��A�<�=�:z��Ru8���>=i�S=֖0<۷�<��&=���7QC=H6�<B�+=F��<}JU=�&+=�Q�N{J=�l=�o޼�uм��=S���x�Irڻ0��<֞ż�=��Y=�/X���p����<|�y�a��=��<2=$u�<�ټ��漿Χ�5�����[�<&���T�����{�=���;Vo�׊�<0���E@=U-�<�6<{=���<�N;=~Y��/�<��ȼo�ļ" =�9ջ��"=��Z���<0�^=�B����<fi�<��+�3Ļ��=��<�L��<��o�C=���C�z=jn����P�����r�0k#��z[=�s��9D�<[['��~�ʠP<o�=ϡ=8��Z��<��Z�yB2�\=ڳJ�rh�<i�]��T��=��r����0H����"���R=�Ti�-x��fD�$֬<&߼� �<���D� =���)�<�2���=�7=�0:=!��<%�*:=�߼���<�w2<.g2=�3m�̛|=��8<M���x7�h��Kb�;T=Z=�>
=�yp=��=;����<	�7�Ͳ=�v=�XV��c��dx�L =�����W<��[<��=�=(K�;�"��-�/<��/=Sĭ<��@=�^�o�A�����ת<��.�M��%Iq=,�9=N
.�Vm �H��<�P�<���BL�����<����d�=�7=�J����_�r3q�<Ap����0X�<�<w<�L��S=�aռp���2�;�sZ���h�x��:�� �9d<��c�b��F�=n�"=d)�<�|�S�s� ��;C}4=1=�:�<�)��^�<\�-=�ZH=�"���5�Z�;0�l;�=�(�<��@��eڼ�@^;��Y��R�2E=���!��=��򍽼���<�,�=q�<FZt;��w��ּC$���Q=0�<z=�TI<ч<�Vs�;a(=���%<!q=�-˨�#�F�Ŀ��;1(=�tL��y�<��
���-�n��<VB�<.�H�k褼�ՠ�(�K<����L�ܼ%fF=��"�g�d�k�==���<�s���I@�D����6r<�F��傉=��Mڼu�L�'��t!� @a<u�%=�'/=��a=�{���`�\����&���R<�z=��R���=�Q=ƹ::��4<��-��å<�1�okp�0�d=�i��9�<G���h:�����<�Y׼@�Y�&��<M]<��W4=�/=��3=Y=z���s�<V�]��iF<.��L�9�	�&�{��yH�D*���!�<�z�v����=�h;����xu�=��j��:�;a<�����<�*1��~�<�d��d=��0�c�߼J{�_�=����	ȫ<�q_�,��<���<�	S�t#�:X��Y���	=3Y;^��3<Y���=�|}<;l�<�?%=>��-#= �<�<Z�m<O�=xe�ƀ��d�K<9{���S@="�*���+��V(;�.<��8�g=�N;kJ���#�t:�<��6���7=����g<?�'<���8��l�_=/3X�O4��s���[|<�9=�rN��E2=jJ�<D���d;�V�x7��<�";���:�Dy�VT	����<I�� ����
<�+�-���f<;]׼�4n����;��ɼ�+=^xm���*=�Hռ�=�0W=�a=[c�< yw�9��<mc��f���m</����^&�hKC=��r<n��&�2=CU�<E�����F<�B<v�j=)�%;�0j������� �|��<t@�<��9^��ɪu�|�1���D�xg��k9�ɡ�q>�<���:�e=����E��<��<ԗ�������.P<�����ߖ=[�=�GH=�h���"(=�o%�\*?�)|@=T�D��	<��4�!�<�Tk=�U[��/T�2���,Sm= x��ke!=�_���< �<N�,<��X=��+<��=[ɼ��/�[j鼜'���s<=�;�U�<��绲v;<I@==�`��Ģ�Ю<U���~��4�<I꼯�߼~�O�0Q��i�kj�<U�d���<���L�Z�d����;�ḻ ,�q�)<�-
=�%1=����8�<�(ټ�7b<ɢ��\���Y@=|��<�<��~�%���<� %Dg=�'<�<v���@;ݺ[�׷����= =2�7=��0��#��5:�w=%);�L�=�#=�}�1�м�6�Ǒ�<bmO=�8)=�<��E=��<��2�:��h���Y[=,)=�8�0tY=��,;�&ع�lY�F��;��I=v�a=/���o=v[.=qF<=��e=0%�<#�)�B����O=`�=Y�=mw;���=����b�<���<�`�a=�<d�v<���
�S�3<��M<�ܼ(�<�m	=E=�T� =��x=,�T��=L�C'w<�3�� E��9=��D8%X�w���Oj=,�<��h�}u�<s6=4�<<�E=�wy��W�<`��1�I=!;=��=jV�G�`��/��P=����=�޿<�M�����[`<�X��Н�<!&���<�Q�LQ���-�<)-�<���;`��?�<�b�<�c��.8����σ"=�1=]ww��-]=(C2��s�����F�; 'R�L+,=�C�
8�r =�=6���	���2=�.�=������Gs�A��=�M=�e�E@j���<[C=y�O��]�!�3�ba=,f#��b�L@�W�=ڒo��d<%�=�,¼���<��=�y�+<��)��=�+U�YN=��W�ˇp��_
�L�=� �UM��4=(��K�S�E��\��=�x_=rH<�7r<.Լ���<�����ż�Rl��`��ށ���<N�����6�����|Ez=����5�;dQ��v9�&^�+�<��*;fsU<�!,��C�%����R�T�*��q̼ɤ;&���IeL<&D=I����Y=h�)=TU��~�<9�=�	h4��z���<�z=֛O���={	L���
=_�Y=�=#�=e� �"�ļ���;�P��5�P�H=�ũ:뢒<&N��L��M�H�C=��<"=�g�<(_T�l�z��5<U7�DXλ�ͼB0�v	5���<h���P����
G=D'%=}ʱ��9=Xj�������B=^;C=�)2<V*��G=ߘ=%<|m*=2O= t
��,�=�[�<��3=;n|;�=C=�|�d<e7$���<E�V��,y���]�5���d;��U���j=��D��\����ٜ;�"=XI`�U��<��=��:�����<y�=L���^Q}=܋=�Ǻ<�}Z�e�5�m�?=A&��γ;Snͼ�a���],�p�Ȼ40=��C=��l���<+Oz�����D:>���;�@�<�ﳼ�füIA_=����F=ť�;�V��^TJ<<$>=?8F=��<q�=�S�	L=4��<.k�<� =vA�;p2��似l��{��#H�y��<��o��W'���M<�7<��@=��a=5��V��y	=�x=�`3�q���97l=~�3=�V#=o<�<�U=n��!4R=b�G=(��:��w�V�A��'˼��<=h���=����n�<��������4~C<��<�pȼn�^��=���<*k=Fj���Pؼ���q�;��=��f=%4=��=Չ���_=���zM=Ҭ���%<�˩<v*����b��g<=+/=�&�C�K=~Ʌ�a�<��9=�0��^�+Sm:��m��W)<6�L=�9=N�?=h����Bo<i3�:�=:���e;��0=n� =�]C<�1��sa�E�C���K����5�;���-P�V.�<}�����8�T�s=�b(�%�*�3���=к���8���V=1�&mֻ_]����欼-y�;3C�<��Ｙ�`�|r=�.=_aM=�"r�W�M��G=�Sx��@R=��e��Y�<^-�:�:c�A�=8�:==��<,�<&�=y��������U�62��?�P��)v=g�Ż���<�̼b4�<2�H<u]=�)X�&�:=�<(�=L��/ ɻ���<���� �<{��')<?-�9�n�K�<=O-� n��\A=�\�<$�ۼ��M=,��-Ez��Ӎ<��P�z聽wl	��'��f�!=�"P=�cs<�D�%������q=w�Y��ɦ�T��6���T߼��Y=7 ��>�<o$=ʡ��~2�K7Ӽ��=�ƻ�,�<)�"��|���(���T����<W��=*�������<3��<��f=l�<h�3=��= #q�Sf==^�ݼ=;=��W=V{�SeJ=jڂ��d= �������w��]�����<�NS<	����{4=w�<�V-<�dH��3�F}�<��S=qhB���;��Jl�S���U�뉦<�)F������R={M���<{�<�����%!���L�Y悻\I	�ob;^�=��ݼ�pD<�'�<���;� ����0j%�gFT��8-�.ʭ�-:=��h�'ys<S^2<�d&=��;r�=+ӹ;߬T=�=�PQ��rr=Sg!<�]�!��1=)�-��BA�E(��Q�d=��I���$�0S<d� ���<�b�:۪c���<Z^������A��h��<C��<�J=U75=2
<<|;��-ř<��ںܐ1�* (=��]�+�7y�<�;*<� <���Ar[�d�a��(�<PG�N~:��h=���;BjQ=}|��D�@�K��<�7%=��<�n��@2<;�ܼ_ͼ�s�����,_+�1萻�� �yK�����3�!=�@.���)�M��.&=�M����c=<�/=�Z=M��<��05F�9�W�S:��lb<���<򂍼}�ۼ�b�"�ʼ�4�$Yk�\k�<@��<p�=�O<�����c=���<n�a<�fh�n�=kA�5:=b�#�Ȋ.=�ˏ�BΆ;�!�<�05<��n�Ww �R~<�*=?߼*S�;L�ɼ��;[?�<���<c��<���<��=����~=i�<9W���6�<G���e�<&���߫��4�=���<��;����P=D���T <�N_���sIt��� U���꫼I�J=�#�H�@=4�M�Q=��	�1<1�=8=C��<�p��ֈʼ2o�]#=��< �[=X�<Q^�=�q�<3*=:(��Q���c>�6��}̼��@�V��g������<	�;W�%�1��=�q��$�Z��<�d�+�<ׁ����^�P݀���4=4�=���<�֡�����끼�3
�{߁<��#�zӡ<���/��Y�Tk���}�cr[=P�<dJV�3A=���<Rg<0e;Z�=�u���<��<�l�;�A!=������|=|�;�<��T<!�D=G����j�,
N���a=��.=���<�P�<A{ػ3�=���4UX��79���=���<���g��<$	�4�����Q� �C=�fF��<�&�q��L�k<�ߕ<Kl9=~]]�����˭<�s=L�a��xȼ����j�<��T=��<D3��n�>��9ݼȨc��ӻ<��X�P������<"���H=C��<z���-B<��<�v%���8��r�����</~v;��2�r�=L65�;b�;�8?�GUj��8I��=�])���=1���ۼu(�zT��=�H��=��]<Qn��ż�A[�#�<<�����yV	�c�w<}��a���W5�<���_�S�$=tDC�Āk���K�IW`=vU�;0��:�1�t�=�<S:�FμNa;�m<*�<x�����:<!<a�K����)�݋���<�Z����� X#�g�@=e�m=�jܻ��I=Ν�<�h��M�:��=.�.�6]�
��<ڳ���2�<4��<�$��
��=�;�=<C��;w���/��U[<�m=�={�=^8=9��(�*J�9K��=�g�<���<����9=��мkk=�*=�q��1�S��iH;u�_=�=�v.���X�PT=Ю�<Y�.�/�;=Vf=�k��������<��y�+�	�a��<n�<�q=OS��l�{=�16=���;�}�;Zl�<�3u���;1q��8���Z=_�/�{:t=�@�;D=֊2=��=�#<\\�;��<ڜ�<"ʏ��p/�p=����>P;�J<K�*�u��� �������PԼ�<��@���j�FZj=�-�9�mN�Ak�(�e=�1�<�*=αf=�+=9CҼ�j��l�G=�yW�B-��u�	�򌐼*8$<R�F�PjB=�e�<5]%<A~�-�=�U���%&�ݵ<��q<o�弟H?:�_s�A~T�G7ʼ�p:=���<������q��!���B ���<�h��j��'ø-�V=�]�<bS�;3��<�\�����)<��m=��<ދ⻫ʞ�B���Ҙ�<�N=��=�jP=��9.B��Ǭ�ӌ=�q��e����A����=��<��;@V=��e=ξ̼����6<^�6<��$��3�<��k�U�+��)<�s��?�Vng���5=�-�2�<<�8������+<vw���Q=j�!=\`��\��;`�����RѺ;�F2<���;����,:�8�2c|�N�ټIQP�q�0� /=^�G�12����<B���F=���b�=�&;Y�<�I�%<}�ܼ��\�)�W=r����L�<ذ=�aa=���<=����m=9"S=�'��7��<����y��	<�)E=
�O��_5=c���[g�<�.��<�>�<K��<P%���ͼ��<&��=��<��<������<�?=�üU�5=E�<Ƣ =J�`=B6���,<�K�&*�<�s.<��ʻ��;<�|=�	?<�(	<B��<�R�qD��j�;N����N����5CV=�L5��_	�=MZ���T<��=)�=�z4���]�� &=H�&=�@�۝�<1�<��>�)�T=�v��.�<f�d<=�C��f����J�=𶑼����U=޹�M���������[z$<Č��d(�:N=y>L=x==�A��o��6=��;J��=�@�V|��!�Q=���<q� <v�#<���=:hM�F���Ũ��<r����<=51;��v��V�==/7z���<��÷к�'K=Vk==�=���;L�;2�!� |�<� ���y��)c���
=�����4X�f��`�p��=�`a���2:Z�"�SDѻ�\.��$��芼���<}%<\e=����?�<
=��G=8�μ�;=��7;4����<,쁽��v=�HY</q�$��;?r<���/ˍ���=��/�A���2�K�<���{fp�k]��$�<�U<홾���<�ȼ]Y�QLb����:*wY=M�;h���to���Ｆ��<�i�[c"=g*e<�$q��X��w$�۠�=_-ۼ6����瑩;;'<=��,=_Ds=L�=�P�;�(̼�v�����;(�5���<<��W=S��S;����X�=;�(=e�S����׭���P<I��;v�e#��r=�$=�ۧ�ND;����O������<[���6������M<�:�ա���=��߼��.�b_�<M<M�z�<�@4=KS�E]�ҬۼTh=��/=ə<�h�Z�<�[F�sB,�<��h[5���ռ� |=}��=Bgc��漑��:;�R<n�=����@�=�%I<��<�0=T�
�Ρ	��Y�<�<Z�7<莧�Nh;X�2�_.M�D����p;w�̼v ����/=d���p�m����.�<HϼF�$�݌`�XeF����]�C���C�;��#���h��.�6ȭ�-d����4=Ś3�ܥ=��=IO
=�.ļoz?����"J=��"=x
�<�Z=(�<�l�</;�;�����p=(x���eK}=H��<���-`�<IӨ��Q<ױ�bΌ�^|�=�9�<'���O��9�70=3P=�nZ�#;�)�;y�U���u<��-��&V=�a��f����S<��׆E=��� }�<�;�>=�C�:�E��)=~O3�YwJ=H&���]S;�9�<���%8�<S�O=H�d�=�=��8��T>=Ɉ�G+=��/�g����-.=������i =�`��Tl�<|��<��c=�����!=d����:QT�[�*�H5C�cAb����<7�R;��T=���<H�"=�j�;��/=���y�i<])��|�=��=�e�<	���Q������z»�A2='�>�,�;���:��2�N�g=��Y=�$ۼ��K���Nu�;��P�/2���:Ѽ/�=���<�Ţ< �f=͝�<A�����,�����<>=�p�<κl=�/�r���2�=��:�	t���"<	��<�=��y�<�]��n��c�F=_�<�=R,2=��;��&=�R=�(="ּu�R�ǀ,�ӆ�ҍ`<�:���]�K��<��d�C��G�<6xO=Ac\;���<��;�o�@e�<�<�<}7=���-03=�-�<�i\�%һ����:Q'�<���<92Q�S]�<�[$<��t����<�� �Ǳ������o`<4����I���K<�%;�݇�P�Y= 0=�X=r�ټ���<2)�<B�o�`�%�!��<_�==����x�u%6<��=��<>����`�[���\on�H0<�0r��CŻa�U;j���=��<���<�'���E=�b=p�!��Nx.�`�<��_=�X[=�[5=Ի�:�:"<ăF��ԼP�R<�=�7m=ČἣX򼔊D=Bt=��<��E����� =�.=��d�Ʌüj�^<B���	=��<\�-�u�L=��;J�<y�<�<Ҽ
\F���4�0����k�ƫ<�S���+�:���ͭd���P=�ٻ3|��<X���K�<��;��f��b��}ӌ��_��>	/=��J=T2i<�D�<��<��y�;u����X�B7D���-=�r�<�:X���i��į���u;�s�(Q���<x���r�4�K!=�Q�d�<���<#��;�>=)c�<��<��h��轼��}�Ϩ,���+=�ϻ�#V�� <�rJ:=�.=H,�7m=A��v�<��=K�1<�	�<J&V<��s�η!=�C�M ���=?����/�I������8���vT�6/����Һgl���
��WZ���!�`��;%��;� V=*�H�����(�ݣP;�=<�|��LԼ�@�aa�;j��v����=m�뼷<�=�s�;�{ĺ�Y��_�<���<n�W��A�:F
=�u==t#='�<z������ռ,�-<�;a�yǷ<r�@����<��ϼ ��<��	�z==?K*<�-=Z��<=92<�5F��2\<����\�7w=�:�!�=��ڼ������<܉�<I�5�R?޺�������<|Z�9�<��S64��56=�]=d%H<x_R=b��Ta�:/90��Ӽ�7<��<�ʼ���;�����(=�.�B�=2\� ������;���<�%9=���{n�;�B���m���;^i�����<�5�Y=���$t <y<�?e���i=i�<�mm=v�1=ܘ=�d��;=�����=�%;�@��:�1�<!U=8W\��yn<���r�	<�I�<��<���[<��N�5��<ʺ�.J�<c���B=�y��K�;�^���U���ib�<�<;�9BļK���16�b�<?�1�@f<JGżD���ck:oa`<B/$=<���Nh�;�
�P���"�Q�<ЩY�&�K���z<#���tq����v�i�-=�6���޼ �6���-<ۼ�D<R�=��ǼX��<����V?��OQ�����ڛ3���d�7ؚ�'�C�\�!�� +=����[�����ռ��+�(d<��]=�f=�	Q=g���.�<{=����L�N�w�>���*;==�o�2�<��
�,焼C��o<�ػA�OO�<!�\���7GL����Gpd�Q�=d�	��=-�=��a:��=�S=��t=V]�8��< :�;(�����%��a]=��=�BF�<,6�<7�ǻ��r���O=H�8������<4�Y;��<=��� �}n���@�E���D:��9<�<n<C���Z<�O��<�=.;i�޼�KH=��O=��輕B=���<6��$�=���,ru=�p=N�#=طp�TB�::�E��M�:Nw�X�=h�;��L�T�e=���k��<�<�Y=#H��3; ���5=�D�<�;@=���*�;4yo�C�Լ�q+���~<��<�):=Q�0�nt=��b=�vp=�9.=w��-p��e�<T����8����C�Zܼ��<�ۈ6�NZZ=|"=�E_=�F��'wR=�6���yQ7<~�l����<i�	���Լ�tm<nW�� �<���\�⩆:�+<�T��&7�4��<��';�C�A?�<Xt	=c��<��`=�;��e�C����0�Av<W��9Ի+X���=C>�XQ���5G=�Mw�w�-<٣<Ơ�:��¼c� <���O��;�Z<����]�D�����.<D�+��߷�ݢR=ɝ=L<�����;p_���#r�Ż��k���dO�F�=o�:;��ۼ��=�h�;!m�;��D<�,<�Q��{}<��X<ޜ)=�HP=
��<l't���)���<���#�H=��y��F���9R+;�¼��|=��i�����+��^{��V=#��<���ֹ2���L<MҼ(�Q<��<(~Ż3�<�_;�D,��M����G�I�K=,C��[=�=����L��Ӽ#r��S�=;�=��u=���,yc=7�d����� �=[)�<���ʕ;x����oE=su�<���<ڄ�<���������=��Y�Ӗ=<�<�� �:�����+�k^�6&Ļ�Z=vP��L���J~1�_DG=�&�%���$qK=����<h_=�/=)�B��$=�B=���<�9��e:�vV9�8����M���)=	~�;� ��<7f�<��h�����۾<��/=)�\=~��;�ڸ;�q¼�E���=�NA=�fm=8O<ֹ#���ya�@h�8����|Ҽ��R��r1���1�_�<P_<��<�X=�i)�7��<�:B=��Ǽ?ȩ�H�����:�a"ȼJx=Lz��Ԇ!���d=0�< ѐ�&^=���<,3�-
t�5�<w�����>O=@01=+�K���f��=Ы�嚂�{�S�`�i�\��=4ͺ���g8=�x�<�g���R= �=�tx=�<߼h!�=d]��~E�L?[=�	�=%�=������:��;�
���Լxơ�W�~<���_�;��w��=CN��@��!<�U�<fZ�ų/=G;�<|�;�df�g=��<$�<{ݢ=a��<[�>=C=��Z;rJ���f=��f�Qf=�c�E�/�<���汿�����C=�R_= �V=V��<gX�<�����Ͳ� 缄��<?�/=�<��<Lns��숼�X=	>�<�HH=K
y�+Wf���E�(�=F�=@ ��ϛ<e*=:BS�a良%|��SQ��
x�w=���9Rr�a�<�^��Tn���w=?��:n�ż!=���<�k�<,|�148�7�����g����;[�=�M���仠;R�./�<0�5=rK?���v��U����ϼ��={�I=�ؔ��
�:�<�S2<���<s�<�����hC=t���;Ob=ռ+�ya��tb0�wpJ��%��#_=��y=�`���<�P���tۼ- �<���<��;�剻��;=jT�|��H'�<�ǼP�Q����;�.=��x<�$��MS\=�!f=��?�����S�A�ʘn=6NQ=��K��*�Ʈ�;��`=��;Ђ���/{=d:.<zQ�<-��KR�ɭ�=hŁ;.�����<AY�Щ�<^n=��2�O=��=�4��)	�g�<�U-<i��8��4�*=���<G�D=s�!=B�s1"=@��W ��y��ZW=g�T=@%8��$����<j���D�����<1!�;�m`����9���<�{�<-�J�D=|�_�<ܕk���㼰��='�; |{��!���<V�3;�Lμ���<�C�хF=�9^<�F;��b<s�<I'�;�=8<9T�:���<4��0��j�M�6����E��T[��.�9�A=#-/<���=���>j=����(=�༮f��M�e�5=f�,=k���*�`�=p��<��1=�߼M_=������d��<���<�"�<6�J=�5;�i<���:~7��v޼�����>;hE�]�<��̼��<�R=fQY��="`9��^=V�w=� ¼�>=k/;#*�ً� 4;:��1���;��h�H�<�ռ�v�U^g<V��g��b1������6�1=<�m<r1�t�<�Pݼ�+<;����*<���1�t�=gmY=��;km�<),!=��=���ڭ<#^H;��@����<K��<��N��(�<�ļɃ�<�:=�w�<����	�$=C�ԻT=T�=��+��=�h=�?=�'&�Ab=�θ�z�����5K=J�Z�����[��V3��(��,9<_���8	�<�[)����N�l<~G��#>�;�g�;pQ�j��;g0;�h����;����_=�@��$����X}=V�=�kQ=��M���=6=_��<�<]=,=xP�<�$�=o�=?�����ߍ�<a��)�<�6���E=]�<v������d�����D��4�2������b<�+=iu��vk�<��=�Z*�pom=4N�<x@���X�мs�Լf�/�
l������
Ƽ ��<=�;ó����|���(<Ϸ8=(I7=c���=����=��k���}���"<cm����"���F=��+�����3�`=(�j�m(~�qA[��r?���(�=x �:ݞ=�X\�z�r<YX�<0pY�0 0=8Ԑ�������<}�6=S	��W�ǒi<�\м�F�e-<�9=!<(Z5�F�<ɹ���;���<�	V=l�c�q�1=��&=C��:�J=]�f=�v�<W������;
���VX��Y�CpN;��<�p�C�,=�;#=�3�U�+�򝯼t_�<���>��<?�.��~����p=��c==�:�cԥ���<��?=.༌H�<���<��c��M�<`(�;y���z==g.N��a7���=�u\=�C1�`;��A�
��<�Q���=���@<��n�6V��;��<-̈=�=�F
�y�=��'a
�;4�=}�E��0!<<`�.P���	=G-�?��g;�j�2=�&&�K��RD>;����u�4M�`ҥ;�:5=���>4��뤼�#H=��=���6���Jy���̼�_��V<�;�=��X=46���!�m��:���<p��<Ţ�<E�7=�e%=���<��M��#=3 w<1ƍ�E���|�?=g=hQ�<OT�<9��<$%�<�o'�˴-�)eN=�:l�O^�	A���S�Uz"=	��h�P=<�=��v�D=ĥ��y��evA=r�"��\��Q�<���<J�&��G��.Ĵ�aW�v�{���<٘u;	�L=�{m��y�<�"=���<|��_I*�ŏ�?�\�r�<� J�;��!=��=��=�r9=,��#^Q��TE�W�(=����Ǽ7<���f�:o���<CFI94N���|4=�A=�/�)g��z*=*��<F�3���Ի�!(=G6=ʻ�*ǻMö<!	�<5���T����i=I�@=� ���O=#h���M���껁��<���<>E&=����B�0h��+��CV>�m	,=�Q�<��!��[1�%=�����8=U�<h������<��(N��d(�<�H;[��B�'y<%��<
?���`=�O�<�}���_3=;?�+���j�;l���e]�;� P���ͼ_�鼹���<�Y"=��&<X@!=�?�7���9�=�,�9���;��(=�&�<�4<<��Z�M��<� =���<�ü�O�<�Z)=:5?=��z�����V]\=fel�.����k/=Qy=���<��<�F�+�������M���X/����<���<
��<g�;sZC�D6=}��<<�=�l=4��<3躍-r<��\=_g��>V����ߊ�bN��A�<��W�RB�<B9=��+�wҵ��"!=��Z=�b�ݫ˻3�'=�'=�)�<40=
j��{Fq�u�I���<���<>�<'�~��R��g�<�Y���(��ٺ�M!=U���{e�<m��;�<B���9=�ػ
�>=�I�<	du�`�M=�͂�D6�<�c =�Ls=�| ��c,;O�l���99"�^I=2/�=���<C*=��D=Ł=D�4���]�!�;0�	=��e��<Ӄ(<\n�d�7�=�\0��E=�,����<7hp<D�e�z�u�_�<������b<$/B� +�<n�v��[M=�N+<t�3=a�<B�ݼp��<��ϼ�f=�Wt=1�)�w�F���ּ3�߼_K2<p<1<߸�;�
�<�O��r+m�������^=�ا��3C���ͼ�r%���A�3F�<p��g�����Q��A=��.��!�=O�o�yk:L�;���&zU�VPG�	�����ڼֻ[�м��!=��ļn$��ed� ��<�.[�Ǟ3=鼺3J�#V��SJ�����t��q[��=��;�����T=��ͼ�D�`��<i0m<�j��A߼��k=�^��]�;"�M=���<%����Hc)��K=�ټ7�=���<�I{��j%�.�A=���=����@>=U�$�5k�(\i=��$=A��<&��<��R<˺Z�P�(��E���+���&�P;֐�;������u��K@�6GY;]����O"�eӅ�(r�<p%E=ȡ0=�,=~�缛����V=�ټ����ɰ�S�мv�j=�{�<D��ƞ����=��<���ߐ�<�l<�H#�2=\����:2���<�n<�T=�鋼�.=�p=��&=U�=~<¼ni�=T�a=�Ѳ��G2��<t�=��<�g��/*;/=m=�9�<��K���ۺS=�]�Y�1r#�d���^�;�R�"��<�uX<P�v;�̐�Τ6�
k"�v4J<�ڠ��t\=�^����X�z��<AI����<�S/=?|G���a<��=�ʼ���h=�?<=6=��:�������Q���
=2��<�7׼3�;��X=�v7=>�a��ı<a=��%=�VJ�e�=��*==�L��P��:��< F+�z�2=��)=�<<��;�SټQ�]<m�_;^h�;�Ҽ_�u��#=�H=^�w�	X�"�C;t=Bi�:�W=B=\�=q-�<Ӳ�<�M�=����UK�<!٧<�<�����5<Aݷ�[B=��3��e`�$��<�?�<�5�ѕ
���<.��]�=Vƿ<����R�;��=� ��qc=��J:���$r=��_�<�rU��^K����!�:!��oq=5Z<P�E�lp;�a�����h��-�<���R��<X�>���H;�������<
�E=�=uwռH�c=���;w�<h�-�܇�<� �;�[
<�<��L=�<��ʼ|N7=� Q=��Zi�:�mT=�3����ۼ1o7=�uR={��x�#�|�i��+T�s-�%,���=��+=L����wD=2A=���$C�H����=dC6�&�/=��Z�b�*ӏ=�;6=��'�_8׻%�G=�nμ�C=�S;�e?=W;��O���)[=}�&=��\�d�<���;DG�M�n�r��!v=��Z�bUI��Y�;M�&�%-	=l%2��9̻8uA=G#;�=L5d�
t�;�|7=�V=�<��;QaG�h;=���0I����h���7s�e����>=[�-��r�<*^1�O�a<4Ƽ3�(1���{��Xq=�M8��T����=�=RQ;	ߝ;�_ռTC�P`	=�Y��Ң�A�c=y���Ү;��	�N�O�O@�<<�g�?�e=V/�O����	�<M�μ�e=��0=vB��ㅝ<���y����ۻdȻ��L���~S��X�BL�<D;m=��<?r�G�#=4 �<��<�o=�(=��<Z��;I�;>�<2�4=<��<���*=��W�΅:="�/�"�#=)����=��� <��#=��<Ϥ&=�h�<xb<E�/;O��<���^k2=Ih�l�;�\=F$A:"μK|K�9|���=ԕ<G��;v=H;�I�8�<F�:=�+=�l���Qۼi <ԓL;!x���S����)�d�<���:��l���f�.����:!��<咑���I<¯�����=��J<.h(<$&�<�2\����<,����}%���"�`��d2=J��;=���<���
9#�L���*�����T����<$*=�|��VCq=r|.��!�(�;�����,�3z�<��=l�8=[/;K��������<�S,�Y�V=�TY��I=$��y�
��9=r/�<wx#<�����=F��</���5#8=�ps=4�<JI<�쏼�醽� =�J�;���;�<�T�J['���2=�r,<�*=�c<�#i;��G�:�r<ZZ=�ż�e'=�L;)��<�<խ�;:an<O�Ǽ�v�<h�=��5<�ae��X��<���R�E;��@���P���(<k��q����<E3��@];!����!�<I>�<582��YX=fP���������=�LT���.;3�L�x�<�"	=�<��[=�<�<}r=w0�; �"�C�R��ؼ{�U��a�iՋ<��;�`r=���:�b=��<4��*�=%C��G6=�������=`�λ�f;���<j�:��=�.\���`�,���<����D�c=1o_��Ʉ�\8=���K�!2Q����zii�`�=;|L=:A=���d��g-�<�.<�h=xje=]T�=���nR���g=6��<ʕ���6R��la=N#��U���<W=XN�<�e����v�]�}�tMS={ټ߂�<ki��$==��]��2�%.!�؊=��o<xd�V;<b�a�Z��d���/=��9��˃�w$4=��S�<��M�%8���Jd�_�0��Lm�Ur_����W�B��X�<��=�Ǽ�Cɼ��BмH����=���:�ƚ�]W�.T=�b<�X���f��� <�}?�w�K<�v9�V��K1'<�nO=��$=�
[=*Ł��a�<���X<o΁;��<�:�=T>��4�<��C=��D=�<;g�:�*A=8�׼Ze=~��<Dp;=�#�;�)�<�$�:��˻h�x��޼�ҩ���%��%��`5=�Q�<bμ��s�*��<U1�<֢�<�Qi�Ò�;#'�`�b<�20��ѝ��C=f��>�꼣��<��4=zJ�<��R����;)t�jIk���;��H=8��7x���"�´��>���q=�1�<'�Z=��|��9=��u̜�P��0�������<�R�<��z��ߗ<w�<=ެ�<�輖������<��<*��<G%"=�D=�1h�n�K�Ǘ\=���;�B�L/��ʺ���;'&�:�!=�2\=�0<iF�)o/���$=V<S����<��i�� E=�<0��X;djN<�	a=F#%=���<4f߼��0�st�ne�<ڻ!=����$=�uN��S=}+=IU?=�h��'^<[gc=���X{;=)@=`T;�ul(�Y���9,��:�L�+S��J+,���,���ɼ�󫼼|�;�>��?<18=#��<�7=?�y��B�����n�<� =B=�_�p=�)
=\��d�*���=�D?���;���\�[�I
=�9O�&a@�A���`~2=�ց=v�<�ӻ�:�<А�;P^H��IP���<��w<'�<[��<� ��.B/�_�8=`�,<.�<;m�;�$=Q�6=��-=�d�8hE��mS=��1=���:��5=0[@��mQ<;�˼/YR�RW����<�2.��	=^�<ض�<(X=�0=�~��������<ƽ=��E�AFu<�u�<�tJ<��|�>M<��6�� �D��Iw�ȐD��g	�ټ�<�n =RMj=�!=x���0�W��v3�\h<��=BNY=�D�H�?�?�����==?�O�!��I='=�[������c	=��^=@��o=D��:�<��V=Ӕ���=���ހ<n�f�4�<h�I�4���(����l���ǟ=.�I��H=B �<�����18��K���9�d=[��J'�;�h�%�v�w7�@/�$�"<�ܼ��!=��<#�H;H���eP�f�	=e��J�8,����1�Jq�;��<�҉<��g=H�7=�4(�ȗ@��r&=.p�R��<��F�ߡ�׍�)<�<<%���A�<����w��K=�����E�;o�P=��2=�|x���2����<��=<.=IN�~�=7n������=���輭���2%�-e��n`=_��<��h<UJw=B�����=���R���c~��rQ;�K�<f���*/='$V�6�)�#�;Ʒ1� Q�<2�e�Z��<Z���O=�!�3�2�����3�<��=a��=��b��Y����<�h��LK=>���fj��P�Πl���B<��;��;<��8��fI�{Z���T=���=����;��ɼ��;i�ӻ
?V�6*H=��;A�R</c�<�&��)�`=�������<=4����;�L�<���	�=2�w;�I�"�8=�00�&�ؼe׉;�<�66<c_ � =�,1=�K<8]�u �<ڰ;iɼ�]ļ�?E<��<���������P<�X�2�y=ks;��I�;DWQ=1��;`��ˇ9<���<ϣ�9���<$�+=��Q�̌����<e���i
;�=����O
�l�g��<�)=2�;����LY=*�Ｅ`$�gmҼ�=H)��h�<��;��!�j���;F�=�=���%�4��^x� [�<���wY=)ͻ��6�<��]:�,���>=�.=wq�<7�P�]=��</�x=��y=&ͦ<�>#�^KV��W=h�:�)����у��?����;=�[���Ӽ�%��%=���<��$=^��;Q�2�W�׼�LL����<AGG�D�>=��<<\�'=�VW��"�<�[=5i������[�< �g;_`��%!����R�3=��6�u�`�2	3�`62�C��JE����<D�<��<�=�<"�<�+�<�~9��Ѽɔ��#��gPǼ��N�;B�;��	�Ȧ��J�Hv����	�n�ݼZ��<�|�&�����Լsl�<Gd�;�R����<��T�U:=��E�o�:���;:�����<��M��3=��*��,���!�S�$=�N���~�ēW��Q=�Ü<�E=6��<$Լ?\B<�}V�d�)�o�i=>�J=���U��;�?=.�,�[Vx�&G=x˼�l�<�XG=]�=Zb��fV��"x<�qB=�;��;'ȼ�C�;`i廍����A�{=<^D�=�q=��=8$�X�=�cP;d��{$,��A��ɼ�%��	�e�ެ=�76��g1�LX?�`�= 6=�?=�.���N�a7�<��=��՗<�ؼ��J=ц�O�=����T]��iL�?����;�Q�<�ϗ<:�f<�`n=�=Y�<��=g&=�Bd��<�"�VO��#��wi��ὧ:��9���G�K:���e;��<���u�<Ƥ��������<{O={��<]0I�沀�����B-F�I\X;a�1�@=���ږ<�s���KY=���<=^�a;�X�E�.=�b�;�x�<��ük��<��D=4 ����<�S=<ɼ#�N��M��/Լe��u���<��}=�խ<t'���3E�Ӛv������ <��A=-[a��/���<�A�Z �<�I�=�?��$~�����Q���M<fGK=��<�ż��<'��:k#4<WB<EF)=�;*<�t=[=�:�;Լ�C��X�<���OuC=�Ԧ<�<=f8¼v.0��,μ2��#�m�L@�=d,%;MV�@aH��N��?����?R;`nv��4�?�=�	<=�/��s�j;=\s���=������,=�M��A�;@4"���b�<ϡ��������D�����7=��<I�<���;��=�,����� <�@�D�H�%=��뻩�����=�/U��t��g�<���;9P���	!�$T=U~'=��f<.��;�Px=�P:�2���N7=� Y�î�<UR�2�<��ҼJ�<��c=`m�bu==G�%�ۯp<1ꁼ�R&����;�"=��=$��7���ϼ�`��JZ=��;�V���HC=���a����b'���V<b��8��<�/k=�̄���"���̻}A�YU=�8=>K��*��$���g��mU�Z���򥼽�6=���=
�4=��#=b-<�޼)�B=����g�t�E=����j=��c�z�˼˪�<��P=|j�͊2=g#>���<O��<
B�����;m|`=�9�<�*5=iW�;����b<ڭ8<�g=eD=z`=��D�Co�<�ZW�%�|="=��Y�;{@������<o���5/I�3�T=VD��f�H����<�с���Y=�'.=�4��'݈��v<h�<�g?�ᷚ���D�gm3<r�T�/&=e���/[�'$a�*��1q�����=�%&���O�LTE<�v:��D=Tۀ�&�<)3=��.=b�3;�<��F���E��q��"=�Yo<�Y��y��<߶��>A���.<6��"�vR&�_l�4�=y`ͼB.��n��
Q'=6x<;j�������<�����<�Wȼq =��(�y�o��)�<k�<Q[5=݇�="� =�<���(�����<�
��d��
����=.�=}u�<g��<Πͼ�9k�G=B)Լ��=��=Y4S�M=;t �~8���f�;fz=Y�
�8]�bD=�z=�{�<���B	����E5_=�5�<��i=R�;�6���`=��N=��<Z=X�T=j?Y=�-�:�E�<�U�<��Y�?�V=����s-�nLʼ�;V=JE��d��`�28=�����x���=�a�9k�
;OG<��<�@@���=0 ��;Y�<�&=i.�<0,=/�p���<����S���0�j�ļ҈��,G=k1r����=N�S;��ȥ�;Û���ͩ<��n=Ede�\�h�q�0=�Y��;�;}#C=�e.=�g��E1��^�_=��<��*��3s<%-=��K=2�<6�#�-%м��ݻ��L�T=�8�;��:bz!=:O��X6�k<8�<=|���V?���=2:�<L8�<�<ĉ�'�P<1A=st=�]y�}=SB%=/2�<K/���V==TE=u�o<��G=��<�߼���<���<�s�v���;ؑ��K<��7j<����O��0=���:yO<�`=�_ :��=S��;���<����X��<τ.������>�v|#��T2��=ص�<5K-�-/<�I;��\=�=��4�γ1=��bZL�!�B��E=���/u޼(�@����!���=�f`=��0��$-����<~C�gq�ol_�Uc���>�h;%��̷�;`��<��#=�ז<��� �s�KAL=������<�g�ʻ=�qw=�ļ=�<ϦI�cǍ�_܊=-Y�\��<�C�xS=`~*�2��ژ���?=��_;�%+<O�<��,���=�"�?�=G�(<p��h�ͼ>E��ah�;/�<czl=3� �=f��dz4�ܞ��C�\������<D���!=�Y=�	2<��9=�i������<I1�SCb=��<NYU�H��ki�cg+�s6j=�攼�t5�Cfn���a������K=Y��=�S��C�<�k�<bk�9m�����=G�o��;pڏ=GVL<�|Y<�\�<�M��8ÿ;~J?��m=%I<�G�4.���&=A��¸l����Z�Q=uX�3�/�5�;y��<A�M<�7I��C�<c:�<q-R=u�<�N���G=?=A���t��� ���3=f_=�x<
�7<!1�]	!=j���$F���!/�j�=� ,<��������\�;;M=x<I�<P��Ӂ5��<�센Y�{�.=[�n=F뼻?^<}(Z�x�b�6��<��<�z��6���<%Z���0��b�z��;+1�<!g<
�Q��L���
=�?���=�`���T�gi4�S�<��<��R=;d+���`==#-���z:�^#�'��<�"����j�V="�i<�&����:�l�<TV_<}Om=I��3 <�l8�5M%�,�W=�a*=J�8;�'5=|�=�˷��K<G4���z���X(=�7=��G=b73=�.<܂��e���g������J��(=g-��h�<��>���,=Fqͼ2�=�X��F=�6���WB=�D@��z0=#�\��5"���2�2�<uO�=>6����i��|��r2�c���=��=U�����
�</Y6������M=�%C=D�X=K=Ny=��߼�����4���{�9 �<e��9�����"���	���K���6��d�ln����<�H==��;�G�<��p=�ꇽk�g=\�D:�<��һ:���e���Y5=��=�ý<�X+��v<���;��O�Q��4mʼG`�K-=9ڙ�̄.��vT=��<�ü�qv�X���O��<���=N�t�>��<7�=���<��<3�Ѽ�0�`�c=��~�C=ҳ�;�t�;�B����V2����<�`<���+j=t��<�輨[�<.����E�<�g
<	*C�Ɔ��袼gKT�Dv��?==0Y����<�����u�<��<�O��Vܩ���Z=;��aNq��%��J�<���Tj=`5�x�y�6P<�I�<Wb*�[O�ܰ�<�(=�-<� <�����F=�_=xS��]LZ=���=Yk=4�W=a˩;7�2�}/4�h�=�}:�z{�=1�=�V�<�.��_I<�߹�WH=�u����<��v������u��U�bhv�ՙ�p���3���6=�]'=�A�(le�J�l=󻎻(���G޼F���A��ڌ���������{+�vUj�iG�<��=�E�;fZ=>✼Q�E�"�m<�T�<�IZ���!=N]�<#_üM&K=;m<�3�<�\k=�"ļ�]���L��=�lx<g��<BwY�$x��ۗ�5tk=x��U�=�hV=������;�""=c����-=��=�~l:b�	=>՟<^�9�tE=?��t<E<���<�9��{���.�)��<r�ѻ�W���:9�dJl=��ƱU��)�b����J=��<�O<��򻌴p�^1Q=1()�47�]t�7���3��܉<�U��܇�<�1�;������J���d=YV�<-r=��C=}c��bO==�'���<,�=�d�<�&=
S�4ã<�(S���;�W=�,q��`=T:�:��H��;�<�)=;��:e)=�H=��=���8��>=J��<��Y�&�G�H�=��Q=�S�=�t��bG��K�|�~=1���;&�<|J��ϕ�p�<,Mi�#_��6�=5�!���)<ӹ���;���<���[�z<s�]=�7u='%�<$f�/-]�RL���c�<p�;�.�rf0��i��%���I<8��<D�<�9,�t�<��B=�4޼C]"=����~>=�'�<}��@�<�=����M��WX<���<5��q=^�4=z&=��<s��,́;*4=��^<�s5����<q��<JC0�/+C=A="�`��e�:� ټs�*��d?;�^=C��F�$=�h:�M�L�fV��i�<�?��/�c��<�z=*���7�Q<�b=A���a==im<~Uh��8:�	y8=�& ;��;�K(�$3<i�'=S�P��܂�jCP<h�-=d���J�0�ڲU<p>�<��<���d�.<��Ӽ��O����g�f�$=Q'7�8'	����<�T\<�< ���ؼ�zn=S���-&;��=��<ŷ=,�?�x�d��F�9e�u�f���2�U"9=����ȼ ��rD���L}<��N<%/׻�y=�y=�MX=}�;�#W=Z��{�z;��9�%�^<�x����?�$=�4c=��ݱM�s�Q<,�0�!U���� &X���_=�<�~�G�*�V���꼠 D�(I��^��E�<9
��Á�Bۻ;T�A�K�=��c˼���(<�=*�<_��<���<H��<�z�Vf�9���� ���!�'�0<�����W=�ƛ�[?F=X�<�_�	��<;�=첒<{�J��f�G�_��"F���<Q�<�N�<8�g=^�=��=O�
�I�=�����36���<���;��<�O���=�G�<�N�;��;��M��v�<
GY<�9���0<�M�<6�w=<0��5���%=E'=�� �<O:��(0=xY�<����$��+"=��<�(� � <�X=�P�;���=0=NgC;�9A=��4<���36�O�<�� � �;���<Y�c�E-f<V�R;���,9	�$�U;	޼a<=�m�;l�	����;	��(�W���j
h�m�V=�\��I'��&��K��U�[�S΅<�e=7A�<�N�=�4(=���!4���{����|f<��e��tE<%��<�YM=�e=�n�*Ƽq��!;������<%��;|��<R���gq��H4�p|H=�u=N"޼p��:%z�<h��;�q?�?�e=E7�E�=�X��_?���;�����,�S8<�U==-���Ǽ��==��;��l��Ǽ�U�<U:��U���=�_��S=
rL=�$�����Z;�<��o=V��<%W���I=�r%=H��<� ��2����\���<sͼ�0��DC�����x;P�|=����+��<(���=�_=�Q�	��<�Lݼ�l�d�8�{�����d�<1�;�u7�^UJ�-�=H���F��'^=h	=.��>ֺ��Z׼�/=&�?�%6ռ6�����\��I	��^��=�<Ĥ=z����<�hFڼ�J��fd�c�	� 1J�pI�<�a�;[��<8�=}|I�4��;'=�V�RU�� �=l<�"=ϐ���7��ݪ�z��I/��C��<j�T=�^=��-�ջ?�B�Z���e=�e�<��8�7=s$�<bW=u�ѻ�)==�	���p��*a;a]N�r�a�	�<0�=N}����Ϻ����<K�a=WB�iI��۹�<�hԼ���<  ^���z=�5B�d����D�!�/�Zm����%=�1�9�C=r��`�/������a<���s��� =H�����Y7¼:"�:���<4�k<��'��I1=bX���=z|)=%�����p���`��d��-;G�js���3�?c5=��H�?�i�[D�<�x������< ����_���_�v;��¼��;Ϲ��r�1DV=q��������/��>s=����yq=��2���v�<�?;�R���c���f�0�<��N�:���V��((��x=�"��=Q�m��[��<
�_<\N�;�P=`O��H�b|<H=�HW=�4���E=��<�|�\'@=��o��H=c�;V�����=hQ==�Q�K[��d��{�<`
��ܙ<V�����<ʘ�z?:=�zb��i��{ɼKüS�;o�=oԻ<Z�=�٢���h=��<�+;��@=d�<^�u�%߈; �Y�~4 =f�<
=��<U|<H_<~i<�_<��ѻQ)����H��<�t)=����{H=j)c=qg�:�)s��o��.a=�73=�3
=�(�� f<�P���u�<��4��o=d��O�c�jPp=���aoP���1�`���h<}��:�f�<���v�ռ�k<=�"μ����Z�t=˴�<,���T=�b=�DM�LѻTfU=F^�EP=�)��h$;��Լ{�=}I�<��/�W�e==�;�1hN��wa�KҀ<�O�<"����]=���<��<m�̼�k�ȑ�d�Ҽb�<���U�<�����'��L�<<R�;_����<x������2i�<q;��ˍ�f��<<�;745�$ⰼ���<�d'<�[=k�������fS<Z��S|*=�i����;�Nz<��Us����<��"=Hl߻��=j�1���!���	����<�y=���<�R.=z�+�+6��)l���k=^�%�V+�<�t�<���;0'�;�,ݼ��=rA�<D�=��==-�<��8D�{�J�
8=�iy=y�D��I�<i��*e���;��2���	��YY������<�nI�O�\� \�p4�<��X=��<�h��q��ܛ9�T=��
O�{��:~�=yM�< q=��;��d�S��/�L���-����d:�Fz=z�S��Jf��;�<�1=�i=��ʼ
t�<��=�S|=�=I��_��9�;ƻ5=��<��2������S�9%?<����|fR=�b��7��K,�2�ļ� �=���<��$=�M���'=�}|��I=�=��<�G�;%��<t��ͥt<�h;�m1�u��:Gy�<�\��	�x��-2&�.��<�&O=�.��*�叵���;yYn=�V�����)�@��Y����+T����N��ɯ<۟�;�0W<� ;w���!{(;��
=V�M=�l��G&=*ՠ<o�-��F�<W=j+���"Y����=h<��s<�����<޹4=�X�<1���{�;Q%�ޒf���L�T���j�"=[�<^$}=`''�)��+2g=�����h<u���`=�C��\��K���n=0͌<+&!<uH=��ںG�K=��h=��==���;٭��е�<m�=��;@'=��De����f��[j=��~=��X�Z��ح��|�<(�;(؏��%=����I=��;~�]=iJ=0��<����%�d��ȳ:�\)=��;[/�����%���=zGx<�����j==I.��d�=fҼ(�T�@��<��m<b3�; �F����<�/���"=��v��>`=W�<�	ü�
�<����3����=��)='Xz<2:�����)P=��M�G�0���;P�Q<	i����<|3�<���<}����<œH=^q�<�V <'�<[y1=%��6`c��=�:b���c<��?�l�W<��\=Z!�f?)=U=][��\=�;l�H'/� ��<N=.~<=����^�ucg<)!=#=���~�E�B�����u�i�\��<#C��	5?=7�.����=:�<O�R��%�#�T ӻB��<�&���:�g�$��<_�- =�XԼ�4����\;z�8<�K=�� ���4<-���<g=�	�C�J�/�@�}�a�<CR,�����T�<I.�<2�p��n�u3��=DEK=g�M=��U=����-��P�<�B��Yм��Y=I�h�i��2���_��Rf:�e��G�仂<��?=�b<S�P=��x� ��<_L��N��.�%�(sn���<�S��}8=����ʧ��t�=rhx<a8���]��J�K����#�<��}���<Mu������P�`$��p�AP���!=k6=�4<�@]���k��X��=��)�g��z��<t��<º�<��K����M`�P?�<3�&<��C�72=
o�<6�e=��<響��N��Fi��1<R����=��6�<���ѡ�;�Hu:�=��[�����0s2=�m�:�.�H��i��D>=V�üet��G#O��d=q�0�Y�"<r�� [ڼ+�~���4=�z��غ
Mm:T��<�\޼��K��d�;�a5<��O��}f��M=�+�;�W<�L��W�^=������<Q�=k�,;8;y=��=K8(����<� �;Eey<q�=��9�<r@����t�<��<B]���M=HC=~P_=��;��z��=Z]H=;=$�<4�D��ڵ��~��(�2������8d=�L�O�%=��;)�)=����:��M;2���=��;��=��<<pT��i{.=i,O��r�s�=�+�<�&R=��,�9�U=�6����<%N�;Nȼ]�ڼz���j�H�o��<����_�]@Ҽ�[����C,�c�h�k#W=yR:��"μ�h�A}�9$�����<6Gh�"�L�����i�8���<UM��`'�<g#����U�h���;1	V�4=U�� �-�<�;��<uQ=�1���Ȟ��&�<�v�	��<�����Ά�� `�6`�<S�$��[p�?}�X�A=1��;V"5= �=��:;+w;b��<�������tG<�P=�')��,����<�4����Լ@�= ��~<�7=���s���<�+�gy��q�l�)IZ��*!=_�,����<��J����|
m��4-=�� =Ѥ���@�<�=����r�<~�����81��X/���<�\t=:3=)7@��q�����:vE=�z�<��Y� �U��}<��;�u���:���0�`�����<c��<�����a�A0�;'���;(����p1<P�c�SV}��;��׷��H�=;�K�d;�Yp��J�a��-�G��`=�
L=TQe<�mF<em3<^���L�F!�n� =tܚ��ل����s�.��'=�I&�w/=u�Y���<��	�]ɜ<-2�u�=�ON�^��S$u�xf=�����8��<�D�<�� =M��]/;楡:�sX=M��;5�<�@b�����.�V=��0�J>���.�<�(�ҵ�=��U<C�K���o=x��<�GV�B=�k"���j�E<|°<K=c���R(�k���+��a= S<��7���:#�b�Y�8<u��<i���	<��+=��f=1o= �	����</�a=+�M=}�޼��I�4�Ҽ�����j=Z�<nn=���*�R=ȃ�HRB���!����;ν��T$>������H�P���F	O��*�<��c�c4A�^XK=e8<��=��Q��nQ�d$9�ſf=�\=�犼�c�G`�;)	��*X��P��Rl�;�k��X��<x�<}b�<��U=��<ʸ����'�������$=HS="M�<���P`=0̀�_>;��Y<�%�X�d��.4=Є=U�=_����㼭==Ӗ�<�?>�K��!��<ބU��:_<�16��a6=�= ={�<q�`<^F���6���m.�_%h=*�o<D� =�<V=�<1�==gS9���c<�I:=�{P<f�Ļ��	��� �A�ἶ�l�8͏;���V<��=�9���N<k-<����(X=E7:=�3���4G=<���Y�=K���g<�t��;6��+�9�=c�<�3c==5����<���<�>��K�?=z��<�<:un<R��زJ=�R$���b<M�<s�< �G�l4]��I�;."�;�;��<Mv�<A�J�5���^o��&Ѽ�i=}�3=W�;�=��<��	��n߼'�����V�19�QᅼRq��a�;��\���'=|������]�@�(,<U����*��`ĉ���T���H=eh�f"��J=�Q!="�6��*!��ur==�� ���<LOż��{=8������;+R���R�N�<�o�;�>f�����`)ͼc��<��!�4��zE�<��N<��<ZDA=d�=�!�;�Iy<��V�3=����$�<[~����fE����;C����f��anQ��X<��0=�2=I��<-,��Q=C��<Q{;����[�g�;����b=��.=^�V��L�7,H<TU<W�c<m�;'Y��IἝ�1��@&�\y����<�m���v=9�Լ4(ռ<�n=����E=ˊ���#�&�Bw+��]X���<D�9��<`�X��w�y�;5~(<�m�<���:��=�V=��[=1R��k#=: =_D��U=וT��^$=�䠼�ѹ���Q;���<,<$=��=ENg=�}69�T<j<�%<�##��5�G�E�w�w=�Oj���.Y@=r!!������l�H���g=����=����n����;c�M=��༭1��;3<S�����1=cD7=�Eּ�(����I%Լi��<��/�4���)��4����޼��K=��ϼ�I�I�=�!���B<ܯ=�������<z8M=�p=="ϼU�q<��d�_��;_=Ek�;It�#�8<�3�����*�;#����Ȳ�+�:H����[�� �f�m���2e�y=h�J=�*һ��<�l��<��<n7=�s����;m�<�G,<��z<D(�Kl<��{<�B�9+rU�5H�e��<��	==/��r��յ�2)��y�i;K@=��<��}<��8�-��-�B�'��*�<f��Wa�<�|o��+����=fO4=��<�|�<Uu=���<�QC����h�ټ���x��LaJ=�<�-�� <̛y��$���B=���;�P�j�L=�<~�.�Eoٻ��Ϲ��<��<���<�Y<�:+�{�u�d$̼G g=.b���:�ʦ�F�����"<k�8<UXK=:����I=T>��S%=�|S��)��j��H�
=ү�<Ln =b�������%F��p��,�󻷞�<R�M�gm=i�<�D�g>���
��샽�f���7#=��{<Oc�<&$�c��<��<�"D=e�!<oǀ�,��PV��I��g ������Ū���E<,9<*�m���6=~�+=B@	=�,=-�%�u�w��<��r�sE�;��E���<��_=���Co=��!�V�<Wq���qg=J �<���|���;���<
�W=�W(=��3<8�=��=��0_<шǼ>����a=״¼C���G�&);�^Ƽ��e��&=����l����;�4>���o�H@=��<tVQ��G=�f;<|W�<�1<*+{���I�Z�<�Ȟ<�J���=4}���<��B=��]<���<�����N�F�C��<�<�k��ytO�����SB=�6�����U�G�C���l=�˘�X�λ�$A==`r��N�F�4�'<[�\�׫e���~�uF��V�xf���6=�q(�r�Ǽ�9�<=T]�_�)<fD���J=�J=4[���<�呼`	�<bzM������)�sa�<T�M�3�F��Fɼ��ͼ��G=���h��<�׀��nq=�M�h���&�^=dƸ��iż��;���%7�<Xj=l��_?=��k=��$�fO��SL<)m-�������$�<]AW�Ӌ�;�.7=��d=�ż��<f*Z=���k�xѬ;E|���<��';o�_��<N3�=r�9�۷7<��W�0�=���<�� ��Ƽ����C=�:��:��:6��j<%����@<��=f	��")=�2Y��m��jp=�s�¢<��.=nRȼ�,=}3��˷<yq����<�=:�D
=a��m��?j��X����f=�!��h�<kc=[������N�q�<2��<@E����<\�==�v.<�46=�i< �<b�<�r�<�;��9/�)�=�W�G{Ļ��w=�p=��/�4r?;JA�~�v=���
_j�J=�]�*�y<�uA�9�<�4��xA��)����x<��=�O�k��<�8�a�=�F<�����<x�S<�#�:��<�$��<�oV�G6d<� �<��U����;��+=%����=ܼDU~�&"=Ii�<�0�<��}=S5<��ʻ�l�
~G<��&�L-�;�i�������;6R;�n<������'�K=/�&�vo<��=��u�A1=�C=j%�<�:=Ǚ�Ktv�2e�<Ƽ�S^g��o:����;��<-y�;��=��P=*�<�{=�/���J�<��=3TS��Ā<�U2�55�<nGȼ�y<4B޼��>:�Y)=\S�<��=E={��<���<�(�8y@�<��=�=Â1=�pX�qm�< ����^��Β�_�*�%ְ�X1�!��<��]R�<ꪴ<����D>�<�Q9='R8<�U<�ڬ<D�K����2�V���6���(��􀽔_H<��H�n==���;�c����;��4�� �C�V�gg���<n���}=��>;cʭ<b��<*'?=T2Q�P6�<���s�C�vX^�\�ռ��9l=���<���<讣<ĳ=Z�����=F@�<^�&�-~�<�ؿ<���W�$���y�C�]�9E=�	�<9a�;�"p</�=bo�;/��6@Y�̶C=h�A<C��&}�&�8

=�(=G�<zc=��0��L��h=+=`���{D;�宼�6�'�p<_���y�ֺ�#���t<=I]<�2�:�4<<5=%�S<����a��`�2�~:�d�ۼ����?=�ET=&S�1!��Y2�=��<��]��ջ�:�<��t���s�W�<��t�v��<�D=�"N=�ҍ<����r=)�1=A��<�^���=]=�I<�P=/ݼk���6M=�Ϗ�S��$:��NN�_�h=������'�I<�IS=�����:�9��v=}�;K<#=\]��<����J���9���;�1�#=jY\=pĩ�B�=��=z7��ٖ�=�dP=~��<Tg��3�;�-;C�0��>�<+�3���T< �o����M�)D�<ol�<�#;=�o;�=�y�ݼ 󽼃$^<Z�'�U=VX���=L�ּgB=�sJ=�M?���*=��<F =X���I�@���u�6��NY=�w����'���������w�G�ـE=!����k�;^q�<�?��0=|H$�b:<�N�<)�!=9=E<�=<l)���@���dzF�ӡ��g�<�g�=+8�U~V=�[���<�W�u�]�&�=_R=�:Q����<Q�=I7=;h��<(y=Tr=(��=������'b�;0݄��^h==~ݼ�y<=N��.<o_S��0<n�v=Z�_<����4=� L:q4;���%=�E��</1>�ϼ�zﻖ��<�Tļ�>�����ְT�|_m;F��<rE=z6L=i�X=!I�'Ճ��Lk<�?�z	�<�jռ�y5�Ka����޻6]��u��<:��;�#��\��<�E\<��)�E++==dt�X��<���<\���:_q=N,����c(%<W�Z��7e��ȼϡ����Q=3�<?M1��C=���:�>T��j鋼p'j��sO=�pP����b@=��<�lR<t$79�{<�N
��8�qa��6��<���/U=s !��p���=��󻀕=[�/�Ƥe=,����J���	H�B�����}<�-<Ŝ=�=���ޙ�<UR=l��^4����<4�<�uL<��]�G*R=�
�<����V=c,c=�o=�-T�s�<B�M��*�<aWh=�ϼyA�<cH<"4M��Ef��u�<>�M<Jͻ��<���<�l�<�X�<Y��<��*=��M<���<x$�:x
-=�4�N�;�2;)� =���(*�@�*=�C���t���w�;�W��{��=+��;��<�/�<�f-���<�L:�;9&��RǼ��`=���-�<ö���Y<�b=��ϻ|ی�P`��W�<����KG=��!��`=��+�u�4�|u[<m=K��0/�/�:��.������"�(�p��P�U�<~(�<�ݴ�J�F=t�=wm9�?=E=�������G�-\<����"��;{	�cK.=V;�=y|�<�ɷ���<�P�<��"��Ё=��:�=�o���_�u�	�m���=�߅<v��/�ջ��V=Fxw=��5��;-F=8#=����k�<b��N2A<!�;�܌���<��<�i
=���<�eT�:��\�Z=��1<���<AwF�xļ��#=a�:���<���<F\�<����F<$x%�?{��_K�<�=I�����;�ݶ<iY��;=�H�<��dr<��*�v��$M.=ӀH��q
���<��A=V����<0�<l�1�T� �)��<RWc��Gh=�=�jX�E�#=pD>=��d=��<;��-�z�}<p�Y�|��;% =��F�'�`��e�<�z#=�k6��˼���1=jЃ=?��< B��a���O:#��<q��<?0=1����<8�g/p<@�=��o����<�{�<��Լe B�Pɔ���<n����l� �2�����p5<�a���M=c�<ϢK����Ym�[��<�mb<d8ʼ0�����<cQ�<��=p��<\}=f���� ��<���� =��b<�D
�����=�>�ԧD;ruH=ټ�]���q=��R=���S<7��=�b<��=9�=�Sg���Ҽ�f2��/=�=�p�<�˼��;;BsG=�}�<D�q<p�5�:�<�]=Ư<��&��bN<'r\��hR=s��<e�j���֊��U�<�e��z3�9����<@���W<3���d�󼒄�R�=|��<�Wv=���*��bX���7<=�졼�<��=�$=��	��T��<��I�������a=!����J���8�}�Z=�mмQ�)�D
�J^*�}��:Y$)�`e]=I��<j�<3�.�J#��PV=21[�"�<�B)<}��<M�2=���<��=t��&q<�3�+|e=V�Y�T:<f?="<�Z=�1=�9��3�w=Ӹ1=��Z�ώe=���T�3=	eV=z�<t�=��ؼ+ ����ۼ"��<�����=v����O��^�x�G�L޼F+W=¸ ==�<P�C��Y�<��<9�H=�P<��5�o��;�q�����<V�)=�<��].N<�}�<=�	:9��0��`e=ng\�-k��������=�^=�`��=��"=����E|�<��9��I=�弾���8�=?U�<3��;�,ͼvk=�{(=i+ּL¼��ϻo�0=!�X=o9�ǣ�<!�����<_��k/=������7=f����̟��;�}+�������#<>{����<�Y=�fD��{�R� =���<i�3��aX;���c~�K��ծ�<ވ����{�;k����3���:=���
B<@.�,�����<��N���=�¼&k7�vZ%<��f�Ӂ���D�;.�N�ϸ�<��t��=�`�=� �^Ҽ.��P"�<��P�q�����&�< �R=�S}�z����=Ǫ�<s�:=nx7={�;�r�<W2��T���7�<��<-;�9{>=3Q6=>����E*'=H�i�^�G@����<�X4��n�<$z;�/F�l+�ȟ%=���;��=jW����o=�jT����ՙ�<��<�>�;�N�<DDO�@4�<󧐼��x�<N��j�<}3�<7���"�Z<�T��k�:�Ƽ7ż��j���a���T=z$�T=l���y*=�AU=�����<0�<�H==�̼�j/=��K=���;$ ����ݼ���"KK�o�6��5�ۓ><V����q�< ����/n���!=#�<s��<�"��KRK��ἢ��<hм�<�����<E�x�k=�Z=�	=<=͐Ｑ�<���<Y=i;"���<<���<�n�<�#ɼ�34=�U�b>)=���< �3�!A���\�;3��;"�<���<aCO��>�=R$=� B���v=��Y����Xa׼*m��p<�����c<Yw�< N���p<�E�9��R=}��<�`<*�^=ۼ<���@!��y���4�C�1��߯�.ּ��=Ĵ��d1`=�/������)�0���,=�ua�w�<����,<�Xx<�0��V=�S�<�i*=��/�m `���!=��:�a]='Q.=�ռf�=�K:4/.=���� W=X���m룼�7��M�<* �7��Z=�y$<��*=]��; �u=+�k2=S���e<��{<��z<���<��<"y=k�뼁!�>0�<8b=���<6�h<O;$�|��<�Jn<��<'��oK!���;=e%<!m=L.=�Y^�o>/=�=�^U=��8=p:s=�f<��<\V<@(��2"�����|����9��<t��<!N�^����<��컶��;צ�f�c=���<�\'=YA|�Ҫ�<Z�+:D�F=�^1=\�<Y�:�?��d�ż��?=�qZ�T�*=��<bHh�����z�Vi������g���f���ν`=;"7�L7=`"(<Ox=��;G�=.)R=S�f=X=8=Dj���7� �,=�@h�7ɢ;��,���A��\p�x�I=K0W=ђ���+1A��w=q^��M</��<k���U�
����<���<���<��=nt���=�E��Gڤ;��=�}���ʻ(�<=�>�1�Q<��ى;|��-�%�==a�;�؂�;�=�Ҭ=�	��6<��/��1Z<��a=�b��6*��`=E4Ҽ�c��0�<��M�И�<�aU=G �;��=@C�<�K����<B�<m7m=-&
=§t=�M<��T�%:��[_<G*t=��Iy�6���ۼAA�;��=g8#=�,<Gx�;�5=���=�\%�w�.���?�ӼbS���;=~N=㤶<1���$I+�Nئ;�OL��=��K�6�O�f͑�r\�<�� =�W�<-�:��!=�Oh�����`�$����/=ڝ��h����y=V�:�R]=�(!�_�=%���Y�zQ=[ES�0���O:��<��=��<�_-��>��K=�=0���$�<Α=��<����T�;���%�<�f��!Z\����<S�ɼ�?=Z.�4��;���<���<٪=;��e�ݺM=�f��L�<"�e=��1��,�7/,=�.=Ȭ��e)#=WNM���Z�9��h���=���<���+���)=���<�H�;��N�ڌ�SÄ<j]=Я�;���<˖�;�ik�����X�<��"=Ԧ�;ԣ�<f걺���<��h���=�5�<:=;�<gò��X7�dP����ݼ�F�<�c����<��S�������pK�<w�:���*$;�yY=۪5=/�Ի���<�請�z)=M�+=��<��=�q��u���
=8�p����3|=Z�=��P=7��-���h:�LE=*�.=�*�_%z=K=4r��!���b;F)@<>� ���9�}� ��J�<5�1=�<Vb;<�㼃��<];G`����<ݍ�;4T"�_�W��a!=笥�`;=Or>�=�J�Z<;��,<	_f<��S��Ҁ�ĕ?=B�R��;=\iv��?=�4+=0*K=�.�K��<K
T=&C$��*ǼO����X�=�6�
!}< o^=ޅ�<�Gx���^��ٲ<,��<�=�0�l=�_=��<SP���+=
c���}}<�="E��t���H
<Yu�:a�b=���Oo�B��;����o���D=ɞ�tj�;E�n<sWt=����q��c@=�! ��/=������%��gP<��<��==�T�s�2�,�<�p&y��X���G���]��@;=�?;=�։;�=�JŻ�8;v�Z�vռ<��7=ںX=|�J���$=1�`�%�;����w~�=��<WV�bZĻ%-�<�S��sB���A<x�y��<8X=Z�.=:ռ�H�>w�2K"���f><2�<�ea�l˩�����ܻ�-|<��V�X<��
=5G�:����a�<��<�45���e�t=��Z<�N�}�
�m�7=�;{�|�%�����+S?=R����a={=�5A<j�/�^�4��N��o?��=[=�7��
x8|�n�ӆ<@=�v��I@?=�M=�]�?�i=}k =bb\<j��=�M==jԺ�}�=s"K;,q��P���'��;K�U��!<��h=P�
={�����_<8:���<���;���Di���u��Ѽ�'/=�O��^=�%�<CuZ=����T;==�-�;:�M�0����޼����.=��A���A��Bh�m*P�P6��ç��hIm��c_=���<Ś�<��d�8C=Z;]= ��k�B=�$�Ⴤ�`K+�I�
=J��<iT;-|&=�1���]��2Q=�����ϼ;�(=gw3���~<:��=�ke�0^��")=h�׼����.�}u���޼�< Y)�9V�S�s<3ȼs�<��=PW!=���j�k�3�d;����1�<=(�<-�&��1�Π����<�)��
��@�R=0�1qW=.F�����Sh=��l�M���nC���g=Q�����ۅr<n�Ҽ�Қ����;��<�2x;�SX�KE<�%F�ċ=��7�E�=u���^=+�=�-Z�~D�ȿ��7;����B�m!�>�=nvD��P=;.	�LHK�rmE��s����<�4S�XH��/=_��<Ht!�Aw��<kup<!z!�K(W������k��&=�NỘ
=f�(�8?�������J��,׌��.���9�p5ռw݇��=@߈��ߤ<p[��ٕ�:��_=F�
���P���U<�|5�.��;
�<�ak�����O)���<�'q�����'�g��Q�5�:=�~<�<�	e=t
<����M+=��;��:=˘�<���<�<�W9<�*&���=���<�+=ȣ�;���M�:�:�H�����s��j����|;ټ��f��G���D=��^��఼��Y=`��=sF���k�W4=�2=\О<�`�`=��<x�<I�\�n���2�t<�,�<�]_�$��<��V<Ue <�w�p�4=��\=�ƍ;���;���,d(�b!0�0�	��,��0�c����sۻ����»AJ=Roغ��k=���<P�Լ�]�<GԹ�����u�#�7<�!,<�<�#�VL!�����!r=���>4=Y�x"<��T=����o=�P�<��,=�=���X=o[��R��T�6=�ӆ;
up=٧e�3&����<u���
��Y�\=�\��;3�t�<[I�O����<���<�6�c�N�x���q��&@��� =�<����_�Z�"=� u;)�=ԗ�<�+���3��t<�a<9rf=��=��<+=��l7�;���o���=�}m=]q�!!=��p}U<���<�P.��
��0w=��g�iu0�B��<wBS=�F`=HV<�T0=L��<p{O<�hp=D�M=�:?:��r�=�}�<l�X;�+="��X��>�<��̼�Q�=�C<��<��<���;y<m�1=i���Ԟ;g놽���<*A׼c8M�ELܻN��<������;��I��we��x<
`=(��<oi���?���/;���<�
@=mvs<�<K��б<K$� �B=��.<v��<Nx,;���<�d�<�R�G����-�� ���쩼�*=r>=�&A�����x*=���0V���]=ߜ�<�9�<��<�,��܁;',m��]~�Z[=��<1�Z=�2`=����B��<�;��=h��<\&F=�*=F��=="b��<Ծ���-��<�x��g �@��l7<�۰�D5S=�b���Ƽ�Vb��{��<4� =5�<@['�̫޼�w��}L
�xW��㣘<6�?�=�"=��<�ּw��_}����=R*=䴟<�d^�9�7�_s������?�sY׼�U�<f�=͹�;���<�?��qټ���4^n�갹�q���'=�����Oļ2����� ��^-ڼ���j�;��Z�j=J�=��'�=gJ4��_Ҽ��K���ֻ1�<9t	�E�;�����F��+'=\=pN�<Q������^�<�yͼ�#=�<D�<�.m���L=�k�w��_�%=�I���b�<1jI=�( ��i��2�\=ޞ���=�L�;�n0�7~A=�9�=G�-=�
 =��<\f�ɻ,=y�ȼ>L�a�Ȼ���<{�.=<l�a'=���<^�g<��=��+��Ȅ<�ZJ���A�K�c�_a��X�'���#=�`=R"t��e����;������<=���<o�i�Uo�:[����<Va<�=id�;��I<p����<��==�t��|=��S=�bR=�H����=<˝</u�0�4=����`�<���:�_=�pC�lȂ��J���R=��?=&6���T��ک�u�|�1��<Ԫ�28q�1m ��EF=�D=g�ܼd=��<�����i*=�੼�Y�;�\��ؠ��iN��_��3�<z�X��Y�R=����]N\���B=�j=�
=W��`,�<������7=�S����<�qΩ��֌<� (=�?�<��d2�f�:=�G=�@���I�<�+�"d$=�bq<L�U�9��<Hn^�u��;Y��;�"��9=%�<�>1��N}������+�"�k�d��V=f��p�U<^1=3�ȼ_zZ��1��q=�<ÕH�4R�;�-�<�=^�H��d�KH���I<(8H��A=�G<sy�s[�<!=ֻ�xD�ٲ�i&s���U��#=P<�=r��
�e�$=��;  <ױ$����<�W�k̘<6��<�T�/����c= 7�9G�	:�h=9�0=�$�<C�<^�a��0`��4�/�)=?� =���ɼ�;���<��=[p�X2�;�I69��<H�;�"-�<$Q�%��<6�%=.5�;Bt<2;�<]ԼiJ<��p�̼�;��4s=��!=
�K�(	м����+� =lJi:#6����<��J<��2=�u	=W|��5�p<{����n=�#A�s��r�Z=�]=$��<o���p� ��<H;y��a�6=f���I�ּ�ʶ<�z=[��<&x*=v4��Ke<�+��=�[�<,S=�&A��A=IP=Hb;|�<�w��;=�>�<|����`�;t�����e�a�@�DU��P�<�.=A�<�4=�u!������RE��'�<��,=2c7=DO��v2�<K�,=�^����м�H9��|*���-��%9;���_�<.sL�KNP<���dO�<�#¼�=�3�<d���*C<��H=��D=���s�ӻ�x1=�����R(�0�3�	&����i�٠û������g�}<��E������ƅ<�c�<jn%���Y=��ۼ��N�H��<�Hż���<*<�<m;����+=��<�Ɛ<�J2=�����?츂�\�t5S�R2�<��=�L�T��;P�;�l+��7�����<g9|�>57�s�˼V���:�p�;[�N=-If��X7�xZ=��q=����:E=�1�W�P��f=��Y�<��=�+9���#=nѣ<9��<� m�j=�=$M4��0:�XS<���i�<���PU�;�K�����RG6��\�:,<$��<�rO���=�I�=�\F�*4d=���������7���<)4��xE=����Y<==4�<��=<�7�y�q=�[���������9!��=���;����q(���:����o; ��<f_�����<��T�3�����=�yT<���,=���<���;,p=��A�h�F��/X=� >=|��E���d�<�Z��D%��C����=|�<�F�u��<3�ּ��B=���}i=v$�����7���~ ������
�(�;ww<�}��D���M@:��0�W�(�x�=ʬ0=k�B*��5���^tE���<:�~=���(^�?M�v�R�����.)=��$�
�.=F�<�͉<�	�<��9Q14=W�=hrA=��)=Ũ��e>=�;z='�j��r�<���k�<9�=m��;R���-<��<�ɼ�3=Yc�U�,��0�<��8=��é��Lg����<𢼨!����<��7=��q�5��< _q=&�F�<����\�/׊;��=	�<=�\���m=��$=�o��~�"�։¼x>=ۼ�E�=�I�u�G�J�<��3:-һ<G�w;K�'=�ta�Gj�<j�<�Uk;�r[�y�j;��,�򒉻�� �7}==M���F=+&!�x�<Fe'=�{P=jP,��ٻc^=*�d`=mm=�g4��S��R3���?<�<�0<p6�O\���7��r*�ho��Ez=&�=C�5='��<�Ja<9�P=G��<%y=N=�,L=�[t�>�P�y=/1H�Dmz<��A<�*<q��<���<3=���;���<�X�0�}��7m��2�;<�&<%Y�<��h�P�J�9e=ָ��U}	=��D<�{"=�fͼۆ|���>��º<��ᤨ��}�<��-�wV�<!�=��J��7J)=r] �u������ވ�<o� =k1+=��=�;�<�B�<}�;A�B=�<���~<hJ
=r�����=Pz<|[.��A�YE>���(��*�٭(�,]F=7w׼�n[=�<�J<F#=w]i=6��<5�x=�7#��RF�������?	�!��=�?=}!��t=����R<I=�<ә�<nT<��C=�s�<{�<�}ZP=��)<IYL��]%���i���b�h��<F��<��<=�-�<6J���.�Z�R<<�j=�4g=B�=�n�</���\K�<�c�b�D���J=�>%<��a<BR�<I�Լ��=��^���<5��;�o�N�<�`��V�T=Z]s=��@=�JN�����; \�],��S����T��M�=�*��Z�<"��@ޠ<0�m�!b���^�>�5�.�6�0��nE��F�ʼ܉��f��-B�<25���7L<��?=����;�=����Ԋ��tp=J橼�
��ּ��<����W�v�;�d�<Na���i���n��٭�^�~��+5�� �۫�L�+=��<�P�O\�<<�)=�dE<Kɩ�ʂ���.�:���<���%���xM�ǢɻSp=F�<0C�Q=2㡼;�<@�1�B����H8���=i�����>=Q��̼=�<4�<�!�<��J��|�Nb1<����?V��r����}�)�1��� �����m=x}�<��M��O��|�<$��:a��<+s�<:n<�<9�<O �<&Ca�|�%��R<�ї�C*u�K=��/�M�ݼ�"V;]tl=�6>�*��<�7��!@;cļ[�<E�+���;�3=N5���=���<.}����y�i�=I%�<hYd���n;�-�<a��<�⁺_3=ڲb������� =����m����coh��� <��O�y��'�[�j=�]<*1R<Z��<"�*<�d»�ǀ;�\Z=)�<��9=c���:�u<H�,=6�^<�[M�6X�;�BL�'��<�+�� ;��W�<w��<���<��2�qLS=f�9�������=�(�;?�M8��K:8=�^e��H/=Y녽*��:�h��4;�+u<|�=l �<B-f�I��<^_�<Y�����:A�<{���W��(�<Ӗ<�g� ��<��0��9:���!�<���<�>_=[�==�Q ����,<Ҍ������<��1�3-=�����z=��i=�Մ�jʼ&�L�OV�<�7���(���=��P=Z�P��߂<#�»V�к9��B��S&�<}~<��=��<�V8=}��<��+<ɥ;=���;�����=�԰:�� =gQ=�a?=���<�r<�6=Sx�;�c_���="д���M;*G/=�����=���b�^�@/��e=��j<��ٻL��<�]|<#<�Ƿ���<wp-=��T��r=��"�) 2��|廼�H=$ʓ�a4�;�Ƈ�a5X�ش��_�<0Ѽ�0	=��<��"=!P�<�O��>}��P<6=���b�.���<��=j�=�>��}߼�e�;q�8�Vy>=�,(�t�<���<����W���M=��=<��9� �<��4���U=n�%=��мTtB<�j=��<�rQ=�Մ=��7<���<��i��j9=b��<��<b��<��2;c���	�Gޅ=�dC�G��"�<y�%��ᙼ�#J�t�'�{/�<�[�=M�h<}Q9�U�<\�<�o=�S�-Ib�r�r<�%���5��+�=�<��<@w��jW�<��K=����HμKT<1Qu=F��d��<ܺm���3<�7"=�L?��L'=m�<��ۼ�*�<wzo<���<l =���<Xh���瑽�U8���<r��KH���(=;)X���A�V�;#�Ƽ�B�<�&Q=���<|�	=�$3�p�<S=�w=�3P���I�O�<�(T�Ks7�M�c����<��9=,�4*W='�7���u=/�<S�<���<�N�;n���.!	�L�0=��	���=��/=��8<���<���<?-9=__=���=&�ԼK>�1'�<2N�=�ON�x��$6j��p��<��<=��q=y�>=���<QDA=!�-��Y���`���c���=�H�<]�����<�s6=��=t!���Q=�/<1g�����PY�<���<3���<�<���q�N=�{P=<(�<�y�<�X#=S�=�K�<0L���B��W</$c��!<�i��7��<�@ļ8a�<��;�T=[L�<�vj�<q=\�<�!=i컼���;�u�5=9n�9c>=��"⼈C;�y:�9�-b��K����
�e��<B_1=4O����<զS=�d-=�'�:T��8S=�'�2� =jkR=��=���߽<��5<�8�e���%�e�7=I�:=�_Z�
�@���\;@�<=[+�<k�=��s<t�<��<�7��z�t�3�>�8 ��C `��3�;�<.=�'�  �<?�\�UOR�+EN=N�5���mxE=S���ZK�W4� D�<75=��m��<KW�<��\=?><,,�G�n���!=4V7=?x;~<�
 =fN��J�����~��H�<��I=�q�~o�����<Rs4=����UۼN�C<[�N��"�F��Q^9`g��a�f=)�7���C=K��qK�=	Q=�co�'66=�s;W�]�(!9�H����9�o��MB�<���;�\����=`�<:_,���;��g���8=�����<M���5�%#�<�i=7_B���EA����#����<v=� X=.)�9)�<n�I=�RH�H��<a��<�������<(��ە)<�໼+� ;ɹ�<��A�IW=����1=T4=5K޼= &���1���R=��8=���;\ϵ��Q�<DK=��4�+��<�^=��<v8�<��M�8�V<�H�38;���=�;:=&i�bt�(����!��Rڼ�*)<�G=��4�}e=���<2�S=Y���==�w<�>ռC���(�9� �<e�K�l n�;K8��:=��<�ϼ<+K�uQ =��<���<k�u<��=�Ҕ<��=d:ͺ鼤�!=�Y����<~��<�.<?*y�����EҺ��<D=t�=ыw=S�<HVt<�X=Z:�9�o=�_=���%=�l9���V���H���<�k��-;W�=��*=X�7=�:�'�:��Q�����<?-�<F�H=[w�8l�)9��8��Q�'�-= 5=�V[��%��x'=\Gü^��<���<���,�<�Z�m:�;b2����>=2����O�N2��Y�D»�A=ട��=��5=�Eϼ(	!���l<�hż�(&=M~S<Z�1��"9=n��;���<T�Լ��޼{6o<$L��W	�B�o��a=յ��ML�#��>�y�Խ��+��<��!��H�4��<��q�<������2?=���HG=�א=��,�0м�W���S�>j��h��/�;=8�<���<�<$I��@g=���<�
�<�3B<�_=�D�<�kt���G=�`�<}0żt�p�����u,=�.=�����<�@ּ������=L�T=���"=�໿��|~��#K=�E'=# =C�>�6[<�͘<������Q�<���k���A<�K=� <�CƼUտ�Ь�<��:f�!�֑����v=C�8� [<��Ǽ�r=��5=4�Y=�e1=s��:[�r=��=�<�(�F<�X�a�=+�@=�;��˻�Y���=3[�:՛�<{���<wȟ�[�]<J�<�do����ڇS=���c+�<�u�#��&��;�׹>���r8=��<K�\�R�Pj����<-�j���<e[Y�M�=���)�=fA���G�<�%��#��覼��+=�?�޾A=�A=�p鼃o9���ܼ�=��<��)���=|�5=F�ݼhO!��d\=�F=�.�ބ*=_�S=�D���N<�/#�*(�����&��I��"�]�{�^<մ�<�t��<Ǎ<���<窂<=N1��4J�2�K=[�!��)=�"=������Ą��q,=�E���L=�=q�ϼ��#�Vy�<�h��=��)<s�R=۳P�$�[<���|��OP =��:��L=��<*=e�<�J[��
;�V���2�<�ʨ;=铼okc�%�W;?]2=!@ļD�L�C�;��m<�M�Hq�縼ʞ�~W��0|�< ��;P$���@���o<�9�#�S=��%�M#=�9=��=�Bw�M�(=8a@=%N�:�Z��+(�g�����<��=�ؠ��8I=ᬣ��?==䬘�:F�&��S�<e׻�Dw<j6�=G�B�`b =f�Q�q��<�t<ȳ��w�P�;����/=��;R�ʼֺ<�Hv<0P7=�Tz�0%+=lp�<b7���0��S�;}\
=B� =�0;l^c=KX�<��1=�yG��Z=&"=jf�;�<Ʌ��)��=�<d3�¹���<�YH=�:�<:%��<P� =�e�<:8=Ӟ:;�=Ƽ�|��컼[+d�d���;m�P��%H�w�<t�2=�
�:�o�<�̼�:�C��<i�P�Ueӻ{�V=C8<B��R��+��	2=HoK;��X=*χ<h
߼}��<z��<�"��,?=��<]HE���*�	2=��M=�h�Un��4�b�\���"�<���/<��b��WZ=i��^�/=
9�; V_=��<$Hݼ�����Y=JG����<���<|�R=K���t<a�H=�d�<�켦c׻PX߼޵�<-<TQ4=5����3$� �1<�]=������7=�|<w��Y@ ;��<<�,��4��<���;���:�f;��=��;�Aj:w�v����7.�<aL�7H�(^=&l��	�<ԃ)<X�E����=c��iW:�{#�͹9��<q���i�[t������5I<N�ڻ��K<b�n�P�񼽅�P�l:�F����Z
���!���W=�M_=�`�<�V���cR�i����@�p{ؼh�(�X@7�;��O���P��6$e��s�<db�<"4�<��5�5G9=��U���<i������K�c���΍<\D�;Jh�<^�S=ǦN=;_=��<F�<�S�<3?��h�<a4�<��:��%=mV= ��<�\'=2'<ш<�8��R8ļ5a=����*`><��=q�&=�;�A<Ƥ&�G��S==���<�3���:<�����Ꮌy���p�</S��g=��^=VNP�f��O���K�!=��,=��８�=���<^R=h=�f���;C�=��;�w=Zʆ�� ����S�j��<�a�@�T<=H�４�����4����Ҽ��%��8=�L;���<�A�<���1j=~#��2z�����g�]
���9�a����W� �i0�<�ޤ��=�<��;b)��8�Į�<��;=���<������ ���_=9�B��K�����B=̖0;�W�7�:/�t=Xü�.=a��;��<�TԼd񢻓�o=��z�3�.�u�/��pX�V<w<��,��{Z���D�"*��~n?=j��]����e,<�p�<%K��+�<!�L;XBX�K��B`л�xq=5�9�*p��{�7������9�a	�Sm���B��}=��>=J�i<bS=�P����;M&��Ĩ<)��;l.<#<^ܵ���&�*C3�"(=�����ܼa�=d�|<&=P6�����J����:@c=�麞a���XC�0<P=�����<�G�<��=�3:=�U��@�I�Q���)�/�k��Ӟ<D-v�� �<� �<�&y�=��;Td�=�� �1�j<�B|=��<�J�<�<w:ּ�Ƽ��5���ܼ2.�.OC���K=�,�"�u��(=p�!���<�W=�	��<�Oq��>>=���<[�9=0J	<r=c�T '�_Q�M�����<F�����@=U^=!(1�s�T���y��fS�)����a;���E=�c���d����6�=92˼��.=t��<�Df�d5,=��<7���<�5�tAW�6�%<�*d�*�ݺѹ�<5s=�(��V��s^���=g�l�#I< ��=���:ο��`��<5$�� =57D�K� �?�; zڻ�-+=�o=ś��V}]�zn����k��愽���U=�V���
�<�o�<Q~=��9��={!�p`=1�<�?=* =�[9�'֍<�p��> �8Z�,<c�d��4�$�/��=z��C�����<�y���;�'���<X��</�;lۜ<�k=Vs ��.=�	8��������E�I=f�5�I�5������������ۼ��j�H=`ۊ�UH-=��+�G��:.=�@�V �<^P=%%=j��_��`�����<��=)� <�0=�}<l��=�O�:u�b��M�}�<��=3s<�O= �ܹ�-M��B������<R3�9g�H`<X�!=2&T=�Ii=�L@<��<QYO�l��;��<Z�Y<n�	�qt9���zn�Yu��n���J�$-?��C���z�Yg�!��G�K=��0���<��3=l3G=��l�&�f<�T�܂s��1��w�<v��<h,�6���g1��u��F|=,=-Eݼ
R>=cU��ak=��3=;O��;(=DW=r<O3�<�v���|��pݼ�f��<��7���a�=,q��U��p�;ϑ9="V0=/Iټ�<=E퉼�6�<�Yɼka�@��<B�=ޑ��������ר=�a���M0�
=�<"e]<��<<��� ������H]=��;Q�=E=��"�q,=-��y2��N=��<.Sh�pb�=���A�6��^-=A6�2d�<�X.;	,��]=��h��Z����x=Gj�;��)=�%M�I�<v(��yl>�Z�=d����=��ͼ��==��K�	�P;éw��<eC�<OT���A3�1�%�$�;ZA5=8�d�g�1��� =D]�<�f�<�i=5_)=f/ ��i=�&};�\�+���U�<˿żV����x@��w�gY����:�<�M=�f黐:�K�;�8:�6���C�®��2�< �=7M�<E<=���q�'��=��l��|��A=�4=Wtʻ��<�T)=f�s����;��;pu=Ё?<��=���;^5g�����<�X=aI���j<5m=:͂�̀C�8�-�I�L=�',<�9��:�|�<���(�<%�<iy�0LϼC�<�=�(U=��.=��� �����W=�9=7���L�h��6�<�������2Z=6��<�-���*꺤��e/���U��6�V�_k�=w�KVU=�(����<�.�����K�B���N^<E<�<���[A=�%�<4E���D<&�N=O�����:�c<��H�������[�݋=~��=�.=g�ݼ�Q3�F��<
#!=��B���;�`X�\s�<��A���)��_�=��=:���s2=1����P<,��Մ<f<N�
����.y��Hp�V$0�g�<�j�:$�ͼ~�¼��<�����<þʼ��A��2���S�\$�<��<ԥF���=!�1=s�=%�T�9+|<J�~����;;]+<�Y=�7=O�y�:!�|{�;x��<e!#�un�<ٻe�n<���gR=�	��]�<��C�^�N<_�����;�	=�=
�Ļ�9<D +�i^1=��})=�h!=�WI��ӽ�<p=��~�����&=��<_�<����<';＞� ����<&j�<��K��<��L<����<N!D;�B�<����.�_ה�.==��K��;>�p�ȱ��)�$=��z=��!��o*�>(=�� �4�R=�-Z�
�����=���<�V+=��6���5=׻�F<�YB�X��Bgf=+t'=m�G8�<a�'��:=>�r״��E��Y�;����=M|=^��o�]��<�?���K=��P���k�ȦU������r'��������<��¼��A<�h伝cb=�)�5���`=��S��;=-�3=�<�=�%=�g�ΜS��]ֻ_�N=�l-:��ʏ��Q1��
W<~��<�L=$I�<h�����T�G�<�_=�����j<�Gd�ޭB='.��dS�so����	<}�]���\Y3���f;��3���<��x;�6�<R�<��	n�<1�ռP�	���GHJ��
�:�=�:D�3��]@A�C�=�F��t
���A=�Ɔ<3�;]砼U5=
��</;A7F<ۯ����'��=r!}�Mp�H�̼0A;b:� T��C#��_��ME�<���������<v��թ-�8��<|˼@^L=A�= no=�,=��{<屍<+�a�=������Yd`<���<R�+;�H3������>���;0�.�`��� =d{�<P�9=�=��H;��=�W��l<K�=�d<�1�L�����<`���*�<r}�<���<zD+<���<L�	=z�C<�|);��a<���C����Wx�+~b=0QA�)�x�3R������żh�0��<�^�=L��:<�&�:�\(=�EF=(��<+?��f=��(<��<4�x<�qͻ��n=z�<x���u�}���͘�+T.��,\=G��g2.����<M!<U�,�k敽 �::���<�����B=��p=��H�ͨF;!�=w�<=��; �5������z	������.;���,<���<$bT=��>�p9� ^�H����A�X�<#r��aq3=��[���^����<jI9��S���D=�j=�d�����<��
��u;��^���5�2� =�G=�Ze=3����8�+<�><q���	�<����2����+��<=�����D=�缸�8=;�=F��<��F=]�b<0$��>=0Ǧ;)�=*�J��0%<�����=�r= ����<�|��cf�"yA��l�G)Ļ�P<X2Ӽ�%
<����5�t����(=��9�^&�;����]�;g�9�	�=�2=`#�;����ĭ|=�m8=6cp��dF<]�.���k=�k=�B�: �?=��f=�[�a?&����<�O��h{��R�0���*�G^V�mv<>�l<�[P�̩��:�<�<�(���lj�i��nZS=c#Y����Ks=R㲼��K=4�Q�q�=�.�q 7�:�3=d�@�7�G��h��3�d�m���)<�7H<�� =F$�p��'�]���H=�����n=W�=9`�<,���p�7����;H�<,�����;�ϼ��<rf=z=�� �����M{j�O����=cf=���<K0=.|F�M�C�f=uΈ�M��<?�2�����n�伂�?��A	=M�C�l��K��<��߻}�w=UK<j�7��-[9�V�#z�<ח�Mk8������B�<���:��U�.��zx;�+=��J��1�;O`=4�"=�K=G�ռH�<3�v=w׻�<K����=� ,=�m�;TEI=bj\��**�n�.=[Jg=�ā=�����9μ�1��P��|=�����\
ڻ|�3=L�j=�]��:=�Z=�1�<�"2<�����7=K�}�����=��"�'�=��<���X����*#=����<��B�<Z��<2x�; h=6��<N����÷��:�Ì$=R̼Kܓ<=C�<�@�:�ӌ;<=�9���C=��BV��ϟ���=1��w�F��-�<QJ���^Ҽ<B���7$�(�[=�NC�X�r<T�=�����2��
˻�>=ϕ�(��(.��c�<j�&���<�߾<�
=$�;���<o?�=fmg�N(ڼ�!�PTO=M�X=��+=��:���+��9=s�ɼq�<�Qo=1V=�G�< q�<��x;��*=)�׼�=��m<�jZ��v	=m��N^k�S�#�l�<���f%=ӫZ�ˌa<6��<=o�<u�+=�9B�.�J=
_=�P7=��Vd���<�eG��2=4U�;6=@�μ�+1=_9*�!=�6�FU[���>+T��X���N/��̹���)=��U���B������Y<3hY��X����<�C�<��X��2,�9��<��><��.�@?=�󚼂7��Zv�����޼sq7��2f���;w�5={�<�����A�<�#=@=�j�<����V��|�<|=�;o���L�noP<Qļ��q��49=Y�̰�<��=���<�β<��W<�KU�	�< -���~<M!��8;=D͜<3`=#\��t��;� =�b!=�K����� T =�1"<��I֩<��o<�]=ߥI=���<S`*=#'M=4*N�1��;�b�<)�A;_�2��Ț��
h���=�t:;�����r"=��W=r�=iX���߼7��50;��=�"Q��0�<��0���휐<��i�8=n ,=�Z��I=�� =��W=��=��<�z�W���.a�<��9�*�<#���Z9=$�;^ȼ֣<�,�<*��<2%=1��gGټۉi�Q�h�7�kA�����s��>6�-��<��]3m<��=�1[=l�n��k��(vR=C��;>�C=C���ߨ�<�r6=�8�<C*�ćO=@��<���<�sw����_���&Eg=|�)�
FԼG�;q`=;l2=�_I=PG��1�;�\��_>=j$�	Z*���c��#�t�ɼ�������Ǳ�Te�b4=��S=�</�n=@S}��ԩ;݅�K����=E�� ��!���;�#i<e'f=[%�<Y��;��L�y3ټ����O*�g��h��=�ݬ;6<�<���
)�{8�<�2�R}<� <�$R�����8�5=���<�z;�'=�dR��1=���M:�ե<�26�,��<猸���<�t?�A?�;����=�4?��μc�U���=�%K=�#�<-�߼װ=ӂb=V�B;).=ӛP�8"u��v{=7?�˕���M�=[�<�\���$<Ѫ<�FF�*Wp=������Z�k�G��i:<�n=�z=��[;�>L=�z(=��u�h�8=�ӿ<���$�,��T;ǝ�<['�<V�y=;��;ϥ�{�j����<G8�9�w1�yT.<	~=�
���.���[�K�B�-����%=��+=uv�< ���=�=O�w@=q���=/=<;S=PH]<�PD�`A=<1ټ�j,�ą�<-�2��Z<*��<�L=�#|��_0=4��;�:3�%�c=�V�<P*��2�&(==�;#k;G=.���OS��d4=��	=��U�<��y=�Y=Q��=F)=G��U�S�9��<�������<u��;$ϼl�=�',<������=��&�������&������ �/�<f����=Y<=?�={��<;(�����+4;B�c=��=�μ��4<	�<��%=ĩ���/�3�%=�G��(N?=n��<�=�GH;�3��|<?�=�3u=��-=|}����K<�A�}2z<���E h= ��AV�<3�<��<�@�=$l�R?�q=7L=��(���Z<��0<�`= }y9��<�B=�Em=�v��^_=A�v=E��<�'9��`=M��Ö!��$==�"1��Y =A��;�j�n�Y��޼��;=f`>=1C���<蜼�h�=�I$�ޏ����!�=��,�U>J����<�DU��t����<L���Wj� ?=��<O����L��}��]�<�:���K=_\m=��A=�(9<gw=��������)��ܘ�<��y;MP�R=��!�n=��d=��ļ��<�)>Y�w	�;���?3<����톼7�����#=Z�*=H��<`�h�<]W=���<Ĺc�"=�20�~jc=I�f�&j8��y=E����\̼|�.�&��"�g<2�(�X�<�����[=E���#</Rw���컁_=5�=���$����>=�����q��ۊ<�e_@��==C��<��ϼ�
��Vs<���9�<y=xj6���;=0	 �8A��[����@~<�
=��<�λ�Ye=AW=�U����==ntڼ�"�H�];pGC���Q�T��W����ʯ<b�@<e;��F'<�y���$�9k	=�:=p��^m�O�ȦU�{~�;X[�p4�<��p<������D��S�O���,�<=�_����Q��<ܮϼ�Gz=��C���<񙃽K;,�\S:���< ���0�=7e���_��U<-邽��;β_=ב
�x�$���@;�3=e0�)G=[� �I���"��]���(�K�J?�<��5��V��7G=�&r�w&���l
=X#^=��=�q�䈈�gG<��w;�b�0��;��4=MZ�<����=����Ƨi<ZE ��0���<�����G�`'&�.D�;�)���=*������þ;�	�<��f��JL�X�{<�0�<�<�L�<囝;d�|<��<@�d=:�$���T=30%�����U=��<�2��.6��Dl�\+����h<U�R<�x仒8==a��<9��:M\X�YQP<�A=��E<��c��^C=��/���e�ƺz�={G@= I�<]E�<�}���Ҷ�;���<S��=]�ݼ��[=A5<O�-<UJ#�W5:���E��KS�i<=kx�k���]�g= �$��	��#�V=Jzp;�i-�kr�;bl�<����#����;�y���E��v�<{��9�L�<��"=���,�Ȇ��䲻2΍��;�<ZmH=�=i����B��NX=��#=�s��sC���<��)<� �'2C=3䰼��F<d�ü�=00e���b<<�<x9}�s1�=�m
\=��˼�漯N���(<���<د�="�<�-�r<J��b=� =;�b;a`�_Rt�!p�<�aͼ (i�*�$<��+�����V<�-��K���<�$ؼ79�;K�<��=��0=+M�<Ԋ�<��I=8�@�R��|#t=_(�<�=�<M��<�"̼��U�(?<W?/��,R=�ڱ<��<Q��]ѼѰI�#����V��r[��#3����YV����غ����l�<S�ݻ���`�i�;d�߂�=1l��j��<��Y=����/b=�D��2����
�7&�kPM=j�1�0�X<$�ؼ��4�p������\�l�չS��@h=P����:=��v�]Rj�)B�<�c9��s=5����뱼��<�I�=�<%�0=�~�uj=jw=��ڼct5����M�箎�y�<&�={`��5%=�܊�xE=
��:w�#=��<1��=dT<�w=�v4A=\z�<��=FI<g�<ֈ�=�����>μeg^;єr����:�/=*ص<�� �(�W<.r0=b��;�=�d��N� �����<"s=XQ�=|[R=�r�<��$=��=��<a��<mF=�c	<��$���q�<5\�8�<��3�"��<�D�P�=��z��`<�?��9�q$H<M�5<�f輙;=�Z�q�q���I��X�<W�;��(<p�s=	E=r�2=�"�<V�j�bV\����<'���({=���<Л�<h�.=j�;� �k}�<g�=	���n�>��>&<�I_<¶ɺ�:�����Y�<�&���rQ=(������<l���'�׼i�
O�;�?N=�6�g��<z��<")Ӽ�~�H��<A[=�5C=���<z!=�-����<F��ќ�<�<�1"~�p!W=��9���<D�r=(%=-V��=z�X�N�u�'�L:��I�Y�+=�r��h` =�+�r&C=cZ	���U�_����=��5�Z߱��!K==d2�m8�l�=��=���a���Ǽ,���p��ݎ�<m�=���t<��<]��F��9�-�u�Լ�������=�l��=��<�<�y׼��$=n���V�[Z=���:���c<O)༤PX��FC���|<70�;�x��w���<�>.��I� om<
��;N�L�m�Ί�HI%�DYغ��W<���^���O�<���<M(�;)�,�V��X�C���>=A�k��;{�̼)�,=�EY�*M�;B�X��_��j<k����=������s������C����<��n=�|m=�\=�fE��Tc<߮[�9X<s�;�)��'�4=� *=[n�<G�U=Ͽ�<"���ѻ�={;�<��f�D�u��AU���[�w�ϼ�7�<;�<H�<��<�ˎ<�|���m��0�ӻ,��<�G���U=*b���#;��}<O����<	��;LA=N!W��f<ٯ��4|\=�H<()��%@��!��;"<�&�<��o=�eL��(�=c�i<�?���h��P3�=�L=��y<J�<�O=��"<ǈZ<i˼�w*���=�j��A�G<b����<��yϼ�-?=]���F�<û�+-=?=�����᫼�D=:�2=� =��="xռ�J �> ��R�J��<{�=<6�-=6P��9x��?�ͼc杼�|=}�n�X��=`�T=���p�\=��=���ー{�q=a�W=����<=,,_�vXq=F�9=�B<��>�M�<�;�����q� ;भ<��*�C�o=v��m��U�i<�<<���;V�)=A1�=#�F���<e����{$�q �~�;�<z����t�v=ML=��<b�e��t<�|P�
#'=��<��Q=��!�3
m���<�����=���<�^�;�RI�b�p;'d�<R#'���A��<�F ="ٙ�{�;��N�y�W���N=<���֓=gN�;:t�<l�����<��a<ޞ�;|��=����9�=j��<�b<[Dż?刽U.*=�Hh=��<u�J��B<�t��� ��N���p�<�����`��q�a��<o��s��<�(?��Bz����L<��=˹O��7]=m�<x�Y�B.��Y:�<�����_�<��B=oc]��A���%�����{�;ϻ=�y=�7;D{A<e|=�M(=aH:��=��?������O�<=�
=�8��{j�L�~�ּ���Í]=��o=�rW=�Aػ+���
=�S�=F��;�)�<mF��Ν6��a=]ib<m�q��P�����<��8=V�����<�.�%�b=�Q=)�<DQ6�A�(�}߼�n����I =��<w�ۼb��;ko8���ʼ�|�&�Ѽ��,���3�84#=�>	=�A��֥���e����k�\���K����x=�v�;v�;6�b�w[=)Xy�p$7=���a�<DIw<O�l�����y*A<��_��j���3H�:�,=�����*�s =��=-M8=3���ݜq��?��C8�W��:�`�<�ʼ?��<̰3=�'=������e=L}=;�D��P
=���;a�=87=S�=�x=/��<�=x�b��ԕ���G��Yۼ�ҙ��`�'� ��V�<ԼK�݀���H<Q�w�Q��;{)��IB�������ɼ��N�Ƞ�����D<�'�����<�G�<|<E=��<�Xg�@��֟�<�Zx<`�K=]�<� �<���E����G�}�:���c;h�l�s~�91�/=aS��Ժb!=m��=�<����f==H�ӼR�ֻBO�<V�1=(�=5�̼���`s��� ���)-^:�ƍ<+�.=�B���b��j9����d��7K���I�m�{=̛�����A�1�`� ����3��Po�oM+=���\u=���N�j��`�rQp��e5<��!�D��BB��	�2=>�:�	P<�^=�Ἓ�J��Q�<��*=ӿ=Y��ٞ��Y�p��<S��<^KX=�	b���<M���|N=)��<R=O��<8A�����[�=X����	?����ܰ<F��+0��;<�$»��+=������<M�p��`��&�<��0=�H�<��F�-�N�H�"<�=;8aT��dO�P;�<K�%=` R=�5G���L=�f�z�D<1�=���<�h=���;�t��>�c�}�<I��<9#�	���8*ܻnyV=o>F�6�O��8���J����<"�<�=�C��T8=8e������L<��ѻ�Ř��b�;f*���:=����ے����R�={+$=]���5=ۖ�;=Id����T��j1=n-=z�T���ݼ��3������S=a|��y�<F�0����<w١���g<��=i]P=�j���ؑ;��F=AI<�� ;n8*<��^<��u�#>I=��;:ׯ���Cl��a=*A<�f�s�#�L=7rE�e9w�g�`��� ��c7�R*<�h�<�=��ռ�%���k�&�9�i�K�L���=��q<����+��y�<��<��8��4��v<�s��O�<�x�`�R�^�1��G뼨>���l��zn=�h�:�N<��̼f:�;Ȏ?�����/� �)�ϼgvj<F����+�٘=�c=
�=K2'= PW=�
�<��<��|$�X ׼�e8=9a5=n=X=^������=�/ռ�&=+M ;�b���<����<�u�����<�ἒM�=��I��k���Z<�=Yd,=�� �
�An9�0��l|�;mJ=�ܝ�7^���Q=�8k<{~Y<<6&��(J�"	�B{h���V=��J�%�;�!Ƽ�)b�*��^��=�&G�;����yߺ�f����=e�Z�'�j���s��]	=᥼5�V��j�� v�<� �<p��!�C���<<2�=�đ������Û����=���<# 5����;�Q:=�`�u�ûZ�O<*�:�9�=�W=�=0�>3�<����9<�A.�&6<%��c�<~t����3=��y��M���[<�h=�|���B|<,�C<����L������(��0��=#�U�������ކ<W|���u<������!
'�@�V�Y�v�Q�.=L�M��E�<��;���<����C��<#_�<��;���<����u,�"R�<��ɻ�u���=�dL����<�q�V�=�g%�U���7W�<�`=J�;�<�2�=��	�Ń�)��=`�`=WT�<7g^���T��
���P<���;)�.�X=�="=1n��Y����<�ڗ<����J��cZ�L�3�2�<2�P=뙻Ԋ�<��J�Pm!<뇪<'�����=��+�ؐ=�S
<UN=��ٻ�H{��S �\)�<Isc<T����B=I�k����P�;(�����.��D,
=����z�r�[��˼���<̴��m#<�~���C�<��4����2��<�#1=�{���Pt�M�<,�3<ˏ�<�2R����T�<��<�R���U<��;=�����xz漊"=W��<o�q}�¶���^��O�����(�<R��z'=�E����<4u��Wp���]=�Y1�}h-=[Ɔ��?�;86h=�]f=.w�F;=vor=�@2���|<F�����h�A�=����]�=��*��0�Ǎ=?��<pi��a�)��[E�Ø�<�A3�XT=d�+��'<���<9\�;�<*M���rr��� W=B�Ѽ�B�����(�����S���}<�@ʼ�#4=�a;f�c�4�`��fL<��ȼ�jC�`��;:|[;g�f�Z�'��V�:k_�<'����O)�z���xm8<*ԁ�V4�;�=�G<>|�1ソ��߼�v�<3L=�u=��`=��Г��i =�̼:2��Β<��H����vU=�M�<k}=�� [��<�d�<aN��"7=�ݼ�w�<'E����׺X�<!~�.�[=}P=�H=k�.�+G.=�����ź 8W�8�<*3λ�����ݼ��c�0��Qd=(�5��/K=��= 0�<?��F��;� �Ԉg=#���5g=S��͘@�����3�<�]'=)ժ;_���i<�C=�yU�#�R=� �������<|�Y���c���>�=jx=��$=#e�y�3=���sּ�p�;���<�g�<�!���*<u���	_��/��)�<�D=�vD=�yL=d����Y�<)�=��W���f�;��5���\��و���;ݶټIP<?���o="u�::�}<�C7=:�4<%��d@ɻ#w=,!=���<�ܼ4t<�0%�vk5�8�>�RX���1h���ż>ʼ��`��7�;�{���<���2�4=��@=-�I��
w<q\�4r��2�����(yl;E7?�q�9��3��M=�$<�����	Ӽ#S_=,0f<i���M=��>=OH���<�$��ؗX=�g��"�F�����ģF=8?~�[Z<�5���t�ʍj�>M7=�\��Hٯ�L��<8�=O˺<��$� s�<S=�М<��2��WQ=�C����#�j���,��m���>�)Ff�:�#�� B���0�8(�<O`�;��<z.h�'==�Ȼ"�����<�� =��;�h=�=ӼG�]=���U�2<�_*=��<�+<D �=�2���S�_<� 5�;�+=�F2��I�(��(+=���-��<���;�,/=?1�<�e�����'�c<�q�<����@�=ҭ��\�X󏼧�g=�jS<[b��	aʼ�/������<�3=�?�����h=�V=/@W�&@r=�Tû��Q<0�Q=�;�1�<(21=��;�B'=ｏ;��	��B�<��<x� <��3<V��<�Y��[T=��'<u�"���<P�I��;��M<�<�c��0Y��1<��b=�%>=��=���<D��;��b=v�0=�L鼾*H��٩<t�P=��=�T= �=x_��P��<�������ִ��2�Y=@$���q�<O�<�7��7C�`f�h�V�_�4=�f��9����$<>K�<L��dE���j�2�\=6��6�<�]���a<��<JL�<�\��?��y8t=��^�u==h�<~�O<4�~�in�=3�=�@��T=��;����M^�J�̼��<��.=e{���k=ғ�<H0������=\�=[_���������c[���f=o�_=ھ�<�x����3=U� =��J�(=��2��ۼ�\�;��=��s7=db'����,<�)�<�/��B�żU8{<�A�<t�E=D���X)<ģ!=D�<�������<����W;_�ٺ��<�lV���=�[G=4R#��<��
=�K_��׼bX��J�=)c�wI!���=6���j"�J;ټ��;�Τ<V���?�:�ڳ<�*�>��pr=b�>=�Y����H�O���������<t�%�a7j�V�
;�
�<�S=��V<dZv<-������}
������F�O�߼.���JL������G=-�T���)��)=�Ʌ�N�<_x<ln=t70����;F�=D<;X�K�SK=�G�=+R<�������<
��������B=g��<)4��D�<q�d�$=�
��6�n����4=��<mOJ��d�<8q�M"��ԣ�:L�<c1Ǽ�aR=�
=��3.=��o<\YJ��� =
V\�X�
�N��;_b(=�Q�5g=�C�)�a���6=adQ����<��;)"<�*�'$��*<��v=�β<&kļz��<
��������,�=��,=&ܜ;�:������Ӧ��J�M�+���<�a��*�����V���?=�=�;�������%=���r�q="v<�����=��<���;紅=�C^;6�Q�y��,F��\�/X���K�</r&=�2���N�5�<��L=�#<���տ��)�I=~����c���=��C���;� @�
L\==�S����������"=��8��Ｘ���BX�c�,=j=��o=�1(=bG*=4���<��4�*Ѽľ;V���LP�����<HvP=~�6�SŜ���d<���GF������0=Օ	=���e�!<���<����#+�E�.=���O",=m{ټx�,�"���~a=S =(����ʼ��=� |�"�m=!�g��S�<�!<���<��5�_hW�.7=ۊ�=�n�<�R^=�`1�;0�R�4=�㼛0t��Aɹ$�U=F�����=K缍�A;�3R��/=����,<i��{;�<<=�=
7 <<"��A�n=��=^�R��f�8�<�c����Ǆ�&�R�d���s�<����9�X=s,�<��k<��]=��e:6�N=���<v������Y��%�� �<eY1<5���p=4��<�aH=Y&I�B�����ȕ��ox�=�G=���<�߼�b�%�����=ћ�<����6X=1�^]Q�
Z����;//�*8��¼�F=p??=��G=��=����;"T�;_����K�"��9=ŞO=���<b=A�ͼz�E��m"��Q��$ݻj5@<q�	��-��j �<�~P�V*O�x��vm��h,=Wǜ;�+f=�7=@&=�ǳ�H-=\�]��/ۼ�Z�s'@=�i��=�s=��;'Y��)]=%چ=Yj�/92��c�gL�<n-���<+�=`�ۼN�8=1I��P��<Ѷ�<�oN=�88��&�;sd=I�6=�n<��=�:=���j�=Wx=T]��Q=el�<�<�<X�;(n!���,=t��<ǋ��q��<~*G��p�8����9E=�g��$�Q���7�O�	�F��={<N�9��e��ʻP�~=���<{��:Ȝ=�����M=�����Z�<��3=�%j�ta�<�{G����<�@6�x2Q��;=���;�z���r=.W���Ҡ;Y���Ĥ;-�;R� �UF=�.b�ʚ:���9<��<�H?���<l]�.�q�K��<�($=�J�<�컢�~<�~�٧�<}�<�==,u�<��;�b<�s��7鼣��N�<Rw�;�7��()������&�2S��q=&V���:���;=�=&�/=_@M���<gV;���N���s�Q�>=��E��50=��P=��&=�"�G�5=�v��T��;���=��>���|o3���:���\<f�ּ$��Q��R�s��F�;�͉�t��;))���w��=[=����.�%�	�	X=K0��R���T�<��r������y<(����:�};=�E;�CἍ[���'=��ԻF�#= 7<~�<~�+=��<n�5�:U=O��=��<qD2;))U<�v=�>���9�����5�ռZDC;�gμ/�����A�l�@,��Ū��bJ������뇽ښL=���ݞ1=�2�<7u�ʢ	�'�<��;�h�b��:��!<Ay���=������$E�Ķ=H:��6=��<"64=���kV=�b��T*�<[m�w3J=k9.�[#f;>b���y꼑]�'ӛ��=��_�<�;*{0�۳<�}<��$={"7��ݼXqu�\�/��^����<spq=�	���;A�	��Hz�Q�}���!��]�<J�Fь�H�G=�Ƥ:��6�U?����<�O��RoS�q�<um�����<�'=��=na��D����;��L�wiٻ}�C�l�S��H?������4=JV�<��+�o���`�6���<�ڼdB�<0z<YA0=��= �<�L;��O; ��<$�-=B��<�f��ͭ��8ݼ���<E�<���\��<�&u=��;�/�;�����; /�\�]��2O��#<Z[�;��v��\�����<U�= q�C}=3=��J<L���R=^�<�,I�Г�<n =+*�<���;����==�Q=�LT��H�.�y��u׻9U4���k<&�G<�	D�����im=\�/=D��c�=�B�;�<:y'$=<�2<����TW��SO�}�0�f�(��=�b���< 2I��fM=��7��ڽ�~I����[=�G��M�Ѽ��\=S��<�k.=?<�<U_�6@�<�BG=&Qd=���-�a�����0P=�=�9�޼���<l�(�/=��<���<��;��<�:�<-?＀|9�d<<#�`��t�Y�Z�&P=��F<��r=�����S�P/=�ց�>j���R��+=��@�a =�=�Լ�h���A=ΏF=�f8����6�< Q\�?�Q<x��<er<3��@�=Y�F=��F<�x<zGt=�Ik=�{�<`��ț)��"�<L��|�N;�i�<K>��ᐰ�v�T=ȁ?=8�}u=����+=��X=�����
=��<$"ϼ-Ö<v�<��7=1K�;0>=�Ʉ���[��Z{�q�y;
�=+��<���<qO��F��I)����;��8��V� =v�B-V=1ݼ��5=c�?=z"=�F=|�L�<%�;��ở�=E�;o>V�$b�nsS�=�=�H��¹�4�<��N=��=�kA;�3a=�r�<���<�>V��B%�::`�sXD���O��=�&y���<��t�����X��MBG�*G=�lM���U�<��s�e�=Ղ��b��<�6K�#�'��� ��O��X��_=%���-M=�O<M����ἷ4��dQ�a�����?=�����=uf�;��=~X<�����55��a���f��X����<�Z�;��d=RE��Z�#�	�<J}�;
=1=�e���6��L6�Ĺ��C���8A2;�&4=�-U=����:dT[�c�l<`��;8��<�<�1��>/��-��0!�<����vC='��<�(�t�<�$N���=ކ�t0=y���N��{6��P<f�W=y`�G��Z���4=�g,���I;�ݼ_�9����<��<�X= �'���,�X�0��CL��񙹰�Q=LEH=�/;=C�<�sE������U��P�����l�ܼg��<:�=�/�<�3;<��L=��3��qg����<�p,�)'H<���˖D:`�e=@�|�Ȉ!=\����)�-=79�+��<pm�<�8v=-����B�0�:=:g�<��V�<��.=�.=�k�<m^�<�a�A¼�`�<r��<��<AB<؀}=�F����� �ļ�TA��3=T�̼��1<��"=��]=a.s��RռϽV��9��ܼ�`�PI8�As�#�a��fL=�Ǡ<��<}3=���Df+=����;96H��YQ�X�gO=P��:<Լc=�y�iB&=]ݻa���ಬ�i�A=7�#����<�I(=�G<������;S9���#=��=o�;Fx$=L��a¹�{㼫�J=&<3��<\�<X|�;U>p��T������=Q��	f���<�=`�<�[m�@B�S%=~��<K �<�I<@iK�m��7���X�<�y�<#�;�Ȍ��h���d�#�z�.��r�C�O֑:�*_���n<o6.�9�W=�:�<m�z<g�:�6�=�_D<[���kS=~��<0X=�=3�<=x|�H+�Q��<��P=�˷�^J=+1=��Ӻ��;��k���%�<O6�=6=Q�zo���l�<�g����@�i����I3\��^ =@Y$�6�<���8=�lW=��;�W\�H�=�	<��<��<Cx�<�~� ��i�u<���� =���<]x=Y�<���<�Z�͢��x���,�<'�����<sE�;�(��Ӽ�W��Dټ�e�<
�-�<��Q���=�Nb�3S���<�ީ��:�'�@����<X�1:���ۘ��=�%~=.�<+����Q�<�.��G���z=g���\�=r���d��F0<6=��+=3׼���ێ;=9
�<l�<�^=�
��B-@��T= )3=�E(=*�i<l�=
;�ŻŔ�����������~<��V="��:5���I%=�=�;Z�E�������;Y�=����N��U�� <Y��<ϱn<�B<��\��]<�0�<!B="�x=E�F<�Ɗ���< ��>ڙ<��<@-_=U�6<��@;�<��<������z��eg=#�<S-G=�w�:yO;K��<=�ż!�<�";=�|�;�9w=��_��Nj��I=����3"�~�<JY=��"���:x)�<ӟ,=j�O;�c��k������<H�t�[b<���	<�h�<�o=R�=Z�G<N$�;U�n��F׹��_����`�#��Y����24H=%#�<���<��u;B��n�<�)�;��<��+=���<���ai��(;���+������z�,=SX?;Ō��3|���j<��=ȭ�<����@���=�����1��WXJ�,SD=�ߔ����<�仩�==�GN=��z�>��<8=;��;������<p���\8��O6:.>�;�I��:	=�� <O,һÃ=� ���m]���<���<�#c����4���H�M�]`=P��<3 �� ���`<�4��<(����*(=a�j�Uż�/�:����t턽��;~����]�׬���^ =��2=����{�<ƣ�<0�<E�y��-�@�k��Ǌ;mER��K�<�ז�C���o �V!�<�F7��H^=AB��,Ѽ�8m=�=�J�&��5��<�kM�@�%=��n�@=�W=���<F\��+�<��Z<�%�9G~I=�v�S��N�ȼ ,��O���?=Xi+�L���sq;]@��wO=ĩD<b���r��"�N=�r�B�=n2B=,8�<�p�W<s ��ud=��T�A�<jol��f�:����3�<E
x��y@<a�\=e��2�����<m��;_G�(f;=kQ=��ѻ
KB=�$�<$=:�3���y�m���<f>=�ȼ�c��#�-=�:1;M�P<I�a�IP�ة�-�-<���c)D�Ӷ�<J��<�yD��=.l.��g@=��R�\�M��S=�6���$=WX�<C�=�j�D�4���=�܊<�1s��[�����d=�e �pU=�����)kr��<��<�l2�
?=�я<R�<��m��v�9����:���1=����;l�X�IQ�\/=f}?=//�<� =��z=^3^=��,���b.=�Tּ*���s= �C=��+=�;����A��V�Z-<��3�*Q6<�oB<���g���7=G�����J�k����^<�p�3�=���;��d����<��}=d��<�}��C҆��0����=/-=�O�$O=u"J=~
=�9�Ws9=S���d��Nb;���:>���Og=^T�dW=Ht���=Ӗ���bd=���<$Z�k8 =KjM���;�4,=Nq�;�7=��+<��:=�>U��Ҽ�=_��<o;^=
��<d3�:��<��ؼcr޼�M���m<r�=HF?=9+#=� d��7=S�*����<�����,1�<�Z�����5<�� ���P���\=�@r�g�U=/�9=ȴ,=��3��/)=uA�aA��0u= R��	�;�Y>���L=֋(<DM�<�U�=�*�; y�;p2�9-=d=>=V�=��vd��D�<dH�<�"�<[GY<g�=�|����c=�����i�.�����<���<[���pN<1�(��i.=mvd�)(�C�"=��p<]}=��Ѽ�Ȧ;�걻���v_��_�
�s"��=�6��\�,��9���<�q0���]=��μ���Ѱ��
� ��w�<@`j<K���o>j�t�B=�u��1��ά:��;Ac =�=��m���q=��r=
4=�o =WV=��'��<gHj����<6v�ى�=���<�ʏ=���8J��<! �<����Ӓ�A�0������b=g.*�k�T��`}<���<BL�_�y�K<�F�;���gǙ<й��v�R=<|�p={��;wDq���"�Dr2�����,�<ʕD��n;=`��{J4=ϐ�<�'�<��Ǽ#>=�:-<����P�<^a��+�5=��)���`=�N�<���
���=w)=��@=5�j�>�=�P�ĝv��������2\<��<}����=Ѻ�<%��<�,�BO�)P<�w<������M����Ϻd<" ���M�-�ʼ��T=��>���;�¿�;q�#=�=�]4=N��4��D=�2;�<� S�F@��>=��=��b=��<�n=��� �=l[�:��<�%�=�|K��v���$<�#�dڥ�w����ۻ��d���<��3=�q8<���=�V;�,j�t�ɼF���H�;�P��M��I �ta;�����G>�Ѫ=��=ik*��c��C��6�2�n<��V=��<�`=�jL�v=÷E=��7=B�I��t��g��=�d�<�K��IU<������j ��>=F��<.�����8�����8:9�V��ܼԯ��Q��\k;��,�T�T�:gI=�Ϸ���=b#�s=b�<i�X���<��9<��1�����pk��u�1��{�?=ގ����`�h0�ш$��ļRꌼM��<��޻U�?< � ��%t�N���Q�<V�j�5W=�����:�	N=g�%���Y=?�;w�(� j&�N����;�	�B$[�8I������@<�Fc��-m�-�����=�K��p���<��;l�#�sYg��T��e�~���=�8�GV=�\�q7�ꉼ���=��_;��`�$H�$�0<;cC�E+3=�(-�O%���;�@,=v�+�MK6���;�]{<���#	�<PZE�1x=���<�������������;�3w=�7|��%��	�`���['�;��_�$Z=C
v=N��=E)�;F�M��'��<uѻ�_�<�ܨ:9T��l�b<��:�(�۹�����BE�<{q��-�9<��[=�=(x�<Ǒ��r���v�����Io�</���P<o�?=˝D�+�g=Q������<�>B8_$,���<�{�����C�-�<�U�w�Z=e�A;��<W�\=a =�d<�^;B�ּ���<��&�b�<�Pa=�|�r N<]�'=���<�M�<�i=�i���=Z�u���f��0I=�O��	�qZ�<�`��	Ἦ�>=�FD=[�M�=���îջ�yG�_� =`]M=9o;Z�\�N��>=}��<GN�����R=�<����A]���k�;���<�^�;����Ğ=�80�z�=�1$�F�˺,8=����gbx�Gd=�4��_H���,<0��;�@㼋n�/H����<��z�����{�=�=�9��c�^<�<�<�sy=Zގ�ߚ���u��H*<��<�U=G��w�����<s\o��)0=���Mf�;g\ =+��Y�w=E��<��J���%��2�V�3�5����Rb�?�=(=o[B<L5ջO��=��<���<��<ӓ`9�Oʼs�<�H=�4=����l|<�܎�)�<���<�/P��n�}A=�ǳ����<� �)���>�[�3��G)����<
"V<B�M�`��:������<^弃�R�s�d����:�"Y=��El�<�R�<���;���<%O ��$`�!�=W�<2�<��<��>���<��[<M�J�$�l<�gY��{�<!�Z�h�
�O/=�e���/�A�n��D�<>�ɣ�<vh��B+��,����I%={D=g�����;��=�s���=&� �O=款<.��<����?d����,��<+ܙ<�{�;�1����I����<Y�<s2�;��n=C9D���g<�'�:���8X�<�9�ubh=�vM=���<&]L=5�i���&=�>���-:A���<"݁<c�Q=�rQ�e>�s�]=^(���g<C)J�E�3�k�� g�C���W�=`�"�a4#�̆=unI=��=dS�=#��;��#=ʧ�<=�ڼ�٫<A�<���=��:[P=P$�<�Z�<�4@=��<�D.�d�k�|`�����M:=d��z���k����;���� Y<5L=[D�Op=�3=Y`e=?����<�_=����-�6&�<�dj�ZO��N���KW�j,�<�e���%.=��<"�Z��-w;���?�:=6��;d��;6�a���Z��탽!��`��� �O=��{���p<�p|�R�=d��<��<�㙼�Vs=ߖ�<z)���m�L)��ӫ�4F>=�μ���f=��$����<�����;�).�D�@����Xa�;dԩ�ݑ��U�@=�Ԉ�[ֺ�	8�<\]n�×	<bT^<�p��. =N߼y�L=�-=��2���A�-�N=��U=^���
|<Vw;U����'�"	� KC�6�V=� =Y�S���<�s;FN=�*={���#���[�~��u/�#���yx;
�t=�����d¼�]2�X��<_f�W<b*��T�����;h�J�, i<��;����h�<�"3��g�<�R̼��;�_=Ӟ;w�̍�p��)�7=3L =��Q=�0�<�)p���=���;�c����)=�"��:�\���=����W{��ur=��=���;X*�<�����!=���JI+�����8=;��<]Y��)���<�P\���7�^�*=�O3;��&=}$=�C��\�2�B=�B�<ee��!��<�=�<%un�ʜ������{��N�;<UL���R;�n�<ܥ#=ù@=����_��<p��=c ���:�v���z�p��	�ں�F=/��f�=��v�� �g�<�1�;C�<h#�q�m<^==V.�_���-,E�"A�<ޯ�<�U=�"��㶼V%�p(V=���;}�Ǻh�� =7j~;1<\��	=���Y�������|��'=\*N�l.���=<��];�h�<������%=�Z(��~e�>8���� �����ƱD=�8)<ߘ�=f�3��j/����<.xd=s�H<F|l="�#=�0u<e�<A?�;nn>��_�<�|=��}���C=�B@�^�����;a� ��D=���8�O��ۭ��bA=%>x�z��^�<%�;�yĻF~%�j�#�0`N=��c=}��;e��M༏Գ���b�!⠻�=��*<cg=)P ��=�'���G=J��@;�<!�ͅ<M�u��"��E
= \V���a��d;�Y��
NT<��9�E�U=���Uή���V=���6=��ټ����n�0�2=3�� �¼��0���G=&X1���<lC< ջ@眼U��;r0����<4�	<sI��I7�;2 =�꠼W����� ��S�7��A<�m��ҋJ�<�j�=�=��(��8��#��<�@����%=���<HO=$"<+��<�����	�A�����S\��|k�<��O��n/���5=E(==Vd>��p�<���:a����M�� =�R�w�����#�j�b����<�=|X𻦛E��<��W���L��}�;D�x����<K�t;���<n�<�mh<{�:<�R)�{�=ݏ�����v�<�K��	4���yf��I�����<r���7�<<�P<3z���.���伪��<�Vk�M���!]=�.;�tr=��4����<�Q(���D��v�;�<��-���U�>=벰:!�?=�ꤼ�Ҽ>b�2d��t=�y<���)��w���B��F���"�����eB�eQH=�J��D5�c�M<�|O��أ<4-�;7�<ˈ*=�_S�[�>��<����S�<=a���n�W�����0��;��a�C��N=�8=W�J��#�<-n��_�<:�	�ʚ=�{���\ �Ŷ�p�Y��Q�;�wּ�\<��n=��v=��<�**=�v4=b) ����<�@�qa�<���N�&<�iǻ���h�Լƣ;��=�S��!�=�=9c_H��_�d(���sP=��g=�"�<�I<ڗ�9��B<����6��<C']=��.!K�hW=�b'<��x�����ܚ��y�;ڢ(=�F��2<t="��<�!?=��T=�~=�����@�<��n�
i�� ���Jϼ5�R�,���+ ��������=�X6=j�<��<��&�M7;H��;a�=���<�.=�h���v<!j�oj�7�b=iZe� :׻�JP=^���	����� :|�9G�z�*lK�D�j�s�<8�]��ڪ�PmS�8�"��0J=��<�2�;ȝB����;���J&=_�*=�̇�D/���E)=;<@ �M4=Cf=�ݼ��?Ӈ:�x6�L?���q��4�_>i=�MY�<��:�4<��i�2�l=��9==�'<;�<�<0�L<�c=�Fj:�vb=a���P�/=_�9=���9�k<�V��-=��Y_�<��O�@V����<��D���: ^�;}1=Ń==ٱ��g1�<s�=ɹk��{b������<]�;�?i�;ٯR=T�:�i=�F�c�<i�:�����	=S���C=� :� [�r@s=D�=�2K=�A��z=.b�(�Ii�v)=�%1�q�Q=�2����W=��<��E���;Ƽȗ_�v��:W<�ӼP=Z����=#{�;�rh;=��<�{��n�<�Җ;gR~=��<�� �� =54
����;����6�E=�B��Vrn=���<3.���?<�����0�YPƼۮ<�j���!o�r�T�d'w��-��#�$�<-%�;��
��ʼR[3=��U�A#�w��<�ol=n� ���W<O�<���;����ܶ��j��;I<���v�G<($;#����j���a<�!(�%��gn�����X/=�"�<�3)=�S�+h
=Sf=^����3�S�e=?b;��r�A�`=���<�����^�<.X]=�ٶ;�;�<��=�cA�Z�<�PA<l�(<^�,��%A;��S=��O���ƻ۳�<[?=	vG=�e����(-r<!Hm�L: <��L�)=��O=���:�	=Is�<cC����<��X=;���̒�m9�<�}9�dQ=���r��<3�u;4=�\�:�y�=W�ɻ ��<C�=�7=IH;-Y��X
;�[���}<P#P�Nw�9�e�<L���U�{<��<��*���	�0�z<�r/���Ｂ�R<>���O�����^=^̤�V��`^���h=ƃ�<�[C�)f=y�"= �=j��<�o=Ec��|�=�끻�v<f�h�M�r��rE��Ѽ�;�K#�$ջ<(0=�'�:f=�'N��=��<W�U=@��:��+<��<���<�xk=�,+�¢`:\c¼��<��=�4�=����7����N=Ak��2�Lb�<�����=ӹ<¬A=��2��	�Ғh<���>Wm�Wy�<��I=�f���e=j�,=�%�<�k���-R���~=�N��sm<��=ӑ=B�L=��=#ջ#{Ӽ����,t=4�a�$�=�{���<A~?�6ꪼ/8=�۩�@��<?\L�M&�<;9?�v8���g�i��<�;.��<�=�[��a��Sz�����}<�v�:��j��|R=�T�<r=ŧֻ;�]���=v�R=p�<����b�[&��8�<A+,;��"��I^��K =?�=��=ϧ��F-�=`�;���3\2�G�;Ǆ��F:�v��<R����~������DH����<��;��%�5��x��<��<;~�Y65�V�<F+�<���l<�$;ɉ��7�lY5=Bu�<j�;ʫ"<��?�ݲ��}=������<;��<:]�L�=�)��=*�5<2����G=�8��������<�6D;E�;��^�%�x=Ձ�ey�<��u=�I�{���4�<�/f=�G�<'�[<WܼIY=T�>=�0�:�?;2SF=.��;ZP=���<f=HR�<��z��<� =='�K��	r=�o"=�%��D=�*:=:l�:J��)|b�ӹU<P��<������E=� � 5���:=��f�i
J�<�~=��B<�8�wn��2�=�<~�%=9����ļ,�;��~<��a=�3����|�%���;�x�;ď<���M��<`�<��==H��9��j=�S�}�:=�����o0=&�L=��#�&w���Ġ;Jj#=Gl̼��J=Ф�<Z��C� ���<���<�a=\�;�
���5P�lnR<�>==ⅼUp�<�Wr��ʼ���<�jy<�y�\�A=�<��u�<��)=�D�q���١ȼ ��;���Aݽ��z��\u���<[�F���Y=�Ǫ�N+�L|E<�g=,<L=���<nE<�9M�<B<�m,=-7"=PAJ��bټ��컀R=i~�lT�ͨ���$=ͺ<q߄�sXH���/�`D�{���Y4��M=���W��Q>��j#0=��A:���=J�D��F�<�fH;|_����\��+�<���;
6�wwI;���<W�2�d|;��+��	���W{�:�<�!��)��<��F�����2���(�<<��;8���<��=Q�M=
w$��Ϛ;�D*������_�h���6�8�^�<]d<�!:�>w��I��<Q�����d��B,<8B��7�N���:���>�S=? �:P<�����<<� =?8b=�%���=�j&���&=�Tڼ�b�<=���eB5=��D=b�j�<�$�;�/���<�P:=L��=�D=��'��S�;(�)�]׊���a��=�L�<x�<��<�
��sD�R\�<e<��J伣�?���O�(XF������?�m�L��1H=Y�4�^S��=�`<�B�9n��<�L�<�틼�N=�;�KQ��uZ=Tsn�m��<q�w;�>��XrQ�h����Q�3z%=�1�=T�<(��=�!�=sEԼ�=��<��<����F��U�ƒK���B�#���(�=�T�U�;v����W��V/<��<���'��9y�L�ܼ���;3��]˶���<�[7�T�Q<�B���2�<�n=K�X<�BW=�X��&E����o=HI�<��9�B�*��M7��n=�{\��he=tq{<{����==&��)C��c���L~��E+<V�<��~=�n��v��gl����F<~��<I��;�p��I��8;E�� �(��;D=:ml��m��70?�|�i��5=���߭�<�[ �BD<5�=	�4���y����<�3���-u��C���=������$=��-�t=�� =�oW� K��pU5=�c@<w9=uc�<�5(�Sj=�Z'=���z�!�����͋�;���<eX3=T&�`=>��:��4��S���VJ<�źq��<Jg=K�
�|W=��<@��<���<�yk���@�N3���g"���d�����B=�$3�i+�<F!g�W���?�Cl����� ��|���De�<�:߻^�
=�Q�;�=����4��������r�<J*�<��;��R�G�\=����쪼=Q̼��f;�R� ���~'�Z�8�����<*�˘B<��k=�g�<�D^��#��b���A=�(�V�r��TQ�\q���T��T�d�
[�<�l��k�=�)��z;�<EZ�����;�7��6<(X�;�Xk=��.��O�<y�e�I��<�۷;X�<��/���<\'"={2=D^<��;ou�<�x���C�h̚�a�d�^�K��$b׼C4=���[��<�е<�*=^G��Y�<{����B9�%3���� J��UI<��";I�<Fe�5w�<U��<v��<{m��+ż��Y��$#=�I=�<�k�WZ/���<���;��<Ov=;$Z�&\���=��td=�	�3z��%�<rW�<��(=��A=;p<��H7.=&=�v�=���<�ap;��l=��F�69
�������<W5�=���<r9T��`%=,��<�I�;����_L������0H=�6��h)���ݼe5r���d=x殼W('�/G�<�P�=���<���<p0�bsd�G���<%=g�9�-o7�Y�T=�U=��˼5K ���Q�t�'��D@=?���vL<�/��Q9����ZdW��4<��P�4��<!�&=b�)Y�<��:�D�;�)�]�/� �2��4��|X<M�!�䢑��9^=�d޻!a�4���R�]�t�<32S��<�Q��8w%��P,<���n�=�b4�gQ���
=��^�9T���c�<&��<gr�a7\�'��<Ǝa�a�<E(O��=�H,=�C�<�.�<�'&���<E�M=#�<J��<��<��I=#m�;�׶<V8M��%������D=��;G{��52���<��D;4�gK����<$�<T<�<h�i<��<0;��<�Nm<r��<���"�����=	�ռM/ڻ�e=��ڼ�O=z��<�莽=~E<�z�<';���+�<����s�<�N-����:R�c��<�0L=G��<�_���<�H=��T��Z�<�]=y��<�P=��=�离��<xu���<���<�4=R��;��<a>���/:�)<4�0��<�<��,����½����P��-�	=ѳg=/`=���<�>x;D�Լ������;�$K<��E���1=[�@=�:���i�8a_<6��}���=�`;�����<s�=��(�2�>�U�9="�|;��!=�c��o=���<�g��s>h�%�)�4Խ:�V��{3k<hq< �<J���+:0�;�<�����=ٙF<p�\=s9�I
�� �<�j�<�x�<I�B=g)�d7O���2=�K=�!�_�=n%��>|n�&29=Oڈ�-f���#��+ɺ@g6��yb��t=�=�^��=��p�,=F�b;y�>�__�:������E����;2��{��[���=��-<l��h����߉<�&��z6<��;c]����a=��=����;go����$;;��;5<���Y�^�@��?t���μ I=��$����:�rϻ��I����m^��b9Q=C�=�[��G�,�UF
��8V���= t�<�!�J� �V��L�<�(��m�<��ἬV.�~���<�t��S|�;K�ļwЦ�6�#��v�<苃�Iڼ�j=U�!�jdλn1�<e݅;h�=���;fO=��?<TT%�
���f���[<q�O=d�=ov3=|l;�/j<q�l<(��<Gü1�}<o��>��<�|.�w+=�f� D��D�={���h^�����ڼ�H#=uk ����D={�:���E�M=t�<��O=�O=6�_=�ӎ=��a=�.˼�D������#�u@�!�<��Ӽ9�6=��<uC�;��<=�!=��;+<�;����$���>1��~w�<	�:��V�U�c=��ؼ�| =K�D=�.=�m,��39<cS�Z>�<>L=�Ǽԁ%��	=�#	=�M�;k��;D�#�N�c<F�2=�H�G/��([=�=��U=B�K�+BǼ��a��Ӽ�z���E��BB=��<I��=u	��<#��RL���=��C�?�]�A%�<b�C=8D�<ǋK��S���d�'�T=�%��TvӼ"�H=�d���o��ݢ��	��;�'��r1�
�6��n:Qƅ���7=㕩��=�*=R	 ���<S�=�4弤�l8�(Ӽ:^�<�S�;��;�򻾂l��b=��>=���Y�%=̆D9�(ӻ�c��2�����T�IM=����;p�D���=�}�<�6=�Lm�j=)<=&ŧ<5�M=�R�<R&�<�t�:?�<�мݒS��B�<��/=�@<���;	�<Xb_�e2=���:�ѽ<t����3=��O=�ؼ�ɼ�F�b�m7}:�Z[=�=��E=�;�QY���X�\�D�R�ż*L!�,wD=�/<���<���<T�_�ԝF��琻�q�<��D=W�Ѽ}9M�jv<KU�<����Ɇ��(=+N�/�!�c�$\��
4�K1@=ie��vc���2;�.o���g=^Z;Q�;<�ς��*꼧��<4���2I?�f�pͣ<It黡`?���V=R=#=@*8��7=�C=<z �4�K=���X��<`Z��':0=#�Լ��=<>A��89�FBT��➽�;A.��<�,������< ��<Wv==O"�<�!=�E�9a���9��=a�����)�!=y�<K�a=�D,=�v���^_=���<�'�c��<�;@��]*�)��<�t���i򻆮G�k�<��F�`=�	���ƻ�YԺ��˼�{"<%N�\�)�=�"һ�r������ρ<��<L���X�
Z:=�<�\�Z�,2��T<�\g;�-�<3E������BaO���[�H�=c����<H3����<��;)�<��=ɴ
=CqY�?�h��`<� �����ŋʻ� =\����jh=#�e<��=�=4��<�ʨ<!0�S���=j=��'<<}W��y,�d�>��f����\=j�=�e�:�<Ȅ�&7I��`�<n�t�nx�<?��<�<��&�DF=#��
��=U�i=��N��?��W�7=z�k�Ml���޼��`=|Z<�1q�E@=�2<M0��K=;y���FV�Q3=k�9=m�м#\=Q;�<�p��Y��9,�	�����==P�v=`Ӹ��x��-9<G=�Ν<�+R���=�>�<�\?��@�<�,�9��6=�O׼8,'=�I�u�)=�X�'/<��5=��=�G��߬�:)���M<�8=�7���=��1�<��V=�����<PJ���iH<�}��k�<��<L�E=U=��<A'!=4�E��E�;���:pK�<��`�4c=@h`=T�E�V��?�<!�>��.����<wgc�T���^<ˍ�>ͭ�+f6=Z���K��ޣ�<H�<@#�A�<�R�ܼ�Z�8�,=��N��`�-g���C�I��*������<�n=%�=v'"= �u=�I�w|�;w�&= L��-7<�̼��d3����;�yo�\���ݯ<Y�.�o=�Ё=�<������ƹ�?�<�P�:�M
�e��<͔�;�~7��3�ک>�����_��D=�䠺w��<�꼱u=ty-=��F��6u<-�*���*��Y�:j��=�=�_=0�SH�<Vyr�m���=N���ʡ��aH*�9w|��))��7����u�,A=���<p=<]s=�h�iS1=DJY=���Oa�He���R��Ej<���<P�;`�*;�`4�f�-���_=)R�<@VU=�_ż�ܻJ�#=/��Ԟ�<��<`�=�B��5�<]+;c�F<��6<�nT=�,���:<۴<>�Ż��-�=\��Bm�<A={�o<K2�P�:��F<�%�<=�=�9�<)� �B��<�rm<��<Z�<'��;s�]=)�<^�="�i=	�:=���<��E�"Lټ���4�<��<�>P=|�H=&�t�dBY�1h�je.���H=J�
�z�]�����g&=�M�<�[,��<�K�Nxл�����;u=�)�<��¼�NN;�q<G.����=_�<����`��%�\=CZ.�}�t��<�6=����B�*=���7i��L=qL"=
�U<���< Nݼa���zy=l��@���%;��_��R=��M<������R��^�<C7=���<X�5�=�2�;���`$=�� ��ye��a��=��<�;I<����=*�K=d3��v%=�it=�B�<��<%��<}3��V��N���ż����,=`�9;i ���M��u�0����E==��9������=�㯼u==��;[G}=�8���ZK��Q�=$����<���<��̼�9s���_����C�K�K�= u��J��l���E=��;Y��;�@(=�O=��2=�ü�V0�J2?��zU=V`t���A��GU=����һ��R=�u@<���<"������=����F.�::w�\��<�4�<��&Ho�ܖ�<,W#�o��<��@=�����H<�[�g+T=:G.=֧.��!�o��g@=ea<4��<�#Q=��<U��;M���z`���$��I��1'=.5=	=%Q<%2!=(e���A=�)<NYP��;�dW�?m?<հ��Dg���:/��<�=^J��$��[	=I~E<)�{<Wx=�O��m<��y.�s�=��:=��)�j^y�z/����h�=��=w����+<�}e��I �9PV��Ρ��������<5��<��;Y��+C�������< 72=�0�8�e�H�=5�1;���<lY������	=(���:��<��7�Zn =aH4�4q�<�0�=��<��h��<�Q��j�[D�('3=[A:=���<ZSK=����y=��=�5���(�7@K=��5=�!��YO<<�n=�ְ��w�<��Y�zH��]@�>�T;�g!=?C"<�����|6=�l<�lD=��<��K����Q���(����X���<��Z=(�(���O</�\=��,=g����3{��`�x"R=���<]�_<H�0=Ö��>e�<�A�=B�=��<.Hj=�CE���=g�w<��1�P!��B];L�<���=��{��'=��/����<k�<�LB��{�<*�7=^�g=�k�<��o��5����G����<�n�<Ϳ����C�1�=�E��h)��\�&67�Z�M<7�<��{��e?=�*��T��Mt8�^\n=��G<��?��J=�Ĩ��~:
�=<��������4�g㼂��<(�=[0m<���;a�<a[\<t@�K=@=�I=�%�*�{=Oxd���<�j;�q����\�XD96�Q��<��<�CI=�� �iK=�{�z���S�)=��v=-z<	�3=��F=�oG<A�,=Io>�iMW�Ф@������=̛�<qdD;Od[={��;9<��;s��<=��<p~V=w���0Z7�F�8�^�U��!=�r�;��i��;��	�޸r�?= =at���_�<j��w��Ѝ<�O�;/�/��<��=O�==K��<r�=�%��U���%<H���y�i����<y=|������`��u�r���=�ͼ.�s<��$���<��j<tE=��<��d<7�i=kۡ<�����G=.��<ū�7#�.�<j�&��B=�/��^�����ټH*��,�D�0>���8<:뇼\�<��i<N1q<?4�<y��b#v�g.=��O=�7f���ټ������a`�:ûV;������r�`���ȶ�B�O=��S��x��ɼ y���J�"9�<����q^��Mf�jް<��A�-��;'�}�-�B�	��<��ר��'>7=�A����;v{o<Ф��+�D��:X�{�󼞖�=�!,W��cM=N��<h�;�A���>�;R/=U1=������X���i���Tp<?f��򀽵�F���V=������;�7;8=@<ΰ=��O=x��5W���¼�j�;x� =aص<��6=M�==YY����<�ly��q���?!=�=אH=�s)=:}%������ϼZ�5<b�v����NG=�U=�ƾ<�mC:�c�<;dh��8<k �<Lm���K=�;�+ۼ��<m'�JLü�Si����d�=��.=)Y�:��M��u��:��!k=�}ɻ�-=A[A=Q�ż� o��X��"���H=��O�V=ʕ6��N����c��<�6=���<��C�<�s�J��;W�c=��t= E=k�=̐=TZ������n�����&=��N�n�8=��8��b�;���m:L�K6�<��<�h<�m���';�*V<�&�<�?n���<U��\�c=:܍����<!�'�XP<����R<����D��gN�8���1`��!'=K*=�`�KN�(P\�,�<�<g���<���<o�%���z���C=͋C<ζ8���h<���<�S<�=P�8��@�;�L��[b<�%�<��H=����n�#�Fr#=�����V=��M<|HZ=�of���J<	qJ=17=N Z���x�����- �3
=y%K���'<g܅<�ʩ<ώy<�9�	^5;��1�;��ۼO�&�_��<�[�;nm�(L����t�L��<yT=�[7=��= ����?��h�5�|;rp<=h�=�X=6"�h�Ƽ �=�[G������E��p=��#�Z	8<��f=��=���<`7Ѽ�uF=s�ļ��:��=�<�')�b�)�O�M=ޯ�;���<�o�;�z�Z���'2�	82��v~<2��'�=/�B=(N�<L;�ʯV��7�X�'��Њ=�<�=�0�<lջ<=C1B��eռܱ$����9}2(=�/^=d 8�Ft<�<<F�<k;��;ؿ<BnZ=`b;��֏��o��B8=�XU=+�v��E=��@=-�=����uO�_tM<Q3=�k��;?\=M0<ga=��'���0����MC�<}:��{ۻ�=�(;�?=����-�m���˼� T=�L��|T�}�b^G=�h<㮨�5SI�����"��*=��ң=�5r<W[��6 ���6���<H�6=�<l���$��;=�(�==/bD����;�{=�w�<���8���<A���"��H� �wS)=[��<y�=7^=O��<��;=�[�<��=�c�NRf���=��	<��e=$/���TM���< &v��1��<:=�|=B�o�/n���=}��<�:e<<�d=��6=TՇ:�k�<�d<ˁ���h���=-O=Z�'�W�V�$O3= nԼ-�J�5�<|�S=+�w<{|�x���<��;��Ӽ}�=�=�n�*g�<��<�!b<��
���W�7n�<�;`�=/�6���<�=�;58E��A&="�c���^<7`�N��b�):��=��D<�<x���(C<��[=s�!=+�6=U?�]\k��.��<PѸ�@�T�tj;�$W���=9U��)ü��<�I,=M_����Z=��$����t@=ع~�4�:�"�;bx�<N-=#�9��<�<V�0�I#=�� ��j4=���<�+�JL< ���&Ѽ�mռ�I=	������;3ռ���ʶ$��p��sAn=�ɱ:�v-�ɻ^�Z�ļ
�=7x���&ͼ&%f���j���<?��<ZQҼ-2��g�U�;/=��=�%�<��; ���͛�J/=��<g�<��P���1�9@=8�`=�
�����<Ś�����;�^h=*�A=�e=��h������2�C=zQ[<�x9<}�Q:��I�q��=�_���8S��>{=��<��;}�g<��*= �G��~򼀳�<����W!�2DS����<�p<�t��p�+=�o��Ŕ��=*=��ȼ��<HTZ=�H��<��<��=O�˨<�R<0Ie<�O�"g�<ڢG�"-�ɥ(=T���~�=�6�B9��,�������Z�<�u#<i��<�U`��Eϼ'�i��?a=�.�7_�;Zfg<�l�NxG��OW=�,?�B�G��DR��-'=7-����k=�� ���4<r�<�)�M�� �Wf���.=K鼖s����s=��m=)m�1}X�ر <���3�sL=! ]=��S�G=(@=�)����6��(7=Z-�τ
��T��`�?=Ų�<.C=(��<�Y#=k��Ù<��ʼa�G�Y����W�p��<ȿc=c�]�CN<�c<60&=�ȧ<\(-=��.�i6� W4��}�i�>��Uq<�n��=T_h=	����L��J<���=+�<=����T8=���=���;�Z8���6� �D�B���F=���<��,<hOF���V���<={��|�!�/U-�z��;5"I�Wѯ<�{:���8���=>�^=4s<�<=nor�=P��0u;k�4�a=��%<D�(<�/=ϟ���rB;�B*=��A��������u�N�S!�ƶܹ���<�q��# ]�_*<��)i\<J9o<�Ax=�*p�Q	��2�=�#W=�W(<u�Q��Z<�읻lV_=��<R�=g!�GQB�e=�(�i]><�(̼J�϶�<���;~�3=���Z<�=S�=��@�t�$�� =�ؚ�;J�<\����?6D��b����;��=�5�;"���W`���V=�_x��su<�3U=`�>=���<&:����Щ�m�:�:�)�<�Ձ=�7�8�(=��=Y�%��6��xX�?�ټt_���׼��f���&�����R@�<���6�V=��=�-<E���u:�<	-�<�*�<�����EGn�M+=����u~��'*=�8���
=��F�xG˻��5�ZL�ҏD�w�c=
 ��0
=�*��y8��^H�<�5�<z&���o*<+$<�h;5pK�]�Ѽ��QZM=�µI==L=�+-�	�-=yEܼ��
=Ν=��h<��B�(F9�������׻\�<��Լ�����_��7�<��=�K<���:G���h�g=f=j�:��ⅼ��˻
r@=_�*��N�NM2=��r��.<�D�<u���&�<,23=�)<ɮ@���6�@.�< �黠$�E�<=0p	=(�=�i;I��=��*=n�E<-	�<��4<E��<i��<�����;�{��K�<��G�z"=�p�<�9&=nl��ZL�s�ļ��='��<�j=G53=M����b=�櫼��p�]�"�U��<C�M�K~R=�C<yhf��,<\��<�Qk��s��]���4<� 7=0Q3=�o�Kr=���<b_;t�=
�̼�g�]�����;�xG�@YE�.�ۻܖ��.�G�"2=b�=��{<j�Z������3�<�����n�m�<��m�5ZA��j=Mi��dK�]��<��%?�`1H��s�<��2=�9c:�e<=��=�y�:vb%=��=T��<��;=3����'�h��=��=�
��/��0)�;ct=T �<2޷�^a=��N=��_:��ܼ\&���=e�j��:�/<�A=�ꍼ�B)�6�*=_]~�V<?=~�v��\=eau<��<�-�����;�N��t��fJ=�<=p-L�(���m����:��=��O=Qyz�W����k���8�^"=]=����D8<�_=�1c:��D=�ꇽ�wF���ѻ�<<�WF�p�J��˹���U=^�0���;Ԍ��!la���D�t��,ǆ����<j�N��=�%=��9��=�����<R�����<;�=p;��M�=�k=E,�;;=�d��2�V�0���n=)Q2<����ټּ">�Q�b�d���Z���f����c<�]�<��n�-=�챼w��<�"J�~==���<.�<�2���O=��`=}�"��5�;;v�<�/�Ƈ����9�� ]�>L��~��Š���*��E���a<_\�<�G�u�<�}�h��<��=r����ǵ���<Uf8=jLx�Mk��Y<_/9���6�VN=e��<, =f����<�<6]�<eʼ���?қ�nL6=�xw=a)L�4��;Z���%==n��=��0�5OD=_ `=�5=X؝���<q�g=�Ӻc�*=����7=o拼�j�:��<0�W<�*��$=�]��j7�8�bS;��<�ǒ;�+�=��P=cq<��$�;oҁ<��L��I��V2��aA�� �<���ڧ�<�d=��]=Bj'=͈T=Ȉ;��L)�����6��=Q@������)���<8�a�B�-���=H��<Nߴ�`���:=�~��n�SFA�o�<]�=v��n[�����F>�V��O�#;J�D�f=�oi�"����$=��d��=�{�~發c��<�U=��=7=)`7<r�=�^��wq��+X=�E���v��:�8�>�=�dỰӮ<E'$�I�輼O��tF�:�ď�p��'�==���<-�<�C�:t�r;�_\�Xd=wB�<���7	~<��=���<%�����
=�Z7�L��<�.��h�R=W:�0:��
6���>�װüE�^�� �<�~<=ؒ<��A����.��t49�Bg<x?�<L1@=S���������ɨ�A�z<��=,������00=.�'<��<���4	$=��1=�Ǽ	=�r<�<=Bc=Cb���@������g�.E�;�G\��ݐ<�:?<iZ��.	������;���U�D�o�1�W:ל�<���兒<z����w��;p+�]�;͐=��'��%=��=���������<�������<<�=�b=��X(�<���<���2oc�?]=(�=0�g<�<��JƼ�7�<Rl��n��������D=M��.z=�Q�sMI;�ݘ�j�&=M9t=P��<�m <籵;5��c�='�%��<���F�wא<���<�TC��P��q����]�<]8=����y�U��� nM<,~�<5Z=Zb�r#�I��
$�;�⣼�»�c�g���"`�:e�<o����@=A�n;�k����8��ɀ=��=2]��PS��M����6<�oR���<�+g�݆�<��������l���2=�R��qs�<ü�<�@�<:��<Yf<q_I��J�H_C=p�T��}6���G=��*=�Z-<�z=�k��Jp0<�}q<���<�D��F�iE�<���<}=��(=ǠW=�� ;��<G��y�B���Z=%x�"���Zr$�=�<=�*x��@��w=V��:�$��f�p�����+�6<�=�7�<ݲ�=��;�d��Z<s<��0=@%%=�R(���"�ն�<��<�r<=1:=j�1=��5�<�}b�M	=�z��Al���*���<=e���p�%�+=�P,=��s^�<]c�<�;:��V��R30�T����*���:���C�%ѹ��)^�]`��F�^=n[1=�=�6<���<e>@=1���z�=�㥻-���=m�<
�=�~:=�|K=�,-�G�;qV���A<­��R=3�!<� ���2������=X�<��o<Ӛ��v=.�K��<%7 ��=A:@�Ƽ��(<�P����D=�~�ul��3��<��u<\H�<��������_��n��C�<�#=pS:���<�XX=��λ�O=c�B�w4=eo0=����"׼�üC`:<�:=o,7=���<,�=�ir<��<|ph�Ì":� �������<(��D�D�vt<�G=�-(�����,���,d��l���0=���<��#=�c��d���C�<}�
=]�S��.<�6=O���m�;�p��և�ԞD=õL<U�<[�޼!C��j���-8�0K<z��f�߹��.<�=��g�"3!��p<�*r��=;��8=�a)=�=���<T\~<�.�</��;���B�=��=�i�<�Q�<K~<�P�d��<�� =� =
E=�8��8o��"K���h=T$�슽+��V�P<T�<��%�?8^=5��������;b�]=Y|U=`��E<��_���&9�?B=�$ռ�a�;wo=�o��g���7���޼�KD�no�|���::L��"=v_�@u���N�<�'<s8��D�j9�O>0�>�j���Ǽ���2(R<z����&�b���\�M�P;q�@��?ּx��q.��{�� =�"=�n=j�<L��<n�<H��<]G�a�O=�������<Z�c==�#=��	�q����D9�9�p�7=%��"��<0�E=e�p�~���R���$�<�{��:�=���z0=��<ۖ=�+<�l =�K�<�u�<�K_=+r���E��􅽺@=�m�;��&��	�<5�\=��<�D���
�p ��B�F��:��Ҽh�$=?�1=�`1=巠��=�U=����)F��e�<.k=b�T�Y<� ��i"�l��:�I7�)�¼ٻ�<^^8�z�<���
���м���{u<�Aq?<S�M<Zu׼�=�� �9�����<^T�:�<kx&<]9c��Z�C(<D�t�$;��<sA�<�x�<w����9�:K�_<����֢<����4R;��_=��9��;�L7��o��=.=��&:U�=�Ȁ ������,[Z=Yr�<CQ=��=�i�=��;;x���<5���w��=)AD���K=)��<4�D=��p�
�M=5�=��.���Ï�;0�7��R5=�	�:�(=��Z=�J	=5~j�	</=Z�G��2�����9����L==��r�μ�w=��;ٶc�AS1=\��<-��:��=k^���X��e=��;���<)8���u<&l�S`�<:j=Ð�<�$�D�&=c���
��7���9
= %�<��<��	=�Q =z�=�Z=�v�<QC>����<�FH=Xa�=[h�УU=���IѠ�V�=�����;�\7�����z=E5|<��\<�mb��,=J9f=�R��d)$�"�p=#1̻�8��B��$�=��u="<����d���Cڛ�M�5<�6S=eO�:�ҺD������˻<��i�&����iμ;������;I)%�^}}�|�*���2�3�	�=S�}�'���<�.�<�G��<է���D�P��<�=Ll/<-R&< �6=/"=0Q��������^Eؼ �<�{=��=�T��]^���[��L=�==V�<eU=Y��;�����ջd�=aO; C���<����S4=�����o���B=]�~����fJu<?}J��� =�=Q�B;J�=��M�
�<lV�WJ�(��<��3=�n=z
���K=��S��B �M&o=l�<��5�6��%��<D::�@м�<�_]=��<�E�������.�\�Y��5&=��<�ԼUL��B�໮�q<������.�,�Ѽc���-��S"=
�O=o�d<m#�=��7=��_=�$��O�T���=Ї�<RJ��b_�J�`='炼��D=���r�AX=[�eȑ��>$=�6Q�<�Z�I�s�ٱl��g�<�J$=(�5=��$�2=�1����<"�<���<&%R��*�<�<�66����R�<<�t	=t.�������<|�reZ�8������_�)=�����{Z<+�".��?�_<��3�����}�<uS==����*�<��U��� =�Z�9�<��͍<�ǧ�!�U=�z=��=j��}N<�Ѡ=���<)�㥼�@�s�B��&(�&E�<���4;}���ɼ��	=�	�<˾�3=�?H=� ��΄�~\=|��<=4��,��׻=��<M�qc�8��v=�k���	�=����|�<�����0��:�F�8;%d �q�e=q�=�=�`��<��w� ���O�g�O�vH˼�Q���<��� �g=��E=k6�R �4A#<�=Z��<c�6=	%F=z)0��j�=�2s�������=z�����&.�m�A:TH�<�=�D;���h=�3c= 7��+��i��Z�˻�B��fE=��`;�y�YT*=zu �1��;�6;aԌ=vV��WX�O���i4=嘄�ɔ�;�(A=�w�����u�<��~���'=�)|=��G=�r�[���[=��;Z�7~l�=�E1=Z�@=��5=��<�|Y��r1�/^A=F��;̑����<�<��=+�.<D9ܼ!�/���;m��函�D�<�c=�=��(<�Oo�0$=|�0=�I3=��<n'�<܅�<�<B]i����͝𼸧3�I2h�(��<�=w<�G=�U��x+�<�k<=5~���6=L�J<zG����I�~D�<'���%�;~��<=N<<|���Y�g�=����9��(��!M�ƎK<�[=T�4��N�<�L-����Ȓ�~B�{P����߼T��R��<����1�-@H�!�<���e�;.;�����D<^1=ٕ༕<�<�y����<��ѻ�g�<D�=x�&������A=�=�!&=0�<)�f������=�_�:���ev��,�'�>�Q̼�t���W��u:=�<�=��`<�	b�}b
=����<!�T�<~y�<څ!=ꅊ���m��2�<8�<n�<��ۣ�YCX��ʼаO<&́=��c=��<? �<a��ֆ�;v�4��j�R�F�4�hҘ;O���df=x��<6i���&_<������<Q�S�Ͱ�l�=�[)��\�;�V���Ζ�������<%G���=�<�be��%=dє�=7}<�=��5=��7���Լ~z4={�Z�⃣<��i=X���"S=0.<@�<F~��Њ ��Ik�~�<� ��ĝ��-�i�.<�@��6=:/�<��U<6ʳ�k�}=Z��:���3��D�=�&6�+
�<�J=0<��)�K=gJ,=��c�WL�`>��I��� �����<&���}�<6� ��gp=�_0=uj,="��;�~<��< ���#=����m�#=���;���<D5�<;�#��_<Fk�������8�=��>�p=�v=��)��&=�c�;�ͼ<�';���M3;=�wֻ���X����F�<@�_=ȴ�<&=l�k�==���<ͱ=/Lq<�EG=�k�=�V�<.
�>�I=f Q=	F����;�"J=���J�?�v�(�=QC=�;X���4=I8L=�����:�kj8��Qx=/̔<���,p;)J�<#g=���Ýj=������97�ل<u�ɼW���� �+= 8.�\�=2�=�����<�(�?�b$=�'=]u���̻���Q$=���<�E=U/A<_׼��=$�]�j�I6z�6��_6=E��:=�<Έ�:$��<|�v���<�G="L2�j+��;����<�]���Լ�E< ��m�z����{�<�du��/G�\�j=/�ӆT��������L�>���̞ �/��<J�漅��=�Zl�ެ༄�o����<��P9���:oGмk�.=&a�t����	4;R�r��%��.�
A$=[��%=�
ԼF��;�p缉�c�	Ok<���B�Ż�&��=6����=܂�;�7�����)kS<
�2�Ͱ�k���^����<�:��3��x�W=n�Ļ�Z=8p>=~-<�6��:V��I�3~=LO)��p�Z~,<�Y�m]M�_܆<�Z4=�s=�^3=oh���|+=�<���;q@=z�<� �|���1�����l�Y�<=O��X���b�-�s=[�r=�'�<�.�ʒ���ڭ��T�9=_�E=n�<��H=���P��b�M=���<r[�<֜+���ݼf��`&�=��9���x0=O?�<�ݏ=iN=��z,=N���yN��`B�(�;��e�����  =��컽���L�<�א��4��K����&<��'=�{��}9������l�<&�<��<��>=�;&9��Gl�`y�;����*<Q���G!�v��<_=yoj=]���H,1<�=��!=2���-�	=�#3=t�U��@����;�m��<s���}?�<#c��C�㙻�:=�5���G#�\*=3�E=�W;��E=O�Ӽ�k����f��z��2��<;Y�5r�<=~
=dDA����=�6�<��=�OA�� �6%�<��=F��<�M���R��p�;�Sm�{\�d\Ż��Ἕ��<�=b��~Ls��Ӽ��S=��Ǽ]�Q��I��ڎ�����6]D���ʺD��<��a=�!<hֹ��;\=dȋ<��=�S�$MW=�C�� 8�|u=��H<���<�e���e:xꪼR#=�h�<Y�E���Ӽ��|;���.P[������<�<��}<̵=�!=��<�i&=�@5� �d��5�<p6=G�,"=��]�!z�<�=Ɩ���G�<� 8<�-�t[�:�@��;�)�^ֺ���<o�#<^����Np����<�%���x3�=]=�B�<'�6=��;�,I=~B1=7`�<��b���"�B��������+=�\��H���t@�� ;=�e\=��<#���G<�����D��
r=���a=�w�	ET��eD<WI���=n�<��.�1��2�n<�]˼��:���<j}�
�/;ol2=?��%vY<�֑;-&�<�����O<*Xg=X%�V��<�q�<��=y�����\�o��.N�60λ��>��؀�x+缂��=ߔy=��M=J��@��[IH=�1<�<F�J��:Q=��Nw<ݯ)<�.=3��<za2=��������']J=�-=\�;=0+�M	3<~$�<�"l��q�?<F�9��r�<����[
��l�1�(�'_׻H�S�d&����<	n�V��w�;z�V<�|$<���㻅")=t�=�a=L���#�¼�^��r�	xS�o�L�R�<�t��g���8=)+�<飨����<��`�S��ȸ,=r@j�P����'=T3�0<�3����<U��k�9=�y���e=(�l���F<��E=�Q>=oF�a���<q8��?�fo�<+�?�$=��!j��-O=���;�m&�9�=s�=���׷<�z	�!�;i���Nl�9���<b��<�?�<֊ؼ��=���;@+�<W !=�/I�����ጼ35�;1��(��;�}7=40=sr=�_U<�r��V:��9�=�Z��s�\���~<&�"������m<��<=�ĭ<T)=�a:=��B�,��<�I"<<�k<�P�;���<�%=�O�<R��<���G���Gq
=�&�<@8¼{!=�M�<@�C����]$���_<���^<�B��E�z�����ܻ^B4=r�<���F��G����R3=��˼�o�ݼ߿�;zO~=���b�5=�}3;�=�+*=v�<���<:R=�)<�[��%^�<��L���`��~�<����U���!=c�=��;�Q=��ڼU͛;�8T���-=��\=I��<���<F��<�?��OT��3��� =�[�s >=�w�:�A��<>C,=qU���Y=)����Ƽ"��<�ϼ	�=��c����= ����(<�q=^\0=&�.=�D���Ҽ���V�j���_�׼���<���;C�~<�TH<-Nm���=Q�������<�wV��7^�5I�<<Pt�JD=�@����*����;ǻ�y���ID�Q!3�'r�-��<A�˼B� =w3�����;P�� =��P�P=�<[+��E�=�#=�7��K;�<&#^��N<��u=����eQ=�y�ݛ<?՝<�;5���<�j9=�I�<�m��z6<d��;#�m:M�1��<��t�|?B�e�=o|�=�e�<�W:�`v�ϼ�Y��<H����'=FY)�Gl�D�m�;�q=��\=�R�^�A��{�^!=�(@��u��*�<h��r�=OP�gEc<_����o��E���<��S=~B0=�|=��=gN�b�n<:��;�3�;�d=�	=,^�<բ;�>�E�=K䳼VC��g<E�:a��J�$=��U�C_�:Z}�; �I�`Kv<s��;�Q���$=�=�;���F�"|�<FW�j�=8tG��S=0,�v;� v��)^=ݤO��~ڼ�9�a<%=���<�z_<���;�"����<�>�;s�4=b�y=�F�ʂ�;{B�K>)=�Z0��CL���;��5���;�`�;�����|���q=���<D4ϼsmT='n0=���c����? A=�<e�9�u��7���<2�Ҽ��G�J���[��W��+=�z<g��Ӗ��z�<��5�����:�9���=s�:=(����y!�t�<�s4=e�j���O�@��<�W�;�B`<Z� =#�e=̕D���z��5=3IӼ
�*=s�J<�Ga=�2y���=�w
���l��/=[�k<��a=����.�;۫����o��I�Ě�<!�W�8=�o;�ϕ<�V���"=�,2=�^�A|���><]�2�{Sɼ�h�-���3<k��d	=�K��
�<4��(�*=��$=Nt���.=��мGʶ<�w�:��x<�x���� �f�3<°'�619=��;��Y��R��ř8��q�o�ػl�-=��ϼ�+3;�f=iL�<iY4�B�S<�c��W�<:�;'M<�b���&�_�-<�P7��2�Ǔh�Ƶ���y;�\$=�����J��ָxz@=lF=��X=�N���AԻ�b�<�����}�<�,����<��u�m����<Ye=�������=��.�#,<|zڼ�'�;K��;�ߐ�+����<�G]ռe�h���d=��D=�ۊ;3�<
)_=�:=��w.=7=*EQ�� �T]�=��	�x=� ����6=�gt����;L�������<�t�1�]<�O���B=�I`���,����P<�(�<�=�X�;�I�:(u!���g�%����<B�@��Ǽ�g��=��F9켈�&��AI=���A�1��y�5V=p伥|7�4޳��[޼lc�<>:x���<��o=��x=�2H=��s�A�z����ȇf��/
�<-]�<Ns�<���{���ƼxS=��T&=H�9���+<� =&y;j[=.;�f~��x��h�=��9=T�,=�O=l�<#��v�Ǽ�7'=N��8=q�߼�.=f�a=���w��InP�Z�[��<������ڧ�<�:1[��1�<)|��W%=B+��Yļ��<p�Ѽ�~��;���'f�<<�<7�<��m�<�=��==�v�I�U�Ù;��=\z���[7� �9y��</#"�?�U=�f<F��<t�:۷q�b)�|��:coz<��=�vs=f����?���E��-=�51��2=aQ���<-�<��= 9=C��<8��;��m< � <L�]�y:�K= Z=L[!<@�P<�$��v����\��<�"�;n=5�>=�u�a�]=kJ�<�$�����l�1��p<��ڼх=9դ;���<���<��$=�K�<����h��K1=a?=�-����&�a�X�W�P���=�>=8I7=�L=�p��z��o�T=�[��2�i��;el��ռB<@<N�^=�9[�����BV7=b�K<�0r���=�v�������<:�<7�ֻz�;���g~�<�s�<��R��sb�0���������&<+�")=�^�����<t=�*=~�C�8T��M=�t��`a=�#4=�^=I����x�<zu@���L;Y�|��=2=3�Z=�Լ�#�Sj"�e�����ȼa��;R�-=�K���f=��;9,�<�8ڼ5�<<�8�E=�b�;��t��hf�+� =p�T�ONk<-�<C�p=��`�a�l�IJ=����j=��b�C�;�*�:/�ż��=ROO�&�|<c�<5MG�G퇼1�*���<��=<`�%���}��P=!�;�,?=놼 _<��[�ݻ�����׍��ĺ�)n~<�8;��¼Z��;^�<6�=h�<�e��=�&�4��<���u=az$=,)<�:,<Q�;=�2'��C�г2�j3=!�V�=0�<�8���!�<��<���<Ҧ:�L+=�	m=��%=��d�ɏ��ޑ<SV�ʤ����<.C/����N)�<�"���=�@I<�����,��ݛ=����N�<�!)=�1I=�=M왼�oR=�#=Ir!=@'=[m��<y�<���0���=;��<�=��?e=^61����<_�^;�rf<�k<�����<*R�<�3ܼp���O�{���／b��5��<�?��Հ<��7=6�����P��V�;E�:��*���X�qΤ���2=�+n�C7U�Ɔ<EҼw�ϼbfj<:D@=�� ��<wE/='!����"�=S�w<�;�<]fļ�>=�L=�Q�L<�O�<c�0�J�ݻ΄�=:=��=�-��������G=��K=V1�С6<P_D�:y�<��^��&@�Evu=����x6�����=��<*�D�7hQ=Q���K̼�J���7=I;==c���_D�Mb�CCz;�ư�AX(��j�8�(�<���<��p=�kA�E4�nN��M���j)�<+�<��i���<ܳ�<���i<M�<|�M� ;�L��ǫ;і��P��&V=�^���]����B����<|�b�dK׼� &=��i<��?��=}%<X�C<��(=2g"=�_ռ�z��H7�t�<��]��;5={�P<p��v��4�g�E����8=�u$����<y��<�eF��d�1 =:�:�7�<�f{=D�[��6�<��<�p@<�5=#��ׂ ��R���9=�L�=��R� ��R�JZ=�qJ�3 �����Ϸ$<�u��*b�:<H~<��8�v��=..=����k<�|A=�9�O�û�u=n�4��.l=F�\=;hR=�ό=l��;�CY=�g=�.=������&����������<��]=_�9��4�<��	=d�=��;�o���H��!�<l�¼.�%<Ռ<6�)�kW���0<���<���(���A=%��F�<�Œ�k�s�|�v��a�<e�	��:�U=T�%�=d��U#�wJ�<�UH;
�.��=a-@�c�����=2�����<�cH��e�<2h��.=�r\=9�<�����6���<I=�c�<�v��,<�e�,=;�f�',7<:9;i��;`�P�P�-��|!�X �<��<m�<�h���e�;,��<U�<#�}�/}4��;�f�<��M=���;�(ؼ����Ӟ�; Z���j=��<�8�H�,�@�N���~�oQY<�%U�<��=C�5=ǩ�:�B��<�韻�7�6�<5z�9�Z�B�Rk���;=��= $b=�>�����d�,=��#=��w����V�=��=y�t;�����Y�I�5=�i�<
=��*=���=طڻ@��;H�<��C={����=���<�(��JE���?�<�D6<`=HR5��tٹf4��a<z)j���GML=�B��H��h��e�==��<9=K
"=�?<."=Խ`<ф-=t�H=dj��5���/=@�����~1=��6=m䋼�UG�`�E��}V=�8=1�a��G=��=��tc��4л����x�<�3;�<��)=�А=�pO=k�h<2�=�'<��=Z�<遆��c=Fn�<7����{m7=YO���1�� ���;��3�<g[��Ɵ<K�S��߿�:y,������2����T�;0���?W��Yg�	�<\2=YX7��;�f�=,?Y�2������{<&�W�0�>���L=�|_=|�<R�=�(�<}	���5��>=^���ۍ<F��<cb�>H=�e�<��<�D�=^�@�-y��^�����>�>�����t��G
;�b������Y�)k���=]=��<�n�<'�"<k��:����$�.�%�ռu�;�<�^��<���:�Y<z�<U�6=.��< ֻڽ=_@`�?�R�*�*���ټ��2���=$�����<M������	Oֹ L='r#<��-��-<��B=L]=�k=Z�X���ɡ*��X�;|�;��ʼ�=�Q�X+�<:%,�n�Y�D�� _5�'<�>����߼�*=�)��n:��C���F�Ew =
I=y��<�0'=��'�w26<��b=E�l<�$%����<����wF�˴C=$]e<w��I8#�C�T<�޼G��έ�<;輯g)=�c=���<����'�;�͑+:Ļ�������-����;��3�����:<�=��\��v=![�;�5�<�r.=~6=�%h�|�S����<���;.�;�=�;=�V-=�'�R���QI="�9�CvG<��\�>�<�;�����=3FI=6K.=(��Zj;��:="/<?&��<8<���<3\F=��=K�,=K�T=1󴼕�=E�I=��N�a^<�+?=>�=����u=���;� �.;��ֶ<^��<�4�=�8h�Qg��K�h<.#��z'=��=z
=;�<b#���P=��[�!�[�~�=4O���n;M�=i5���s=�Ch="V�s�<|qb�+(��5��nY#=�=��;n�B=�G=&_<�
]H=�	]<�\$�C4�<G���鍼�c�;b�;�蠼Zc��d9����H=��<�^����!�` =�J��u��<fa%=	=�r�tJ��8��1=��=+=��:=�'���j����<?�e�o�;]HI<�ż$�&������x�ˍ3=8���[d�/�K<��E=W��!�9���h<o*�1�<A���|λ|�ѻ�(��@�x�Wa&�ļG4�1$s����<K$V�KN��͢)�I�L=ɛC=��f<�T�5C���ͼ��H<°���f�2��;Z��=RX=-n!�=tIA=���v�7<pK6���*�,���5ռ��l=F뵼��==��,=3�<3cd<�x>�{=���<�-�<NP���q�^��<�9==���i����ev=�����<�� =�� �h=�L�<��X=9�;�n���n&=0����,�/��<��e�8�	�Uv3�*y(�*�%�� =�i�0g�<��<ddi=�l�9b8��%�J��<>.��E=�$=j�n��L�y���Ӂ:[������em�R�<W�;��ۆ���<��\�.`��B@p:1�=�<܄<	s<�B���ї�:�F���C�r<\_.���<�Y���&= �P���.=���z��k�;�������:�X=K�[�Y�3=U3<�|�<:{(=A����5�g=/���F�Н<���姼(�)<�G=��<�����2��>�B=���<�]�=¬<a��=',V<c�p<�N��-mb������;=�c=�f��.X<�i� �^��aݹ���� ��I�9U���h+=bE����*�QG>��a��ຄ�¼�� =��;�I�����H==SX<w��)I����=�|0<|�%=��<Ƣ�;+eW;k@���4׼��<����劼|�O���<�s��i0=��ؼ�.=�ԩ;�`�-F:�-q�<!�==���<��T=�i��bm�P�/=N�;�&Ӽ;��_�<=Z�R�=fv<�G=��j��o�T�J="�w�S�Ź<�*�ז^�@��<�����O=:�L+{�=q�#<�쑼��ӻ���9�0<=:5=Xܲ��m�#��:�킼�]j;=B=g�P=|�� �;P�M��1�=�~��N<��;��!=��=Õ�<��s���'=�i=8䁽���<�ؗ=i!����<�m�<���<^�����͏'��4=08=��%����@��(� =#�����<�J=)��`V������^��N���Q��H
B�]K�<��м�&�q�ԼB=��u�?=+:��ή<���j�<F�n�]���(���H��j�<�s���^�w��=�2����M�?��Z�<	�<�7V��`��wǼqs���O���n:�df
;m�����<bb�<C�8�< �=��R�YXE=M\�$���7��4�l�L�8U���p��eC=~*��%UL��߼�&�;m��G��;K=f	J��Gϻ*�/���d�k� �ˌ���ir;xy�=��=��<���S*=�k�����<]�=���2<cIR�i��,\�
`;r~n;q �</P=������{�E=���<��<YJM=L�*=v�(�>F�� y<?X5=�Vi=8Y��9$=��1�&+`=�)���x=��<�ZF�*��;[�� fY�ꋼ:]=����N��aQ5;cz<�6ӻ�h����<��¼䇼��:=��<�j<0w�=V=�ͼ
�B��&=��:=E�_�Ye�݈ =d�s;g�!��{=�m=�ę�<�j�~�ļѭ�rh���(<K�G=�K�<yd�'�t=Da���9�<�V@�Q��y�c<@ͼ�=G�=@��#��=\��{�E�V�	<ִq�f��<��<��'=QT��u���m������W-����<ޙY�q)��	�'�R�zP�<4Q=J@�V�軁c��-��q>=A�0=�~�;#�2���Q=�q0<p0�<|;F=��A���;��:=R�<tʅ=B6�<�>�<�'��I=�����h�X��<E�R�߻d2;>.`�e��<����ky��5.���7�����1�l=sJ�<>��;����_~�?)ܼ�"�����<3k�<�g$��B=oC�<�>��z�<.�$��ؘ=I�л�B��&�ѺE�O<=&=ĉu<O�
���=����GD;Z:ۻg#�<�54���;|�L�8_��"���<?m;�M�rZB=�~���{"�g��~����z�9�,�<dA]����<p�="$l���=���<N=^i���_=�!ͻ"W�<X��<-� �J���{s�<8[$����	��������c=F
:=X�=�$=��	=M����<��D=�1s= yy=����=�J=Ai�������.=�;29��u�SC;�v"=�U=ʼ�t	��=��LP���;=/�v�
�}������y=ݶ���2$��,Z�"E׼�"��/�?_�<�J�����{'=~o���A�2��:ʏI�/�O=%�$����13<��_���;�P�<_.9�fVk=�6��hg���<�5=����`�=,ZJ�9��<�w�;�b��=g���q�B=T�U=�>=Ed%��=������:6CY��&)�������<�-J=�<P��aG�A�v<����z!_=m:H=�;�:�]z=��L��#�'Vz=C��/��<_%�O&�0�꼔|�<��<��-=���:�=[��<!���a��.�
mB��A����n�Е =�(<�Vv�.�Ҽ6�_�[ia=�1}��C%�Խ��ȼ���=uu�=�kQ��s<��Z�� ��:���X���R�i�z<bU����_�i�A;`#h��O=��/���S=}�H=F8�<$�u<#'=�Qj�L��ťg��7�S��:��z�	vg=S�*=��c<�^������M=�@D�?ɉ<{ƿ<�>=�/�<~	9���T��H��c�<N��<e���m.~��9T�YS�<]�@;���;
%�<ȿU<����nN=��H���;�?�;1�����=�
=��<;��dhG=�|D=;8��Ǜ�<�<��	=���� Ǽj�_<���;j@=s
n���;��=��a=M�@�C�_=��c�.b
=���<��7�KL��.���4�a=|�D<��~=�R<!������Y A��"
=�Z����'e&=$�������c<Pc��~���*=�!�<�G���6=ԳF<F�B=�;\�<=0!1���T��8v��8O<r&�Չ=ŘѼ��X�i���c=��I��;
�<.�@=
�.�:�X���&=�v>=t�<�8��d�=������6=d���P/��"=LW�<�6�9��׻"��;�ڼ�G_�}Cy<��
�b"=[O=
{=�Z�%!�;\-���P =q�Z�"����
��r���v�n׼�����먼}4�<�X<�I=g��8���I�<��$=�=��l�
X�<hJ=�ck<Sl=Q =�I=-u�Jd�����<= <r�|=�1=�H6��y\��w�Ub ���7=���<���=�1�;��<�FK��g�<��;��Q=���4D�=��-�fW�<�$��S�M|=Q�}�܉=N��<8{c=�z��P�<3��q�M���6�YFt<Ӣ��4nҼ�Z ��0<�ѼI=��4�#
�<ϛ8=�k������UI=�U�<�==��=��{���F�8���<�w�������:=Qã<���=:���K8�<jw;w>�<���=�v�<6˝��G��#'=��k=Sm=�Q�<�.7�Q����:�k;ꣽ?ME=m*�;| �;��<�V�=�%p=U~=��M��]���~���w=���푯���<�࿻̫2=���;F :=e	�p�-�F���8�6=޶I<��=��L:�1<����<��=�R<��
D�<����)��?�=*�]��Z���N=��������/��<O�/=�ܗ��}=-�\��c`=��F=��	�@]�<#�g<?֗�E��<�����;�p����A�_�w=�807<Gl<=�0<q�6�~�s=��<w��<���]��,�e�j��n.=D�<.K=�5ۼh6E��^��=�l=�#���%=&��<����Yܼ��u<�t�<�;���9;66��d�m���<�G�<s������+�<�:V�`�;q�`����(_㼷�<-Y-<�v�<�2�<�L=�Ɔ=�ľ�
�W=����2�;LG���<�5=�=�<�I�E$<�-ϼ,�S$������<���<~@:�H�P;3�;=�&#=������=����!�G��<^
����F<"�d=;�<��b�J����=u޻���G��<+�T�aZi���x<��d<�X�<�H��������D�UJ���`=���<�C=Y���ߣ�O)p=��׼V�q=/�=�f=�\y=N�üC����,�<�r��}�=��,=܂ػ�=��R��%5�]<��`=�H)= ���X=빴��X
=p�a<Mn�<<�P���@=i����!:=	L���>=�-@;�=R<D�S����9��S�F�>=����H쁼v��<!�[�k�<H��< i7=������<��m=���<�l�;�=d�J��H!=�4=yH��Vn=/��;CL��6K<,B�<�=�+��bSN�tuQ���A�|`<�Or���һ͔L<�F ��M=&�9��&:�)�<�a�:��'��e�"qZ���-�� �<pw<�u4��US�:gP�FI��� �=�;���^M<{"�<uJE�U�<�FF<�<A88=�WO=0;/<�,=��ͼ� ��s�C�=� �'�"����<�X�����;%V!�r���g�G��yX;�T�<M��ʉ�f�һYE�<\��<�}S��Q���/<�Zf;z�ȼ��L���;r�R=��'=�i[���#T�|"=��l𼄀�;�����.;SQ�c�o��ϼ��L�$<�w�<�P2��㪽����W=���<W =K��OD�<�a:�,#=3���mF�S�=�p���1�Dj=�P�EeJ�
i�A�=k
==T<B=:�c���<:'�<\(�;h��T����<2���;>[=`��8�|�Q��;;�[=�ք<�른�K� �< �$�o��;��<���<��f��μ��F�|e��4�8��~T�;���<E�=K�ؼ���������<��=��@;��=�5d=Q=~o漣<o�g֋��8$=��8=��<"�e�3Z�`<1ӻ�!V��J�;�l��:�Ś;�������B=�7�;Y��<u7E��d�=
{>=x^=�7$=�w�<�{=[�|<]�¼b��<���<v�&��U%=[��;69=�OBL�nH�<�|+���p�
�=��P��&�<�X�<���<�ׁ�!$Z��{��}�k�钐����<Y�=��*=t�U=�*b;�P���i8=}G<�N_�O�?�a�	<�`E��<8���]}L<W	�<�e	=��!<���;?��t<�G��(�<���<���=�<�<�y�l�����]�<���<?l=Ys|�~R<5V��F�N�<>�+=T͇�� =�P��-2�j/�������h�?�Z=�<�RڼXu=�j������.=B����;3<��(-t<��G<���;���< P�:-AE=�e=B�$���K�[��<dE?=7᯹�M=p��<Y�=J�[��f5=�=7W������֗;��&��T��V��w��z�μ�C�Weܻ��L���=�tj<�p�<y0'�5�,�^Z�<a^==8^�����^
���'=���DgD��j=��-=/���+��S=�A�D8"=��0��Aռ+k{<��8�:�#��<y?�;J/��a��+$�m�~=�J�<��<���<8��$�/?�ؿ���'��@Y?<���<�W�<-���?�<[ϻ��q=��(=3Z�����<ƣZ��/�Z	��IP<@�<���1�<ӈ"=];��u�F�O=5�==�u=��(=�����G=�H=�~,���L=�N��ge��z,�r��;�4�Nq3=D=n!=J�T�^�Hx�G}K=(�}=�)}=#�V����<x0=z��<T����=�"�ӏ޼�ۻ��� <~q�!hh����H�w�H�8���H��qϼ�x =��;�!���.�Z�+=M臼�u=��P=�=e�<�j=�s���T�=���=eͩ<Վ=�J�;�I"�p�I<tx<��/=W&����J=�=�H;�6^�§m=�� =PE�<�kI=so�<7�j�W-u��!$�;i����A=a�=��	=�su��C�; G}�4Ř</���=�s`�L4=�����#=Jx�g�=��<�]i=G��`
=~¡�B�<�I��؁=;T<6=�@}<M�=�J��.��=�����N9�>�P=������;��<�5����<�鎻24=��8=0��;�2C=Ҷڼsd�=�?n<��<��<��F=��@=쥻;5��;�S=�80<7DJ���#��@�;�N���;|�+�ĝr�̬켵/o��I=��V<�Md<q��K�;F�=�Z�[U���!=b�<�u��c�\2�<,�1�1sy=K�ܼ.#�<��<5�C<f_��Xr�<��*<]~<ۏ�OkG=:L��XG��_��j�<�|J��`�z�R=��v;�	�/:R�y��<�^!=i�.�GFF=� W���<���<P<���K3=>�P����������Ū<uW����W<E.�5�D=YF�<a�=^���ļ�5ż��Z<�?b<��<�<>�`��2=��D��4�;Z#��Fr��5��N����;^X*<�K�:�\��=��AR�)+F�j"���E=]���2-=..�<1��t=O��<A�=�f<��<�{;�g�tf�pT:��v=�=,���4��?�����=D�ɻ6c=�0�:<m���@����<�Լ�]�;p��U�<�|M;5�=/9��G=R�]�o��<&Ѽr�P=wj��j⋼:�:Z|�(+�K��;�z�JQ�;��<<X�K<��z�1H��}��A=~tx=�wR�/��dӼ@Q���ǡ<:d=0iʼ˅�<�,8�"=��i����E9�����Z2>=]�%=윚��m���G���<��=�p��v�=��J�
m	��p�Z�=>��^�=U^�>ST<-�u<�z)=�-"=58�<�J����-��i�<=ۉ=��=��<l�8=
9��=WU<�3g<699�\w<=����t�<LL���=�8-="�E�;����3=1��;��*=�fD=pл��<J={�$�n����s����<j���D�=�`";��-=�h�<:� =+R�<��6���<�˕����<JN�;z��<�(=���<��<�o�<�H?���5=�u�<�*8=J��U����y����g��<�h��؟����V4R=�����=*����=Z�=�N<�D^�*���6ϼ�$�ƽ!�$��<�x}�39`=�sn=��<��-�Fm��џ�;s :��w=\�:��g<����Yh=�=KA�U��<��B=PM=��=f_K��c����<=�����X���L:%s�=M	��i�<}HH��cu=��(=BE߼k�.�`b<��Z=�|�<m�h��<_=�`4����<���<�<6R���,=ؿ��,k�&dZ��A[�F+�i�^�b�ڼ:�=n�	=�9<���=EN����<񒆽�g�;���<�gA=C=�^<�O����<.V;=b�N���~�s�I��]�����5�=�|�<���4�]�4'N���=O��4@�"��;	7;������!�<��<��q=K��;����*���k1���=0D;�u=�l6����M=�)�<bR˺k����,9<��T=��=��=��N<�s��~�<����u?=�6׼Rk{=�\�<t���FY%;[�=B�+<��@=�S���=R�6��	��D_һA��<�4��|sA��I�<b��<��=���<��;�$A��Լ<�gy��c�<��<C᫼�U���<Yf��l�<�W�<�Q�=�r�;�v�<�o<L�;9M�<-�R<�4����<�;�m/�vj3��V�4��<�~U��<��<�.�<D6=�}P<;��,(<ɔq=E�ۻ0L�<@o�<C/a=�M���9�J=�Q=�
�;�vv��]�<pAѼ�؍=z㉻g�=a�0�lx��s<觠<��~��/���nF<�J=Pw(�:�<����9s1=z��<�^=Sxr=�v(=h^���L=AX�<��=ߤ=�����%�ď
=�wu���c���5=�'�<��e��P=B��<�[����=��g�]�<ݝ)�#��<_Wۼ�s�V�=�� ��9p=Mq<~e=�Իڏ�%(X����<ikU�*T� (�"���W�+��v< �F�&��e�<NE]=��:�L����!��G@���V=K3����<��D���7< ?=��<���=�0���]=�/-=�̼�<=��=��c}�h�<X�<�CݼS1缠�O�r��+=��B=�z$���<%��d��z�<�I�<�|��Xk=�=y"/����<;��0*6��< �$�f5�<�E�� �ڼ�U���U=4nT;\e�o�$�;�k=t�9=��u=Y7���z�<?������U=��&= ���"���a��v=��L�<�
	�2�<���<�e�<��';r�5<Pl=G��<.o=�X��㟵��x^�nؼ17R:\!��ދE�3�=!��?�=+E@<<�n�� ��6�w<�3=7
�kX�e�/=>d=x�[=
�m=!���e
V�a�=��P���� =M��Q��6��"^=�׻'iϼ�*=2A.�3==�5D���g=�:=�LI��fW=���9�b_;���<i�;o�< =��;Uo�<�&0���5<+==���5�E��i���P-=;����!��1�+���Dg��<�F=J	v��jG����z�9=��b�։�$k���I�h�
<�����_�;FYT;��<K��:5�Q���=���J=C��XQ�<��<�M\�Ib��.==Ys<e6:=��<k�y��Ͱ<�ͧ���6=�K3�,p=���}:��n���Y|9���̼����9;qm�K���߽��P��O5=�9S=X=�<� W=��=�7}���������t�'0x���a=*�Y6�;�a��B��僛=tV�����|#=���;�z
=1i���*��7��p��<�wV=-� =ף|��7Y��V��<�<}k��/ =\Fh�7���ݩ;84W��������<ytk<WG�	�7����۽<��=�_L=ynI=Yg=Q=�<���<�	=M�\��ʼ~T=�腻�w�;�=&ٺ�g�<ׁ=�^=�;=�em��kɼ��f=72�Lj��J�W=ي�<vmj;��<�%e��n0�����4�=�9�;ʢ<�{<4f�<n*�kK=�_�<���:�}�<��;�v;�.�:;�N=�ܗ<o�;�
y��m=���=�\�<!
	=RHf;�"�;Ƶ���]=�=�:=G5<����� �<Nz�?���mR<����E����m��;�$�<��n=l�*�4W<�@<����<�8r�A(O<>�c�^2=ɑw�7�Z�J"ͼ+|S�k�;�T��$c=Y]�<O~D<G=�k��Pm=T��>`�;j�<��l;a����p�;��[=U�ռR��<�!C��S=e�<�@=�_���*=D~d=�h����<��C�=�м�5b�8yT�.�<w�����<D~e��H^��
�<��=}9�����J����M=�(���8oD����~A��z��<�(Q�@"��()�&�6=�%�<S:Z���?���,�u�E=F2�<���;�wɻ��<��]�]3�<lTJ��^ ={�8�l ټV+�qx�0E��(k<K���V=�+2���;h��<��<R�����<M=C;&�R���5��)�cG�<��м�])=\$�:���;܃ټ�H]=)(�P"K=���<�=��<�<���Ѽ dK<C��==��A��d��ٰn<�n)��="hZ�j����<(��;������<)f���(���h=�jV���+���R=DS컉��<�.���+=J-��0ػ�J��:�=v�R�F�;U�C<8����Q�R(B�)��<�ռfc=���<�6=����E��_?�o"=�ʠ��Ce���9=��=�t�;��<�ﺼ_vl�:�~��
=�咻Bc<��A̼��#=�,.=��c��L<�ď�U���m�(=�g�;�6=~���t�A��ڠ;�Ǚ<<���;"s&�����I�T����*=��?=Ib��e:���<�u��'�+R�;="H=�}�<��@׶���:�i�t=��<:>��%��ɼ�E2���Z=XG&�zv<*b���U=����/�<6	=�^{;��*=�����9���
p�,.ջ9�0��S$�Gq�<(�=�G=�I*��x�<��=o(4�~��Aϼ�F<���۰>=�2��F=Л0=/SA=��=ù>����;��=�����3=r���g�=����C'h����<��*=��|��~P<��Ǻ^�<?)]��;(���*<�P1���S=%U�I�i���`<,拼Lw�;��=Y-�)
�<DQ��;�V=�n�x;	=bL�<�3=�=�FY�;���Y5���>��X���4��g�<-=��������*�����=6����=�Wj�<,5=�Y}��}�<���W�<o<���R��o�`��<��,μEF��+G=��C=�
!<6����Y������d)=����Wc=�g�<�O=�@�<�%.<`56�fx=qV�"�=\�6=�;B=��;W�B�⺻�����S�<��Z�z���c�<|��<Λg���˼�_��T=��=W"��ut<O�?=�x���lE=c[�o��9�=��==Y��<�;xj=�%ܼ*	¼݆��O`<����;����[���Ȥ<��;E�==^�"<�b1=nv=���<c��<s������=��f�"&&���@���2a�<�$�Wp�=�Qλ�:�<��m~�<��`=mԝ��Oû��n<lA�1�<�<=����+�<�����3=f�E�|�H�9���/=	x=I�<"7?��9~�V�����A=�������<�|:�����H=|�D;�8�;�Y��q�:ꈑ�|[E=�&�<ۨ�:,u�<Mu���<)?a=w�1i<= Pf�c�;��0�E�׻��v�j��<]]<����G�<��<n��<k	=��x�V�N��wT=�怽�����=�L!D���<hɼ̀=c"�U:�~-�<�MR;��=`=����c���f ���=.�%4M���l��/��ܢ�v�6=�
R</�=�/=,*�����<j��躎����pN3���<=Xg'<���;GOF�lU���ؼ�R�P�=�G��Fr�(!Ѽdab<T�/�r���&�o�μ}{
�	G�-�H=p0;I_�={!�<�G�.7�UA<���<��'��^�<���<4�P?�<g�c�2=f��<Q��a%���'<m�t=�5<4I=|5�&㦻6@=��:�B`:�Sb=�G=��5��v���<�%�;k A=�,;�=-��1����	v<�|=x� =�瑼.���.�<�HO=?L�À�=�0A=�J	�B��<=��<���<_���<}=��<Q��<i�<��}�̴���9��!2�'�T%��N<37�<	D������	�:�D��ϻ;�Q���#=��G��a;=���;��j<� �<�J;�O=>Ҽ�h�=�\
��[~=�w�;،/��}�ͫ;>�R��"��@=����+X��0R;��Z����O�D���
=S�f=:�*=x/@<k�=/J}�U��<�\<��W�x6�m;=�=�.T���&=x�ۼ�P�<��4=u+�B�=%�T=# ��PA�s{<� ܼ��F=��7=ԋ���"<�UJ�E��<�2��7$�<e��;U�$��^����Y<���<�K<T�����F= M�8�0��s>�7�G=7G�<u�=?Z��%j=���3�����`򁽰rV���6���{�}/T=��b��G=�`�kma��� �~����n�TP�<I)P;E�;,*�a�9�*��:o�ʻ�|��TA�������:R;�#�<�8���r1:�#��J�=�v:�[7�œ5��i�˦Ƽʊ�<��伥����� <I�R�Zm)�Q����\������޼�]�3Y�<۵���㲻��=�G���q!=��;�r�<�l�<��<�'T�$y�<�\�<�Z����;�y�/[<�6Z;
 3=L��<zǉ���/=�++=�&�P�k�7��<LR���<�kh�;*A��9�Ve�XW�V�=)¸;k�;���=���<,�����v���q8��g�m�&<�̻.���y�<��J���=�.����7��%f=#e��y�+���Q���+;��)�i\Ǽ����5=�;�;��<��g�<������<J�A���d=W�t=B�*=�9<-���1g=A��<� �:j�G�k,�<�g#�$�}�r/0��/����'��j8=^'�<jN�<7<P;<s+�2j����-= ]�<%��)���_M;n�*='�;!3O=�����a<��j<�ϻN�<:B���:=u�0�M�|=�C)=YI�<�)4���<��C����e��=q�`<�|�<&� ��kT=2
���=W�!��� ~3����;�+%��8�<�Xz�a�.=�{�<��+=b7����Z�����:d��ls=g�=�rȼ �	��AS=[�漱�c�o���Y�h�'2�����ͻQ� �e�L���R�T]�:l-=�����L����<=�U<�v=�c�3E���"<�=q��bL������]�9�l��8��6�H�U�<�@��5����(���H���<�.=:�B���=W<� b���>=�C��p���<v�E��O�<����� =�R=�6`�%�5� �,=I���z�dIX=��o��F�<)J�����z���;8WƁ� ����W<7˽;��,=�=����+Ά<"?8= �λ�Y�;��R���;`(���X��+<&�J����<{�]=�ǟ��)&=��=�I<�C�Ϝּ=�D=� ���~�<�x�Pj<���<�!��$м>)K=��d��6�<��K�)=�u�<#<q�-Gx�N�üL��<���<In��U�<��=>�=�cCm���a�n�;a��<�r$���=Ԉ��H"�SO=��!�P�,:$��3�޼\'���!n=u2=k߼� ����"V�Ҡ2�p�X��z�����5P�!���0�&�N��-=�<I�;���N3�9#�;]�&=�1e���g<F M�;e�������[=�9<絰����<��W=R�Ѽ�Z;�8�����q�7�<!r��f(�ϊռy��<����vw
=��	=k�;S=)FY�J�a�7�<�́=�1��<��5<��zQ^��K�HJ=�E�!�J��m��'[�@���6<hS��U=ݚv=���<�)�}ڑ���ȼ�(H<����J�<5WM=%�ż��l=��=���<��żpmA= G���S=��A=1�<ʨ�<7�<4Р���<+
G��,�&��<��v=��.=�2��Gq�<%�Y=�"<!2#���:=MWs=�br=?�]�~�<��`����;��E�������<w�Ƽ^���gc)<'�Y�q�J��U#����8y��W=ӝ
=9�</t �;�<���<Z(�<�9�;�z��Ѿ��ON��=�������(,�<�6C=�Er=$e\<R/5���s�=W�i�9T=_�L���=KmX��Ǉ���=��';�d=�;�o_=-�*=�!<�,���$����=~`�;PR�<>��ق��9=��,=-�]P=}a=B�ou;�[P1<��e�9�<��_=�Y�;�e<��9���\<�� �9l��j���s���f=�=4�<;󍻑�=��<�"�>�<+)���B<�;.��1]��n�$�,=��ļ'0�����<��<��4=��!�N}=�=��C���<��<�l<Ų�;t� =OZt��T�X�C��#�<�1=�z�����X=!��:���}�
=c�L<3;n=�B�:\�j⸬y�<���<��q=�l�# �C�<�lB��y�9����j�1��<Uo.=��{:N= Q=^���;[{= M�k5h��\=���84=n=h=�E�;�&��Wмh1��#2=�3�IҊ��5=�HN=�w/��ᦼ1c��.�"=�Z��nϓ<KK@=�;�r*���=���;�m<\E=�
���=�����)=ur]=�C�Gт�5Z!=!=�=���$=�F�<��@��	N�ge<m =x_�=��]9f�/��pq=�T����"�(�<fR��N�Z=pj����h=�0�<v5���!8�V�J���ּ��;�n����[�W,���<V��pl���9��s��Sp���"=���r��<Kg����2��,�Ex[=Y�{�
K=�y ���<�5j�#���ݥ;�=��<�e=`��;?�P�ބL<����D
мw�7=�l-�Ϙ���<�:l�v<Ä�<�UA����<T*�2=^=ST�<�M �X-=(��<���<{u':c�&�����y;H�d�f?=Q�Y���8�;~�8�]�=?�0<J��<�>�� ��B�t=��<C�=���=�L=���<Dڈ<������Q<�W='~��*�8=.�<1�9�z#h�R�D��&=A��=��ڼ�~=}VT<�Y=�D�ѡ <$4=�=)��<JȘ���A=R_�*�Q<j#<#'�; �5�|yC=�Qu��e]=ݷ�<��x=h)����lz��!��IY�<�����]&�բ���ڼ�ZD�܁��Լ?��@��<V�<��l���G���F=鑈�i�X=�
]=?r�&'�Z{�����p{?=~�<�����.=�
P={��<e�	�k��<7��<�[Ѽ{Ο��v=:I���p�b,=߻y;5-=�0=��_=�n-��V���Y<�+<m���,���J�n��c;�Y�~<��j=40�<XB�~<�
/<��+����ٗZ=[F��n��㳚<5B<���W���}<" �郖<�/==���� <���]�H'I=��V� ����=��� ������ =~0��F5<�o�<_���&���._��}����*+�=�?B<>q$=��,��H=�0AD����<��ϼ"ߪ���r<>JH=��M���|e0��{<o1��~���\�)�=�2�: b���<ыt��d�=
�F=K
�<�_q�a�&=!g��Hǔ:�f��o���-=��Z��_q=��<W=���'=��U=gy;=jՌ��휺E�i=ꭊ�8 ��漲��:~뜻o�G�<Ħ���'<R�0=R�k= nݼ/��n`�����<��`=J_�<�r�<4��<T馻�O=���j�; ױ<�N	�����ڋ���	=�=�'X�d:m=8��<Et;�ja����˼􊍼�~��%E�K��;��<*Ss�R�\�,�����<
�% <�<�&J=��r=�Sмӏ����<|�Z��j=0"���:���\=V�<�2F+=�=2]���1�g���)��ē���E=5H��(�<��Z=�2�<l�;ņB=�K@=ߙ�����A���C���G�/y@<���ڱ�<@����zi�aﻈ,����<@�̼�8M��H=�/=�ۼ��<i$�q@����=���<WƱ���X=��<!�.�B'�(�E=,B=bL=?�H��g�<A��<�+<=�]��{U=���<�.3=����˻��V=+wJ=�#z���=�%.=|�ֱQ=VB�<�)3=�� ��g�,�gr=�e��Pȼ?-ռR�*M������m�
5%��Br=[AF�<�c=�ɻ׃�8np��=n��%�:���������=b�޼���N{�m�ӻ/��!�û�0:�����������;�1u=e�r=0�l��� <��;�=��v���N`$=�Z���Q��p<��=c�=�����;�=&�|��=i��k2����8�����O=��E���[�f�d��GO=��<�}[�|�y�)�� ļ�*=�	����;O�s�5���<��k��	1<��5�@�w�0��<W(0��l0������<=���c<���c�<�<o����K.<m�'<l��<�6X=v�<D;����&�e�E�eO~=�Q�<�μ{UA��.
=Ѡ:=CJ=��n<�4]�⦥���L�A�6=�o�<<�Oi����<~H�<-.=����fE�<����'���<��	;�zL<!����<�4�z�i�<�a6��[<�E�ڼ��L��iq=+$(��yR=w�H<C��<)V<`�μ�<�F�<z=�;�S�r�A�	Em��K�׿'=\�=v<#XF=/d�d5=M�"=�=��F�㉣�o�b��G=�Z1=oqt=4�<E�=��Q=�W6�\����I<`���k����<�s=Y(=�t̼��,=� B;)88=Uk�;v��:`��\��<��=x˨<�]h=B~=��=��N=s�׺�W=�wp�!A�<���<i*ټn'Z=n�=F�"�) ⻉�<B�[=9|3=]+Y=q)=�����d�G�8�[,��N���<%�;��=��DӼ:�<�+*=��;���<��;]v�;V��<݊�D��<���qK��݅�MN����<�J��?�<QU=�t�<��k=��]�U=�(û���<0��</�u��6g�7�o<{H0�L=}�U���D�&�<i՛<�t�U�=o�r�=��滬c?��:��l���.��� ͼΛ������<��E=�4,=~W��5��<�6U<���<�U�3#=�R����<�ݼ�J�<6�λmY�;]�7���f��=�rЖ�L�1���!=�v�< y;=%�� �6=�`�<r�=�<�⃼�]?=�p=��7=�8R=�1 =%	8���/��>���*�XG�'�W������ ;�xD<� <N����<�=�a��������<�M�<I:�<) �����<��H��O>=��K=�Bu�%0�#mT���<l��o�5<��H=��A<n��<UWH�EB{�A��<���{d�<:ἂ����x�!��*I�;n�r<o5	���<�����b�:� =��#����<O�<>R�<^Ǩ�r�ܼ�2�ﯽ���;���<�=��i^�3��1��<{5u<�_T���i����<�<u�!�[4���B/��Q\<벭<c�����Gμ���9�X�~.��R�;�K;��	�%<�a��H���-���?��k<�m7=��;��ͼ�Cg�;L�����[o �/�N<5����2�<�<=�%2���0�b(０fX��o:�p�{�:�4T���ݼ���<�q��㋽h.ܼR)=;;��Q�����<�<L�l�_�K=G�߼�V��hC<m���q=)A�;^�:�o<�@���|�����;u�+=�=��g<��<i���?=X�%<ֱ�<D���)=��7�D2B=�;���މ�ʆ�v��,Q����D5<ɣ�=��;=��P<��c�oon���缐I�<98<�9���3�<Y�'�'�|��os={C�<E����XB���{�@�=�%<K�E���i=�Z�<M��v�=��<�nf�z45=�M=�e¼�VѼ��ռ��;�s���چ�mۄ=�|R=���;W	>�����M3�<N�<br��0=9��߼t�8�\]4=�a^��q�<.�u�k����������E�@�����:e�/=�f�?[=�?X;�5O��O1=���:�2@�?���.�;=���*�
���ļ����>ת�/� <����*H<���=+�ټ�0���Һ��k�����m��U��< �B�<�mJ��yQ=�&V=���v����;U4���
=^D�<t����5=�}��<L��]=��=�{|<e{�;tD?=F�üC+ <���<w&n���0=�Y��Mb�t�3����:GQ�,�����2� �ɼA%l=}�=�X�<�Z+�x.���;??C<=G�����<io=:.�cjA���X�+�b�8&;=ş2=���;C�%�#��6[�<M=��H=��<X�5=$%���Ĺ�K=l�<�x�;�>O�L�U��&8=\Z=�O���,=� =5z=�}Z����~�]�2���b�<s��;=L�*<�$=eΓ�y0v�+�V�����8鼒�N�2=M=�CR�5�&�i�|=�=o�IM.=�z����Ӽ\+~<5�#�2c�;,Q=l�V=�I �eF�<�	=��=�A����z�YjS�/9=��X=rY�;�S����c�=�z��aE=��.��i����<ñ�<��d��#[����c�:
`l=b����+<iT�%�!=��Z;~Uu=��A��\=Xd=�_P;�֍�|�����;�� �8b*=�<R�W�P�N<��<�A=`�=}/�<��ؼ�̙���;=�����9j=�9�k0���w&<ڦ.=t>��p ػ0�	=k�*=�O�q���5��fx���8��K�e;&�1=&���	�<\Ǽ��ͻF2m��g�=,yH=&��:�M�<5�D=����߻Eq�R:����<=n��J��]R�Z�<�����<�hT=3[�9�Ey��Hc=ۥ%��!=@�_\��.�<()���S�<�P���k�?�z<=��D��<�n=�̊�]d�<�[e<X`==n~���0�~����S�;!G��-���!�4�6��G(=Wb��� !���t:s�<d�9Ӧһ�#����������M�=��<:�2�!���bC��6���*= �Z<6�"��g@=n�!�xn�ъR=�2=P�c�(�<�={������'=�=<�:V�=��;�}�<�>V����|F=�:;��*x<��߼��7�nl���
$<wǹ�Y�<B�f=�h�=6ᵼ������!�L�<��=EA�;��	��1�<��#=����;;_���ռb��:�	=h�����88��8��*��J�5�ꙟ�䎂<F���Mi=�I<=K���vs=l��<�e@=�����V�0߼�Z�<�Q��zn��v�<W��ncؼ�����Ĭ����hƨ��P��J%���<YW�<i�k�e�::�)<w�<�!�<I(�4��<�槼�M=0cu�舼��5��<����j=��=�Q�=2�<�Y�;�|��<)�<�LԼ/
r��;���a&<.��<��<�����=9R�<���Y�P�=�3�/��!1�(�1=�O�{�����<��c�TM�<��<coY�!�:L�<��U����<H�O��#��-�P=w�<M�<��7iy	�1h���<iټ��`=��_;X%D=|wL������O<=�x��L=��*=
��<(�.��y��������hh<������C;�����<���<���d��fe�g����<��<�Y
=���0�"<-�=bT*�U�e�����b���/��C=���;dW=8�=�g��*TK�a��D!=�*>�[^�<:cg�m���u(����5��(y��O�5�7=ݱ=�������'r=��;rP�;�%
��L6=���<m���K��TN��5�?<{C=�5N���-��<o =gRG=f�<,<PS��*x�S����i�=�_l�d�f���`�o]���2=�3�<�=���<y=�"���@=$~�#/<����xO���:���<�[};�[=,T��q�l=d1{=��=�K���1=5x<\����o��{7= ��<�d��Q���ټOU߼�=��; �׼��<��I=7>�<2Q=��;?2��U!�;~�<���<�٣<�t��U��s�;��F�zi��A��<Ly;=o�s;�h@��Q=��`=�w��.�<!rc=g]=_�9=��O=zpR��==�g�h�=�{��q�$=1|��H.=�|�;}����*=\3=|p�<˦.<ލͻ
e*<�I���<��;�כ<�=�Q[�?� ��=� ����<���<��;0������F�4<:��<ѕ���h
���<`a���1=��:���c�Z��k�7��Cһ����8K<��j=���:�H=T}*;4���G=�ǃ��_$���u�3<�Q=�R=�둼�F<�TS=�+F��B)<�C�M=��V����1��U�i=
k��
!=c�==�
�ȉ3<��p<�=Z�cWe��*%=��C��Ě��5�B�@�خ��=!�sV�T0�fB�<P��P�<Ð=�Z=�U�<�r+���7�g�<ߠ�;sxV<Ө�<,d.����<Dr��e%=�2�B��`D��w�����=��p<	�<�2='S���4�<�o�BE�xF=!B�=���x��:=���:C���{=�=/!���,�<wz��*�P���6=e0Ҽ��� �����<n�)�}w����������;����^����GƼw�~<��Tv"�<|S�1ļ�*�<�
c<�E}=	9�F��<w�=��~���<���<K��eP?<'A��=2�'�eӞ=���<(6���L��LC���N����X��< ��9�]庴��<�����w=?�� ����_=�=��\��=��缥�4�I��<o�r=cuf=s�ؼ����9�:4O�<Y� =������k��+H�[��;'���eg��h�=���;�%�����<MF=�{V�,.=�^>=�@�<�/�<��t<n>-=��:=	S<���<I�V=���<�ͼ���<UJ����0ݲ<�J8��r�^����u��h�<T7��w��]a�;�[:=|��;�M��1��<(�켕c��s�;@@��/��\ ��Bf<��k<{��[�!���<�O5�흼�0O=�v==�U�;�k}�S䞼v�?�#�7�S�==�A�xR���M=��=�Q/=0�;;�<�w���<��4=kp<X�:3�>(��aZ�=����Pռ�>��rB��$=b �3�#<�ϩ<��U��x �7�w����r��<�ag=i�����<8Z	�8�|=�U<w�D���_=��=����nN`=���<ݯt��̙���<�>���rT���<C =Ruμ)���:=��̻��D=�U4;D)?�O�X<*�9�����r�<̡8<�ME��_�;6�=+���݀V���;;�<	����8A�N�=�ռ�m���O�<��S�j{=ȘC=����Y��F�6=1H�;���/�&��g��z���<�7�:ވ�<4C����;��<{p��ƹ����<1O��K�T=l�=¬�'R��푼T0=mK=��	�@��r9=G!i=/D[<���{��d��<�����|=���<.L�Y7"<�6��:az<p<r��<,�����<%��=��<W[<���<G�咝:^��gQ��fk�2�;l>�=bB��k|=��ɻ�5�<�s�))�d`���߻�e=.��������<�C=�M=�9^��5�<YL<+d?<Ɩ<=Is�v%W:b!=���;��M��a=�lμm9Y=���<RF���܈<� J=�
�:�# =������U�`=��<:?������<=�Q�����<3h1�� f<� =�``���v=���@��ʪ2=쏼��?=�8P<�����o���#M=-�R�d�=���<��a=�O=��	<|�<�6��;��/=eH=	�l���;�&�<o߼�׶<�O4��3��|��4C=�3���,i=��`���>mۻ��3���9I.=)��5�� <*1<�ֻ�M=�r�<���<	�;:��<� =�*軣�I=��="�=�P��y�I= ˼��s��(�-H�"�N��q�(�e���_G��'���¼��xżtes��%��Jv=b��<^]o=��B=v4��&=l�<�vE�L���J=,���U{�=�=u�X<5J=.�0=�0߼��8��<��3=Q0=�-=��B㨼qO+�ɯ����ɼ��=	�<���=�/������84Լ{��oɑ<�چ��`�;N� �0=��л�J<�N1<$<�_A�;6��ߦ;�'=���<�g�<�F$=�Ӽ�~V=C2<=t�f=8FZ���@<J�h��"<��<���Z��<�Y�<9�G��\�Q�"�;�=��A��A=�����k=�I��P,=��R<)r=+���,7`���v�B�C=;I�<3��<d@=�L��=*�<=t*==���vK�K:]�[���ӍZ�v��<(�=1��*P���L=��=��R=�v=w��k
���'C<t0<+�8�H =0s��09P<�z�={�+=\삻]_໴rG=_{2=��G=1)u�7AS:��f=YA<�:�;�z�< =�v=��U=���������<��;�����:D&�w���(�=��<���C`�<�B�9koH=	��̎^=�2=�=��%;Al�;w�;ٔk=RZϼ���<��N=��=�N&<�W:���q<��<z\t=:M��%��N!=�Rռl>Ӽ��O��u�u�1U�� ��]�oD/��\�\�=X(�<�S��R���&%�R�9=v��E��hL<J��<h����ZD�W��E��m�*>� �[=�:���&-=���t0�q��/<��<��<��<�eg�k݈<i$-��"=	=*=K�;ǤV�*=nI�<'	��#�;Aw�;Y<=�q1=�#=!5^�3��<$4T�s�һ����k
�<t�?=��j�93F=�˻�=v����:�]<�v� E=G��L#�;���=��2=���|[=�O��F+��8�]�@��N=�ߠ��-B=3B��(�;�l7�R��<����2�@=`D��+��<��=��=��O=���;!b=�^=� <�)��u��=�K/�������
Sü��.���%=�����t%=2�3=l~%��d�<�h�<���3�;�m:�0�TLL��Wn�+yB��G=;�W���w=���<}?=d>=��@=��T<�y�N��@�,:!=-;��q�'!�;+�'�2Ĺ�H:�;7Ta<h��<&�G��u�<|ϐ=+��9弉��:��<�w���R�]�<o�S�l$>;�+l:�J����J�g�� ��M��;�/Y��=&S��HK����<atż��;%#��~#�5��,f �T�����;=���O��P�,;X�9L�=�ʬ<��<�*<�<�ri��	6�p�*���<�Ҽ��=��<��!<F�;Zf�;��A=�:,�	NG������h�%��W�/=�a\�E#h<�t8���=��==Y�=��=Lc�;���<�TM�9{���<v"�<��<�'�5a�:p�V;}��N�;�ڢ�ۭ^����:aP{�����ƻ���t�L��/7����_����.<���<�(=Oe=�]��=��g��/�xT^�J������� :!=�.<��2;LC=��W;!, �D�<��=_��;J�l=���<���EcʼO"�+K�;��=�:-;�:]=��㼧& =e�$<�a5<��]=&��< �x�My0=6���Ca<�S�<i�<=��<6�n��[�<�ٴ<&~ػ�����=�@7��R!�d=g��<�<��/=1�G��Y=�?����#=�c=�
b=�[<=	�_=���<��3�_�H��܉��$
�/�Ż~�{=N����K=͆Ҽ�0o��a.�&Q�<?ʉ;��<̷ �&�m�>H^=$q[�q,b=�R��#D<�L�<�]E=@1(�mb6���4��m`��_���?=��<�9�<�Ǆ<'V%���ND=S	���=u&�Suh=�����^����%�m56= �l=��W<С�=���<9^�?�a=��<��*=��o=xZ�%�o=����*=Q������	X�#-=�%B�H��<�,���`P��U�����2A��&,9��a����d�輬Y==TPl� �==�$�Ȟ����~=_x)=�v(=�,��c�<��ulV�:%m��{�=��=6qd�x������v��^�<:N6�n��;4J:���ԫ<���<����G;(��<$m�#Rp�[M���C=�;���;gZ�� ��R����*��3=C�<�0����<.x�<��
����<���<o'Z�s2伒&������P9����瘺�6�H=��y=�K=�=k=uH=��;M˯�����B���=��<� ?=W�=�4)�Wh=���<��yA=�d��jF��AQ=����7�<����B�a=��n�1i̼�l��yC/���<_�@��	����ϻR��<oҼ�*d<5(�<�|3=!��<�)=���J��<D6�<ŪT��%�<%P�<�]�;�#���G���H��n�<�д<�9>��Av��ְ�?P6��
]�����lD�<�4>�<�Լy�<&N�=b�t<'�������� ���=
=P�5��l<ƳE��	/=�C;�_j���$�G=�N󼤮���w6=�X=�=mʃ���p=p/�<Q�E������:��
;[�]�V�/<�o=7����@��c|��@輙 	<F�T�~\A�_�Ѽ�k�<Fq��;4e;�Cd;���<�i'�e��<��9��I �b�[�6�<���3��������G=p��<��=���NP�<�#=�`h�c��3�<L\=�x7�x=�..;�r!��` ���%���4=����~���<�4漾E�8xlO=d_ʼ?G���<�>��=2�+=~٢<�����=����=:�k=�~4�wɪ<E�&�B�	="ǼJX1�;r�J��}�D��(ػ<�d���|N;��l=�a<Z�;�WN߼�T$<��ƹ��<b}�<sG=��ӛ���Ѽvf=g�@<��=i ����X=�	�X����0=�q�<B�0�I��;�O,={G�<�٪;+0^=x�|���<��<�'=5Ǘ<����{V=�N�<�N=��>��4=�G�#�%=&�<C��<+�<��=W�U�;�-3<'@8�^uK��"=/�O���[� o}��b�s4���{���<���=�n�C�<�{2=5�H<��F=�D�c/N��d�#����y"=��;�C=�f:���;=� �%�ѼAꀼ��a��\���<�<���>��2S��裼B�J;%YN���;����������;���=����l��;r༢����3�t{�<ɂ�<�?=y =���q�d�?���q�lė;#;���| =s��*=�e����<#\M=!�u»�����<I�y�;�[�;ׁ�<���֩&=t`	9~�)=#ځ�5��K0�<��=hG�_W<rA=+D��(JO����:�ܻ;�}=�ڤ��E��5W���3�����L2/;�*�;l<�F=�2�3Ӻ(�`�t��;<���c��Nɼ�/"��X�<��;7�M�-�C���->����	I=28K�ٸj�Od��Y=���;���n�R<>�.�ȧ<�	�f�L��'ӻ_�4��n�<^x��s\<Z]	��|O=��+=�t[�L_;����7�&=��	� Y�;�Nż��?��%,������i�x��:A�;U���
J,=�Ę�Z�P��@���a�UV<h9�-�Y���,�==&�u��t�<��/���;�i8=�V�A�<Ի�=��<��7=��*�a���r�:�:p=�:<Ҕ�;�!%��q<�� ��f_�Q*�=�G7=[Q&���Y�ڼ�;6�N�2��C��<�􀽍�j=xy+=��o��y�;ʇ�k�)=a
�5,=�� �=r,��l�m���м�]J=�� =f��y���<�)<�󴻐�R��oW=�Ԥ<�H=x�;=��=�~��R�=�.:�Rg{�݂)��%�<���5��<,>|=�* =�L�<������ɻ�ݼ���<�=�=qW<
_�	wA�>�׼\�c;�y(�c����ļ��6�{)U=E�=�5L=)�<�լ<!n�f�`<�_�!��ǭ��/)�<f�k�抑�I�-=D���S=��/=��ʼ���<�E�;G<=�7��c��mY=�}=�]��᪼��8<��H=������F����&I���V=JY:�J3<'� <��<j�<=ʎ5��<���U���;�����$=�{+�Ѧ#�9z�����=��<�[%��4�<u�����<�S�<d�I=j��qn�<PO���9�Ⱦ<�E9��u���XK�^P��y��<�D���N����<��<�ػ�����<g*��}d=�Y�����Rx�<�>P<c��=���#��u����<�E:��n�<W�$�������E=�V��� ���<)tA�����)�P<�2�1�O�Z�:<��7<
�A� ��<l/G�rx=U=6���X=Y{%=E΅���Y=�Z=��ۀn� z�<��<o>�;�����h=�a�<�<S�F�K3b=�uټq�<��=��E���w<p���i ;o�g<*�p=@��܈<�gl��e<�'����x<XW˻y��<��v<�i>�7�;�X�<�[�<_Gp���(���<�lػ<Y<�[��������;�=�<�:�<�j�H]�<����}��;�"#��J�<��\����<��s��P��I��U'���_=��^���O=ӧ$��8�=E�!=�E�p�5���弽�<��(�?g;< UP=��i��X~<2&-�)�����<=�:�;�7�/=I��<��f=�-e=��W=��6�V&��gҼ@�L�biE<6�-�O���*��z,���;�-��nqU=��_="��<��]�q؊�fYJ�#�<g�μ55��"����<c.�<�\���"�;Ve&=W"�.���y�8_��p[<���<�}�;�9=_/6��Y���%��%I���!=����������[�I�����ռ����z�&��J�<*�k<�,��GR���2<��<'u!=���<��;=9����<��=ޒ9��=%���=���N�&D<m ;;+]=l�;�G<y�P=���;��d�3='=����_<B��<Wφ<��=:�J=s�.=�H_<�e_�}?���v=I�-�.p����:=�Q�<�v򼰊Z���D�W{Z=,��<P��j�8�]v�<�' �fD��Y�C�@d����==1�3��٩<N�6=3�(=t�A�I7��G'Ҽ�};�\=-��~Jp<ӿ&=}��<3�����<����c���[&=�4�&�<�5�<aG=���L42<H*b�|pM=]ڦ<-g==�=;�4;&�#�<8m	= ��Z^�B�j�/=D�I��P=�&=o�7�����#�$�V=�.̼5x�;��ȼ�˱�8��0=�>����ʻ��0�|�̼'��<p�;��E�h��<A�$=��=Tm��|;�ԏ�	�Q=��<�W=�F�<UN=�p�<V;��o=؛H�cP�y��2�.<�# ��)�<^�W,O��C�"&�o����= �j%:�zƀ=9U�<]>�����k�;��B���={Z=~�:���I���=�Լaݻb�d���<����#��u=��D�v�X=>(*���=�9�����<V]=,�<�"C��R�<VXF=[�&=É�<�����<�黟W[=��3=��<�����<�,`��� ��e	��<1�;��=_�}='{�<}�X<�O�]�/=�W��S�3<�@'���E=ޮ�<a}<hr���}�Y=ap3=�<��+=Q>�;���7�<��8=�[+=����:>=H��9�l��qu���b=�|�<Ao=A/��r=j�����<��]=�Dy<���;�J=� ;A�F�O@=�%(��%�n���DP=�c��ڣ�<�4��H��<���,��<�cü#=~=��<��C����<�빼���<vG�=�5#�ķ!< o���<<�h=Z{w=ަ������R��:�+=,u<�Y�V�<wK=vV�<���<f��=�{{��(t=GP=��ѹ�	 ��ּ7�=��q¼��2�F�鼈�<�Tn=��w<��
�]W?<t�<!������*��o�0�ɿ%�巼Ը��v9^;�@<�@=֮Ǽ3�l�;##=?�(=���<�Y��������=���'<%��͹��ǤE=�8����<�����<����*�ʷ#��:��<�=0<p�����<*�;��{�g=)��< ��x�<�VF=@%H=�s�<�x��!=ӴN�.qU��Wm��W�8B�<���
%=dM=H��	<[=����`���w�+"����9;n
���0PڻvcC�����y.<��Z�.0=	bH;:v=舗=A+$<��t��*\;�T��޻|��<�݈�]_6���<��7��OU<�U;�0��冼����Jf={�];�
<~[=+=z��dO6���*�k��^�;<)ԼE�=�B�<�"��J�h<�R�9���I����<���,+=�M=��ɼ	�=h�8=�u{���������]�<I��0�;����tn�<T�<zL��(��<��9��h�����<�^k=� =�c=H�<��<�:���=�ET=7Ii=��(=d�ݼ$=��g�gk=q,@=nOH���*�j(��!Օ<��6�L��<)g�<N�;b�>�@m��J���bv�=N�՛>�7��;h0�e�=}u�=��<�8_�V�=HO7=ro��E���.�<��R��}�<�G;<+��10�=�=��%� l�:XF�; 	�<E�<̺Y=� ��?�<�~�K1-��Xx=bhY��'���<ۗ����p=�T<�'h:�r<W�*=�T!=�<;�R�Q{=_~��ف=Z2I<�=3=Zʼ��<�N�3x��z
=T7<����0=W֮��C�<���kļ��q�<�ļ���^F,�'h��Z�B��<���;�E*�����,?�;#��	 =cX7��7���F=H�z=�I���C�<�-<��k�)/̻��p< �<�؝<��^<h�I��'3����<ݪ�<�B=yF-=.�&=�p�;�r6=A�λ�=_�k=3=�ap;�y��=u�=p<�3q=z邽�/8�6��`��<x��Vl6���ʻ��^=]�?<�A���$���ռ혍;0�;�;RG=�*��3A�u�=������;(nS=���C�<����+��}�;)=jN=��I=Q���w�T�ާ�<,R�<�=:7=7fv;P�=7e��d*�掻o~==(0ػ����?��$p����<ⴢ� ]�@Ԩ<�n��z�=rne<��	;�{O=�8D<��;>:	<E)q=��Ѽ�Y׼,,c�<���ۍ$����;��<�N���G��t��n�=�o�2W������=Hl<��=D:im�< �=�M=�T�<%L7=�:F�<�JO<�ټё��x�<� ��P=r�<=:m7=r	���6L�G�o���$���<
�F=5#��^�.�<�ӵ�k3�<�8)�h�L������<#d��e!&������%��K�.<��O=��;S>3�d�)�u'x���7<����1���ڼ���<����2�j�N=�s��|𯼯I�0<���+��@n;���]W=� X<���O=lv� =�:�r4�B�~=�\�<׬���w,���A=E��]>X�k�G��K=��'�+��|iS��y�<����2ꩻL}=Z�I=Ի_=�2=�\�n"�<y�� ǉ;���K=�ㇼޚ.=ltp�<T�<��~=?)��So!=�:���=H�H=R��z�<N�����<��WI��y@���M�|��<�<<���yz=<q�����W���<�� �P=qt=^u��ÅG=��==��;��>���:O�<`@f;�5���� =Dx����<�5�l�#�M�4�Y�=��S=�����<��=^T=�k<à
��۔<(Hx��m�X<����@��&dnf=�)c�T�?=ҬP���'=T�ݻ��ZFa���<8ͼ��?����;ֺ���D��� �x"=�D�<p��=�،��t �W/==<�G�O�������Q=2;�;���';�,�G(=B3�"�a<3ϼ[-���;�½<�u����<��=N�E=l�N7�;gY=��=n��<�w���N���Q<�A��Nm;/I�;�Kc<�j�2��<�ŻM���i=]Gu�0����<=�o�+=m=��Z<\6�8 [�ܴ6=�4V��0=���N�D��
�����z�;�;���8*�v� ��%<�Ns:r.	=�:<��(<������=�=.��<t 6�=<�O�=�Fd=$r}��|�<� ���搼�����ц=D�V����47E��Ƽ=�4.�T[#�Q=�1�;�-=^�＼�
�-�5=��<�{rM=�~<Z��
��Pۼ�;�Ӭ;�<��ϼ��]�A��; �=�b���L���޼��I=̙=�K�"+��D��<*~d=�ux<��9�Z�B���9��Z;	g�9
�-�;��<�l!��r,=��H<(�==��
��e�<�=\�r=)@=�B=X3����X�#{=�Z=
ݮ;Fy<G�f�шD=�󚼂�=G��� 5��؝<�'=^{V�AQ\=�Pv=>vm:�諼�[=��,=t�=pk��;��z�X=�<(� ���<r�9=h�=��;<�����8�v5�n���a�L<�*2����<�] <�)=���<Z=���<q�b��RV=�?::�X�<a(=b�&<������;��J=,�K�����U=ͤü����#����O���q�b���h�r9�8>=��<-�$�4����6�=e�=�E��ޖ�<�kZ���<�M~<�Ǽv�H��i��y~U�Z*�;�=]���+�<��@=�⻛H:�"\�<(���z�_���*=U�<t���6�<�(E�+熽s��;%�<\�"=Ӯr<� =78�<IM�<b�w���-}���]�JÊ<��h=i������� =�:�8iy<09:��
�:��A��dm���?=��<=%{ �9J���	=h(=<���<<���S,l��E=�h�	��<C��<OI�s��R���b,���<
0����=���u+8=>�˵�T�ϼ��f�XAy<��=�v�:q6���G<=�	=?���[���r	��0I���==([=PF���\=�\k=mv=߶��v�T=y7d=�<�{�=-���$&��r3=7��<�S�ڿ<���s���K�ټ��+���$=uD���<��B�qP�����f���d?=�#��H5=��-=�.�<��:=�<�u�=T�1=3��<f$�:DY�<-����g<�p;=�T��=�G=Cy7=u�����'={�h���m�T�LI�=�+�<�Ҽ�ބ=��a���L�'0�<#�<�&�u��;s�<\9?���m�UWZ�"H��Z��\(�y/�1==T7=��<P�Y��FP=!�.<&>��X��q]»�D�<�?��?/=��������j���=I�I=wl<]'߼d=[{¼?i���G�P<�A�<xA��
��Q���\-=��D<@�<���<�,�=E�=��9��A<
�<J�y�N=�Oy<$��ok���<���UF�zը<�׼��w<�d<I<���]R=-4��3\f= ������������h<��;��;
bf<�{ż��L��[I�ېb<������=�i=� ������;�o=�"�<�u�<��=�Ba<ȟ�<��л��<�;�<W�^=��E�@W�C4�<"��<%�C���:=x��9����ؾ<V�<�P=���<�9���׎��Qc��ݗ���X���
�<(A��5c�A�'����<T�C=���;~@�<N�9=���<?
P�f=�����]�9Ֆ���<�W�<�-;��wz<r��<�X�<a�7=�N�<��/�M�ؼ�c:=tiջxB��I�P��n�);j6=�!�<G�Ӭ���c��<v��b��=1�ɼ��M���/=�%�<=��	Vϻ���f/�<�s�<�s��Kb9��(��w��<�`�(�Q<�R�R=l[e� 
$=剄< '_����<%��U=�ʼ��=��3=��<���<�\=I�U�� ��zG�<��e�/a=
R={���5�=���</�[<yUҼ��<)��<�9��e��<�Ӽ+����2;k>I=�o�<C�7���;֥P�V����=��:��t�;7n��L���Q�Y<3c�w! ���<�&{�<��j��=�@�o��;Gc&<�ᒼl��=�=@=�;=�)<AJ=��U=w��GV����<ʩs����=�X=�?5�����N�<>�q��?w���;�qA<���"�<��U=E`=I9�<��-������Y�y;@��D0�%����f(��� �|�;Ob=�Mi�gf=Q�=c���ռܧ;=�K7�+�=î8=c`�<�;0��=[qV�=;V=ǥμg�W=Ʋ����~�w-B��7����<@cI� 43=cȻ�$NH�l*��A=���~�a�!�,�N:'��7<�S��{%=;�E=���rv��6<T�.=*�=�Nu�d=N슽ɤ1�֐<\Ȣ���;@�-����v��<�]��R(�0%�<ZI=�\�<8���U9<�h>���@=������ =&��Y�Z�M��wu������r�V<�B���l]�LQ= +�<w�<�YM</�:����G=��<��=��<��L=O�h=���<�u�m���E�=eN�&��<��[����u�*���%=1�<�����2:=[�;��d�up~�0O�y�?=6ؼ`i.��ے<�<׊<kr�<��I=��<{$�k���v�K�Tz������'�;�E����N8��{U��}8<��P<��<�ɼ��)��Ա�q{B=7]�< ��z�k���޼%X7����<�B1�1%\=�me�>=T=��ټ��e<��I�8f���J���u=��W=���!ԩ<c=)�ǻ?ί��,I=1 ?��j��ռ74ؼ\�����<��'<ۻ�=�Vj=�gw��m=�Oy;<LX=57=��߼�P���<"ڼ�:=���:a����ۼK�<�t+�P��p�ļ���<�-=�Hs��R��u=M�7:$Б;�1<=d��<A!�<��<R�_=�H���0�������<R��<�l3=TJk=n�Pi���J=����=&.j��Cn<��)���<䁽��Z=�!=�����|<z(�<M� ��A輅�=����T%=�� <��<�9���<��v���a�V�l=M�#=04=P�����X���:�Os��DRQ���[��S�/6�~P�diU=��$����"�J�0��K�(=��m�<L ��f=n��=�T=f�U=�0g����1Fr=�*��pXG=��K=SG��1H�=.j�\	=�S<��E=U�<w�4�׋!��wy=���e���$�=��L<B#^�uE�&)h=�Ƒ<�� =��'��	�R<�<�ڟ<A-H<�t2���3=f�o=a�p<��'=�E<��s�������>�}��q��ʙ<�21�fD=d�!�O��<�~Z��zϼ�\=��Z=����$����{�	�<b2/=��:=�7�=;/=m�������lWA���6��ἆ�R���A�F�P<+HR=)�<�5�2�(�q;�u�w�n�=�˺<f��;��@�D~�*3�<���bu�;��¼�X�3�=T;���"=�C���=��=�[>��oT=�������;�*+���f�\f��s�S=t\�<�\<��QY�9 G���i���W<��;񚉼�⌻m���(=�(e=bY�<�Z<�\�<t�F�Z�\[�����
F���/��g_<��[=��:��i9=y!=M=�L\���(=J�<�<==�����<�dҼ��<Qծ�|DR�{j� 8������[�<�,=�y
{���(�bݹ�>��:[.=���'vS�S�D�DA�<��"�J���
��G�;h0�:���Z�<j�p={|��t�<E;���g<+�����lgp=(��>*�� �$<4�ἁ1��B�#=��;�%����==�|)=�5c���L��T�#�.=�*�����=r�=<FA�=��:.��;8�|=��=��_��K�;�c=�Q�K�U����V;�m��Pf��n�%=J��;�R�K
�<�7�<|l�<A;<s:����ֻ�!��Y����C�<N��P�`<�<*E��f㼚��<��<m������;���;e�q=Kl�]-��N�Y�j
����PN�<.�7=��<�r���:�<��)=!���D=�]n�8|-�����!�>Z���&=x�(�`�T�%i����?:ˎ;�#o��O��4�8F=�n��K���<�b�]�:�և���$��$�1WI<�o�<�=pK��F˼��.=�ᙽEI=��<���Rn@=�o�=aW�<�;�5f�(���h�;��\� �:��u�M�!��ƽ<�<��f=cܝ�,A8=-=M�z�,�_H�<D=�fӼeS
�����<�C|=��<${�����=!X$����=-3�%E�<�NX=�,*�1���v�r��\�wA;��>=�D��d*�<��t=�S�;i�S1�<�,��̫<��B=k�f<�@=Ð9����8�Yi�~l<zS=i��աZ=8��S7���V=A2��y��0P���j�~�Q=�*-�x�=<��;R=�[=�[�l�D���<��:@��;�d�=-��<bbD<{kA<�3�;/��<7M��f�K=���w�v� ��<��<r�a=��;�z=u+E�$�&=	/i=ꥯ;~�G=	۩�ܴ�<F�H��<�D�X�����<E�=<ڵ��ҏ��=C▼xi�<���]�輒�켑'�1(<q"=ߪ�� ������<> �=��s<��b=GՌ=�μ�h���<��6m=i_,=�e�<n�;�,��Y�<�8�eI]�x�����;��\=S�R=.���<jk�;�6�<�=ǧ4����<躯��(�<�A0���J=�3<D��<ju<��G=���<��������c���.�v;�T�����ʝ-<}���5Ld�I��/�C=8}}=V����<�� =���%�=阄:%F�<��=��E=��:=��=�
�<��N���2�P̌��
�<�7����m=�3�,<�b=�T<�M�pּ�m�=��>���N�*$<�Ǽ���<��d=pl#=\�<��^����Y�f��Rw=�U����<�D��XǼ��q�T×�b�Ӹ���<4")��`�<n�]�f����Ǽ���<[��`C�r�P=4{�<�MC=_��<�-�U�㹆5Լ��<`�X��s0��zX�H�<Ѳ��H}4�Nd�����_r%��y�;��l=
�Ȼp4U���B�Y��W=�=��=�6=2�<�a�O/�<�6=<b3=/@ɺ��<EV��2�R<M8��� =Je��q-�+����<���O{!��Ǽ��=��0��\e~;�����C;�H=��<M�=�틼��Y=B�:<� <�Zr<���S%=/K�Ju�<�F��$�<r�����<ڍ=�!=�<��;���^�E�>�h��<�:[��-C���z'*=��=�� =���M�=2��K�ϼ%y�<�`�"�:=�=,�<����<�i�<�������<��� a���{�����Ǽ61�<��+��dg�ë$�C��>Q���`w�R�����μ��:�5e��Y����W��w����<�<�%��r!�<�gp�J&<�c��̮�m�Z<�*=b�;z�i<�
��d<}L��4c���K�<'F�<�O`�lڄ=���<Xs	�]��;��6��s����N��bW=U��"͆=��<4��<Y�=E�C�y�=Kcj=)�Q=>�=�,��M�V;��K<0Oȼ��^=T]S��¼��=���<�m�����<H؂��.m=u�-�N��M-g��xL=��"����;���=����>� ��m��?;��#L�xi-=�)*=��<��u���׉=�� <���˾컯�$<�`c=7�z<3�P�m=�5ż(=ü�:=�1=y�;��Q=���<�0p<������<أb���ۻ���=�
=�!Ҽ	�?=�;=�w<�N���z���=��W;�>��c1�pD��V�<��߼;�\��
�����O����<��;��<Z:"��
���E=���<�⫻��[=�+k��EW���+�wcJ=ym�#�t���K���=o�)<G���b��S��<ٽ<$ټ�=F~%�������=Hg���Ѽh�5='
�����G���[�<�A=�C�=t��<��Ƽ��<��̼2��=:%=���<�4�<,f�<�B��Ad���=�7d=�l�;��V�me�ӡ��W~=�7.=a3=\ɦ<	(q�C��:/Y��1fO�lj����&�<�I��s𼮪.�26/���K�8�r�*=�,="=���;�~Y<A�=��뼃d-=2~�<ة�<��Ӽ�߼?�9��TX<��<p*�Ζ2���J�\�4=KSպ���;o-0�ɼ(�&4����<�ׂ�)�	��:=*`Ѽ,���"=/�(=�Ż �8���=�Ѽ�|�;\�=��==�VF��9[=�P@=A�P��'�=Fr�����H=�p�?U�<�=!d��9�<p��<�U�<�lƼ�H�<�6�� ���<ai��˻�h��{;j�ٻ�IO;������Y���ЈZ<̭F�tܼ�Zͼ$�,�!%Y�m~�;��=�8��R�L�<'X=�3<�9=Ug[�6tZ=l\�<(�!<�i=M��<�Bt��ԃ<x��ǹ���'L<-,�V�"<���;-�[=?4���0�Ϊ��=�I���&�Qsr=[%��E�L����t�L<M�<H���K��OA=8뫼��"�}�ռzcR�p��<��T=�.:;�Y�n�6���2<����YƼ�[��$Q_=Ļ��^���
�!e6���v�;c:=�%��9�<VмJE���	�� M�<������ĺ�+=Z%�<k(�;�J<�:���4�P�<��<��w<2�4�Mm�=h�t<��q�����g&>�	�d��$�:f~V�̍ʼ;�j<tfR=���<c�z����ؼ��	��<��<��G=��=HY=Su�<����m>�>S�Pᒼ� =��=�?,��ȻL�q=�=��X�7��<�s�	5�<�h���%:L+=���<^��<��=Kǥ<$˻9=�V=ot6=�:�=?���yT9T:<	ļj9;�=��<�,K="�����+<����]������s9�&�L<!�L=>Q�<0[�<��<~Jȼ��wf{=4�p�%= =��X�
�Ӽ�G<��.�,v=��@�u� �r��$����<r�(�*�ؼʶ��C=��=�F�<Z���]=�Jp��⏼
�Dy�g�#;��=��|���'=?%=��=�)�<L�\���;�ݫ<����48��禺����."=�J�<,�;�ռ*������T�< \��^�$=�=_=��\;=��P�=4�o<��U=s�F=�-==�S<�� =�/?=׾�:��b:/`��f��xe�;U)E�<'���!=�}�;��ܼ%<��@�	����bs��]��<}7�=�%C<� �: M<��Q�����'<P�b=x1�<wCE=9E]���_<���~jE<Ws>��|;��A=n�q��K���Y��?C�C)-=j���Q>��M�K��<q_����<r�	�R��<|�m[	��$�} �lԼ��<�# =����!=W5J=q�=�P��Zl�!�ڼ��=���!- ��?��?<�޼��<6?���|��<��w=0�ܼ�Q�<jLD=�݁����=�4�=�n�g�=k@b<��;!/����<���;�L=Ű|��2D�.�d=�	<*�ļ���;�1���L���?=FB=�K<޾E���ּ�/=).U=6�4�T�=��V<�w�z�<���j��E=zҺ�`'�<I�<��=������q��(`=�dJ=��<~-A��fA=*K=�;
o����<Q�
=��N=�	=�x[�r0E=��T<Vs=��;���ռ�m����<�&��b��<'�.���F��^$=A�y:|�`=aQ�#0=$C���*<��W=��<+�)�Q'=5d.=z��;��ֺ���,Y���T=*i/=iE�vм���3܆=�a��}�XWk��'�<m8��/���e��hd���h��=T!&<��5�8扼�k= s^�rk{�y�a=6P���eӻޏ>=�GT<�>S��� =����������<&?
=kR=�:�z�;� =�W0=}T==K�N����ǼVCs������I/��-�<�P=��<�ؼS>H=y��<�e<<�9b=hb,���P=g�2��x�<��s=��~��d������s�<v�ݼ����?�M5�<�^<�o�U�;o3�<��7�^=��滹����@=���<�<G�ļV�f=�E>=���{$)��=����W�A�q������_�;��й�M������Y�Gw�;�e�< X?=��7<�^��;��<��T;�tR=��<x,*;�=Iz��{�2<��<�-�;��v=L��<���B��<�Ҽ��n=���;jQ�<�10����<�R=�<SW�;�� <W���J�˻D'=�g�<���<M�=�Ԗ�������`<���ނ�AR�<��M���7��#|X���4�*R�<K/���<�e�;5�+�H=o9,�쌜��:Zqu<����<i0=:�M<�K�;��;�v���O���%���=���<D�Fw�<�.]:0��ȘQ<<e켥AI�"u�<�vw����<xR��_��������+�U=�T���&��=V�Xg�;sLüsK���m&��e==ˌ:�oR=�_�r��<�2�</�g��Z�;��:�)
ͺh�Z� �&�&�
=�n,�W��:�pZ=��f�\YE=�����^��<i͆;�>�=�[��&�<���<}e�݂h��Ġ<��=�&�<�M��Z�'��|��7fA�kG=rP=�y��tͼH��D�V<��<��b�O��;O �;v�&�]=�):=1J�<y��<ri����9c�=<%�<�=�P��%1�s^�<d��P,�Xx����<�陼�$=�˶<��Ҽ��a��9�<���<������T=��1=a��2�<W�'���=l�`���y��m(=$�<��mK�ҥ2=��<��`=�8X<�S��j�⇨�Z��F�o�I�� ������»I���\�����<C�c�y6�<��^�?y=.�<�L�5��k<�D�`�<�Z����<Pt�t�(=��f��:��MG=�K�<��<��>=t�S=��>;�<�w軉���"w<�y={==�'$
��v�<�Ҭ�(�\=�%G<R�!=.�<�� �v�7�F��<ķV<��!=�F�D��;R�=R@��;�&�A��W=��,=�l� �e��@��
�;�[�<�`�<p�:H�^=�[�Wo:�WK��Ƽ�qZ<��,���2=8��<䫔��LK=|����0=es<��P�.2<m��<�,�Ժ�<�@��,�<9K<+�;%��<���<��#����<�f�I���3��<`4-�H�g�Ӽ`�O���X<��<b�J=�b�<RO�<��;�t�<�<��M=E�:���Ut2=(>�<�C�<mh�����I�8<���,k�<_�w��O�:�V.<̼{�;:��XI�<�7f�!�=���r����t=��"=VPX<���\�<�z=�&�G�*=z�8���;`=\n/=i�<���;��><8$Z��#H�Q�<N�-4���5�����8�2h�<�<j�U<~���������L|5=���<�Na�;��9q;�;�0=N��:I�v��[��m�lMe����;Ns =~r��ͼ�`5=ϼ�^6:����<��<C =��:�`�=����	�<�w��<�=^��"�<�]ɼO�=K�
=j$$=���<�!D�A�2<U�Ի:��F0�<C��Z@<���<��><׋��զ<��1==�q=�����Y=����<Q��<+D��O���#&=b���=��C<{j	�M�7�B�����;��=��t�7�==��O=n�<l&r�U1=��<��>��J�;�o�<`����2M�#�j�:��q�q�<3%<�5��L_<�x=�^=�.B<q-s<��y�.-��<�$;����:���װ���A=GG=%���=�v�:��Q��v<Ԅ�.�:�6^�<�D=�+=MY�<�< 	༵=&Y��߼8��<+=e���1=�Q=W�e��pS��;;<?�wL<<*�.<|D��+Y=�� =��g��/;9]=�p <f�C��"=_�<˦k<�����WC=~`�,�D���!=H�n��CN�?0�;Y���q4<��1�2Y=&�Y����t�U��(�<��;P{�=+��R�=Yӷ�"��<gP*<�P6=V;�C���'=�;�<�j=�
�g�=+Y��O\v��OG=�W1=]��;�n0���Q���漊5J=9:=0e�<�.'���<��;�MqP=D�;#,�:�Ed=�B=V"��R�ݼA��<�n=dx��[�������<�<��=G�;�ۼsR��pC<��<���<�����A�Z4U��ﻼX ���R�<|J��E��Ɉl=S=�L6<7�w=G���DK�E4=��<5�r�`�-=�U=F����Ѽ�;=��&��%;C�<�i���CO��C�0�[=���u��X=7�k�hz���B��ڍ�eÒ;�8�Y�U����T�=g�8�;i��!�*J�V�<��!=2�|<���=��e=TgO=EE:�X'=%i�7��<E =
���CF=/k]=~�s��6�Tt�<�-=�̙<f�� ���W����<��h�"�}����<�ѻ�63<h� =N=E5E�Ύ��Jɼ��=J�3��{��8�<�U<����x#ؼ�΄=��<�{�<�6&=l�Y;��A�3؉;m��X���5 ���X=t������<�?��lڼ'��<�ˉ��B=�����=?�K=�6����=T�<�Wt;����v<=��<!H=ܪ׼�>��h��9���؍�0'w=n=�P=��,=A��<ɷ�ݴ�<�m�U�k=��4�e-�<�b=Ϯ(=����d�:
?��m
�ῌ�P>\<V(�18�����]��<K��~H��^�T�
�8��=�:2=�i=�1���%�h#Ｉ��;'�;<2ǻ-+n�o<�<sI�<�h��*r�;�3�7��<3K<���{Y	=��;U��R������Q<?@=x((�� ��~=%���`�܉�:��<(��a_a���6=���<Y�y<�D=�.���i�%��E� =I��\��/�D�xG�< ���`~x=�0:�U�e�@����|u=�]=�C=�h!���G<K��d�h<w��հ&=�A���6�az=~�S=Q0�:��R=�!=EB���0>=�*N=FFE�a�T=�u>=�R=G����T�Z��;DA<��=��x�wD�;�=û�� <��R��#��rp����<H
�=lfP:$h=��O=�*�~�|�<�{< �K=V�S���!��<=��S��2����1�<4�;=��O=I��<��<n���`��8D�<�wj�L[�.TU��5=9ʹ���q<}� <0v ��g¼�i�A��;joe���ǼYZ�<eP=kLK=���;Q�����<�b��I!��&%q���v;d=T����<f�g�/ �<}��W=V"���O��f=&�N�S;6ݼ�����,C=�p=�تO=h�I=�-Y��솽=Yn��� ��"�f+�<�E'=�|<������W<Zg��_ȼ�
/=���r����c�c
�;UG���޼��:!��;�(y<�5=ޠ�;��Q��&H<P4�<���kk�d ��K���o��!�m� �m8k=8>�ߺ�<���։=��)�n��<��F<6��:�����F=�Z�C�u�Tf���<4�_����<㖂��%\=.]���<�O��ۉ���6�<����XZ����y<y�[h+=��=�ez�H	*�F���G=�h;���<�#h�>��:�֊<���<&i[=��=S+�<s	�<�k���g����=��M=I�{��=<[mp���9�Mz�,�A�2�<�<A�<�Y7��f��	��c����F=����ɫ<	켭��<_�6���<.>=ex����<�ƅ<�9�=�
=T�0=��
=VS��<�7��K��/,�=�3=�ټ���{̻<�'m=W5< jȼX^>�L��<t>�VV;o�<&����ԝ;�TǼ֍�*=�~_=�<��Q�!���0=���n�!<�eB���;��<��g*P���;�!=|+=�.'���<>� =�lM���d=��e��!z�?J/��/߼���=Jo[�f@T���?=攼xs=�n=$����9��a�=T#��c=i�}=P�="R��FI���*]=`J�=^�A�3<:YG=�=�v�N<�Z=T���l��T��i�K�<�$�=��;��N=Bc�<���<�Bs����<��h=K�<��B�S4=��%��=�<�����g=&��<1��<��$��gA����[+Y=�z���y0��,j�6ں��!�����}!~=-}�<�F��s�߾�;�\K={A��=-=<�*<6ȓ���.=��+<ff"=��T�g�<0�����E��U��0��d�h�H�.�<��e��<��<��D<+l,��
���@�F�E�2<-r���b��ZoV=1�5���o<���<�4C�z<�7�m�,=^�_���<zwf�'Z= qJ�q�\���B<3vS��`=B_6�r<y�	=�k=l�/���F��w��_s�����`�<}3ݼt4=�ѻ>=��<��/�G_P�&<�����:<{;,���F���¼�a���e�4�Y��C?<%1���=��Y�^\P�ޒ:=�q��eY=�����&���=���;��𼑪[=���6=���<��=��=��8=�놼%ϡ����<�)��2��<]�J=��<�@2��Y��V�G��<�n=9q<��g=� �E��<������Hl9=�?ֺ���;�{��"�#P=����M�-�<��:=<Bh��L~�7~�:�=<4M=����ͰW<���<ʟ*��1��0H����;f�ϼB��ң���|�Y�����:�M�g4'�����}M�M����;�-�4��;t�,<I�7=ޙ���><��#<��E=Z�\=Oee=g|V�x+;�$��%��$�6�j<H=׼T�y=�eO=r����y����f��T�;L�F=��鼿lS���a��t<�_� �<^G=L^;�)=`����)!��M����<��׻�!<��8=t�O=��< �	=�8=�޼�p�:������;4{t����<�6載�3=�G�J�<P��<`?��%���4l�T"ּ'B6�$�i�U�»�>8=܁�1^���@��R�<���<	���"1.��N"<>���=�R(<M��<�Ͱ�/5=*�}��<a�<�缇y��S��DX=���K1<s6o��6�vD�f��<Y�g<�SO���%=rh�<�$ּ����bh�3=ZQ�϶M�ƞ�<ѡ�:K���J%��H�s�
Z�+f=Ǵt=i�!<�qN��*��
=Z�T=.�=����3����L=���$�<��<=B�߼�Y�m�4���޼';;��0���ۻ|�'=����<Ǯ8��߻�PP�x�K=Ψ�<�@V;jC�=�p�<	-	=�w���&=0e=}G>=_��<w�����}<Pi�x�Y����<U� �FU�Y��;��A<��;�>��^L��'=Y��;��Լ�ZD=n6c�N�<t��S����4<5��<�M���<�1C=�p0�sh��N#����TC<m`�=�뢼�+<AG:<�]к�<�{>=���"7�<�	)<�E�m)*�U2=�=>�<H�A=�4W������=U��<��W=�e[�!�d<�[��=��<�%V�_
����<�z�� ��B"=����@�
�~��Q�=ğI��+p=�):�;�<��6g;��6���sV�<=��<aZ��b$=�.�9�	�E�?�@���.�%~=8�=:�h�U��<�o=Vn����켏�'=�[�6^W�!(��X�^=Bf`=�����y�0�=�J=��Q=Zy_��[ѼK]��;/��F;d�C�cd��=з<���<0E�'8l=dWD=��!�W촻��L=�4<�C�<d�-�
�b�� ʺʙ<�� =�sa=��<�%k=�!q<����
=#5{�J�<�#j=�8��#��d=pIR=��X�)�e=�֙;j�<��F=�C�ͺ(=�e<q�F���<)f��.���m�	<\T�� �ɼ�2�<Z��<�m��u��<��Ҽ�M��ǻ�`�"��3���ve�!�`=��a=h�<iƂ�n��ʔ�<҃޼��=N.м��o��Q�����Y(=#�S��c`�Fc�<c��,�<K���S�O;肌�g喼+�j�9i��8\�iE3��I;y$A=#	�<#r�M�k;�V2=�:���a���J��J׻8�D�==Y'���1<ж���i<~̈<��T�ĺ8<lxE��7�\i]=��<�i<m������mx<#U���<�:�'oF��{h<�-=� \��,�<Dl��)>�K�a<]��?;�sN�ɶa����<�:7=�+n��V�:��<�e7;QG�:� x9?!�;�V� �#'=��m���<�Ɣ��PO�LD7���m=F�A�<{\+��<]���R= ��<*�<���<X�=�FA���b��k��݌}�F�=���M�=d3$��&��el��wn���C�AD�qr����a��O=��C���=�˼Li�Y%������i=F��<��S�^+� =V7=2x2��h�<��|�=���c�9=@�g;��
=��<�����<�h�e{s<�~r���=g�2j�<�w��m��=����< F�m=+�<D�;e�:�#�<�=�o�s�S���Ҽ5�;=K�=NQ����<�z'=X��:��y<�������<��=k
;�X=�=ؖ< ���qr�9N-3;7�ü%Eڼ$��;%8������%�:G���ә<���K�)���m=%�����/�u�l<��r=�;�<>��-9<N�I�Q#�<���2�o��;p�K=��<��,=�I\<G�k�m���H=yPڼNV$��}=ep����"=����<ek������Ư<�*�<��<߰�:�b7=�Uu��� ��]�<}�
=/$(�N�=k������<�y<N��)�(=���<�(=����<y�ü�[-=��o^={&=��=��6<~��?F^<�W<G��;1�<5�;=�/�ڬ���7��(ʼŭ�<�|8� �K����;� T��L)�O{���;j(T�[�<Nt�����;^ j��=y��<��LK������X���,�69�-:v7W�vd��<(l9�2}���O���==Y���!���)=�p��� =��+�î�9�O<iB���|�<��5=yA=�v�<�:л��He��kWy�#�<=c���>�=� ;=i=/���$/ <f��*Gh�����dH���C��������1=5md�qp�;6�~��0�=DH����<�u=0ib<ҷ�<�!=yq6=r���g����)q���ͼ�����M.�n��;�g{� ��=�N�<�����G���u<K�j;�k�<?o=��M�����+�<K����Rt�@��)�E�Ֆ=x�?=�.��v�~;���=�v�1�o<cLS=ik�<��<�a���=��}�@�o��fǼ��h<[o]�AM,=�?ɻPP���;���?=���<�U<�%M;�h�1�;)5�9Թ<�O�,�[���i2���=�H<�H�K���v�2<JƊ:�
ƼX%��ٮ�<�Q���Y���n =خ<��ޑ��� �K��t5�<A8�<��e<�2�<.!8<��<������;?��L����~;#k� �<u����x<:[#����?�M���RhA��^�Ӫ�<"��:ڤ��=L<��Y<��/=K�M����$��<�d�	����2�:~ <�0� ��/���v=�N<�
=�=	)�;7v��t��s����_=�;=\��<�,=E'�t5�e�9I	=h =|�Ӽ�p���D����E����3�[�4��ȩ�x�n=˨|<��<;P�<�=ǊL�qL»1��<��k<a1�<^Z$=��=*^=��<�$���/��8XM=�*�;�׏���=iö�`�;�I<=�<%![��E�< .8<7-=���<�{�q?�<s�x��IC��IF�nqJ����<rU=�6#<�U�6��;c�ܼ��<M�<Q�(=�U�=�K��Y����<tb��k�<ī�;�^F���
<2��<r�Uk���D[�;蟼k�	����<���a�����`o��X�R=P��<FE׼��<�E׺^�P����$��<� �<r�r=�"i<K&����;���=a,3=G�㼘���$��f���-��7�<g�w=��<��<iR�;�U<�!N;��<��L<��-=��<i:���	=�8��m�<U&&����i�~9E����W^�<s2P=����(�c�t�@��x=9n�<^�P��I�E� �8q޼�_Q=؞"����<�㼧�\=ae���W=��<�KW�E%=�<�$A�5������)�<=](<��=YU�<Gӎ����tLa�1�=yT�<��<������=�&�:4�)�;W�����}g�<L]�;d0D�3a=���<�C)�\��2NW�����C*��x�;�'=_���U��R�<���<��=�	=:����i�����
=z�=��
μהs���}=�3;Y��k�<�g<\r��v�:=�ܼ<�\�<F]'=�+G:Z�E=�b=���G��;����6�;�s3=9��<|�}=g�<��<K�����<ME=�vU�'��;z�m=�k��ݼ�)���O=�6��@�<�3����n�;�n��v�X=�<a�Դ@�x�<͟�u6��B;[`=�Ge=��_=�:��p=)�e=�,��-�����bM=��&�ſ&���1�)ʼ+2=���XH<�(3���=s-d<A�u=��;a�=]tU=Ds���/�s��;M`~�3�;��߼
e7�S������<b�-�@r��R�R=�(r��1�<04�����=�ջO�C�w�S����<0���*�<p�.=��[�_��&f=
x`=[����=�=ۢ��3=�W�Q����3E����<�@'=��<����F<��=�i�<]g���<�,�<��<��j��X�t�;��9���|��)�<�bS���`��p<��#Բ;(N�<�'<X��e��;rC�<���<��~=�
#<���<MG=��0�
(����Ě-��5�����aϙ;�]��p�E���>����<w;X���=�<�8�<�	o9��=u$�=X��2��<��R�R�=�O�A�p=F�[<���'�8��̈<&��;�0M�XmM;y-�<i,1�~����̼��;偩�+�0<U�M��R.����<���7ꍽ�Z�<�� ;�� =�Wf;KS=g���[�ʼy��<L�;�E=0��<�~�=�p=�f=8����<D@�<�P�O�}=�`��9V0�Z�<��ż�{0;�fC��2=�O��(9��w�7=�v���C<����<rz�*e��1j༎&=���;�i���1\��4;!�2=h�!=�\P���<�Z�;̕ݺm��9�G��p�B=~�2�׸���-=��-��S���򼈾��(�=.j��. ��E�<��"<s�~�!�D=-�̼K��m�4�[_�<�;
=6�;dVʼ2�����Ck��&�y<9uS�wG�;��N=ʩr�y�m��ּ U����<��=e�< �<�\S<�Ga���==[�+��x_�y�<�0�m���jm�-[���7��3�<�50�]=�w�<���f�<���;'=μ������q'Ѽid=�w�$��+�%�5�=�}��<���<�#=!&5=R8=�=;�C�;��p?��<V�@<��]=6��;��<u��$�;�-�#�K�t��<�^�Y�;��z�<p`�<�ܯ<�(W�i�o�=�Hm���+G=*�<wL=>�9=�Ӽ�����f��w�=Ӷ�=]�L=�K�=�HY=��x�r �C=VG�;���<F�=�`�<*�<bDȼ�D�<�$��6����7#�3�����Լ�'==��:�r�,��g���'���<rMɻ�M<�T�3=����U=Hq
����<���;�G=��=��;���<�b="�:Ljw�3�<$H:���<�=�P"=rk<�c�<)��;�k =�5��_�<zW�<멗���'�!�＜��<��w�/S=w(=�S�ҳ�7�2=iF��h�{l"�:&�=ߜ<��1���6=1�<��I�X=�Ʉ���B����L4��	+=���2 �W�;�z.�<�>�7淧�.9%=38s:�c��6�V�<w�$��R弛���i�y���-���W���&�� 
�M�]<��� t�;��&�-a�<&m�I�<Рۻ�H���6���z[=犉=��<�K=�m�жb�`6i�u��޸p���=++��@�J=��=�FJ=2t���	=��缼�!�v�O�����<�����HO<�A�D����^=�)Q<�02�	�V=�= C��(���U�g�f=Ҫ)=����~K=�<v�^��]=�0�Td+��~�����;�Q!����'�.=e��x=��μڼ_:2�Q<��<�`=B�,=| 1=�=�����V<L���8�� f�0��b���/=���;����b�ռ;Ɂ���=s�K�J6�;4r
�~x{��>T=vYL=���'�	�C̐���������@�<%1��ͬ<㈭<7�N;��D=k�X='x�<ވ�;��_�0D=�5�%�}�*����<��3�!.i�Z8!�<a<V�#���<A���o�=���<��(�������`=�ż�"=v�<�v�J��l<?4�<[F><x�u<� >=K�_<zӻ���<��˼�=�,M=%\ӻ�RѼ�m��?�.,T=q��R��<k�=�-+�_�<(JB<��%=�RJ����<�f'�Bο<�=N={1��5�'���9�:5��8�<<��<����9>�e�'�Np���4�9�<����t=.�d<A��<AE��7�;3=���ͱ:��s<�r8��J7<�l��Ȟ�۬9�`s�<
+r<s�g���E�P:�Zŧ���A=��ֻ�l7�U =ٸe=UiJ=*�*��J˼4!򻻌����7�=�Se�����<�}�<�'N��稼9s�<�={��Y�=t3�<�G�=��<�s�;ߥ���m���rT�y�	=`�X��!f���J<�k���k��5<�1T�R���=�`=��7�.�<��<3�O={X<���FOR=@�F�mJc���%=�B!�B�B=�Tݼ�Xy�)=䟄<�l���F=�#���+
=�����
�<m�,�1=>=7p<����,=z�^��K�b��g8i�4)!=02<�=�����R=��a=���X�u�=+z���N�W*	=�C�<�k;y��<Ν=t����NԻ�U��D���J=�z2��L�$�/�D':o�n�r���&v�%�o��9�M^�<�s�<����=�4���a�P�a=�[�8��L=�1�;��}��Ӭ<* T<�z��ѰT�뱋<Eλ@��<4���ؕ�-r@��k�<9�"�|�!�=���"؏���(=(����؞���LڼC�W=���B��;��5<"�'��Hż��<��
=ٍ�<��<�f�:�V�<�5=)��<�F@��<�<�(*��.���3H< [�;���K=���բD���M�r~^��介]=�Z=��<L>��w����̼G��<�ϝ���G<"�=�1��"Sй�/�ꡥ<�����=|^<s)�HY����;�0�, U���<1GB=�0D����<��U�:�;�|�Ȇ�:���<FX�Z�������<�;���<������*�a��p#6;�,��2��oQ<@�7��>z�Eh[=@������<}^{��i=_�"��u�<wc9�(�=�/V=���<���;��d=�<��<}$;AS><� ��E==�,���%=��3=�Ĵ���T��W�������"<�Y�˜�g`�u�=K,_��7<�5,���N���u��5�	=A�=�x='�ϼf6��0b�4L=-
�Pv�<����K=Z��;��=<&�'=M�U��3=����<|R?=�I�<w��<(�=Q�ļ|cg=D�OZ5=�� =h�%=�W��X[���w��#�2�S4�E���3��}F�A�0=�s#�^e�<�m�<�:�<$���	<��;��2w=�ϡ<���<**��Ha�<�X	�p2M�M7ּ��=��<�	<����0;�.��綿���<�=��#�<�C�xV������l=ب��	=��=��&;���#=w����WżT��CSr<��[=}��<�	�<; 965{��{=�nY�m'Q=�b����u=e����<��<q�/=�3=� =[(=�G,��b<<W�"=����#r=���� �=��K��=��F=�������13����< ���3JU�*\�<K�D�C"żq�m����<�bX<�+��U�'<E�;9u��8F�X���/v�6�<��
=�"@��{Ik��R_=�͸<R?=�۪� �0�R�J=��A=iE<pq�<�	�����ĩe<�{���	U=O�ʼ��P==�ʻFPb��|"�+d����J=Uwd�yz`�M�O���e:3k�;cS
=¬u��L�i��<i�<K��LO� żY><U�<]��}�����<�=S�]}?<"�Z=�m�.k���<E���K=Q���
x���	=�=1=�<?�l��zd=�b�<e�����=�v`�� <J�8=g�<�0�N�	��g<�Dc<��F�I}=�C���'v<��n<�R���&�:��=2�ot#���E=� �׳	=BUE��+/�X����!�9��<�ɳ������<UE=��׻�@=d��<۲k<Z��Z:�H�3<���<�H�wr�<�+���;E�<4�t��7μ�hp;'�4=��N�I�i<�(%������5�<�b�;a�=�.�<U�I=��=R�H<M���^�����<�=�h=t/�=.P=7�v=}�:�)�<}�<�ً�h_3=H������
�A<�@=ٯW<��9�;ȼ@�h�[����;��-�e�2���<�b=ڑ����%�u��a�=��A�>L��`�o��<?�\=���<)�мh[�<�M7��9:=k+=�5��!�ȼ�R��P*C=]k=d�m=/��<���T�H;��M����<�	���2f;$�&��Z=W���F<��d��?\�Ÿ=�@"����ۙ������=��)��T%��c=
����G&=-(���!���v=�5=Sؼ��=����6= �=Q_
=CjU����<�"��g�;<�ʝ;�=��T=�9 �T�m�������*=�&��=�!�<z]��)��-�B���?�<i;V
��}�;�`�y�̻RW�<�H����><�(�;��|=.�ϻ.iV��s�)P�;{��Q��=�;[s�!mY��}E<s�����%=�|�<T��<��+<=P4:�^��@@�E�"=�C=ƕۻ[K;��dļ��<xX0=�1�bz��Q�=>��<;&j=��<��	��v���t(=�Q��T�(=�-9��1S=�P=���)F2�����̫R<��<p�M�tt{�k|���.��+N�7�I��L��Ih��$Y��@p��D�8��<�'=h�O���<�����c�Z�<���<;</ <�
\=�MG=�W2=h$=WnV�l
�<#=��h=�|}=��ʼj��<"�����|<ر����=I���l;$��Ⱦ���5�</OO�9��<��=��r;�ܕ<��P��G<�,L<z^0<41��WP2�1�����<i+n=.�<߆�<^E=q=�|[�ώ���?ju=��Ի7g�<��f;�o6=�i�<;iD<��;�ۉ�����VQ�� ��g&<���;��a�˒���8=���<��G�J�<<;f��<X+��#�m=�x�<v�z����<l�<�O=�A���c==�;ʵ�<�0=� <JL��x�<Bp��8�m���0���M=v�W�fO���<��|������<�c=�8%="�;L8,�J4E;�t*����<l~�<+E�<-8�<�Oi<#Y�k�=L�H��ب;�(Y=�u�<� F=���؋�;�-=&�	=K�~�/��c=�l�;o�;���4M=�a��:����<H.�=T�=�a�<ؼ>h<�J=��J�|~�$�=Ax=J��;q$����=7�-=�hP=��>�c�׼p˼Z=}�=�д<��8���?=XT=8�� �<Ӯ?�f�1=�V=7���2=���B��O�U<U��{[=i�J��	D=�s}�y�����pU���l)=�S����@�Su�T�;lм��U=,u<�
��=v�>��D"=fՠ��8�y� ���$<Y�|G��{)�<�s�QW�<̽)�!���>h칟k�2�<�qX�8Б;���Cw?;��G=WV"=}uP=�}��^# ���J���H=�6�;��=4�k���m=oz��f.5=�W���X���Q��*�<x�|=�Q=�o���N�<���cV������~�W9;'����Q��S�Y0w=�@Ǽ��<A\X<�^�<��<��B�m!�<$�l��ȻD�59�=.�-= �<����E��.P={�X=&0G�2E<��}�<7U>�w�����=��<6�8=�Լ���<�/�_Vp=%)��
�-=Ɨ��D������,�0=�[����6=� ='�&����<x�;�l�<���)�;�#�=>�<�;��C���Iu�����������"=�E��㦼P�<�`[=k0���]G��=輇�ּ�,�:該��3]����	C-<5�<<�QF,��V�<�׺<X�=a�9��3������Լ�|=v�
�YK=�-��<�t/<WIN���=�	o�b�;c7=H��;TR�N��<w=-�?���!6 =�b<p���˾=b�м-'��L=�7��@�<�sS����<�T�,P=��*=)ԧ��(*:cn=7�<��@�Q��;�S����=��<,�>�Hd�<�$�<Z_�<%��<�W=��:Tʅ�&@y<'"� m=�R��8%6�b86=l�;([�4<=�6=�^����<?vB=�O!=�"�<\��<.���<�J��J����;u$���=�l���M=���f^A=�~y=W<�������a,=:y��=�
�<F�<��<J&:7��<�l�)\����!=�Վ�E��<��'�b#=���{�<��<c@N��m��*%9���L=m�M	�}�ȼ�\��Ta;����Z�=�	R��t�<�����"�;j0�9GC����T��k4<h��<;)����
2<F9=����F��RV���W��e=#��<E�Ǽac��C�4�t$�<�B�9w��<�ia<�	�hho=��9����5L���+=��=�_<� �<�	3=������B=�%�<�/�<-�ϼ�޲�8�C=��	�#���=%7�;����#�<�j=��S=e=rx <C=�.�a��7�<��.�fI=9��;�C��0�;,5�<kEռ��'=��R�!']��=B�ռ��9=�x��+�X��Y*=��'���=O��y=��f=ف�<w�L<wr=m��X�<�G!��(<o~k;�ٜ��B������-=l������,}߼�1�<v�#��?=�t��=?���=E=;dd�i�<�-�<�`�< ${����<9���_%=T
�<n�`=ɘ�<J=�H�<��=��K=J��_�����[<�T���;�Ǻ�.>��q0���T���\���<�4�=&Q=�6�<�B�J^[�e�L���B���<�1=�?b=��b<'�����<�&��������@_�<CZ�e[�I�����;�s�l�,�&+�<���</�<z�`=��%=�%����ؼ��ȼ���2P��x3�̼�$�	�>=��<h!E�*��'��<��O:��a=ÿT���/=A�5=X������<��;�\5�^��;_ =>t�-�<����X�I�=�S��s<��F��
=��<Ğ$�%�;=eKX��}/=� C<FX=�.=ea�<~+M��6`=�2i;�bJ�2*��-�O��8R��u<�<5c3=`=�<�%=!b�<a�ռ��N���ܻ��=�-G�fJS<t�;ş6=�&�}�=�l�<���;�y�������⣻�"|=�쮼 �M<�'*=���<��D<b�c=��;K6�Bm#��-ۻD�<d����L��'`	=X}=�MO�ķļ�1ڼ���:xX�����`���<O�!=�5�;�&�;�)�bg�ٰ<���Y�
:=�==�+*=�e�<�����\�<E����{&=o[=�O=>y˻ʑ=u듼攊<b��;갶;�D�<�A�?=7�V���`=�T����%=��ż�Ɠ��x=�����=؄Q�L��<+]=H�S���3<��=q�<m�M�6��()��!�����'=�)�<����r =�n�|D=
܌���q����:փм?�<��Z=uvV=1�L=�ꔼ1a��漢"̻]ᬼG�J��� <?�C���	=��F<�=(=��3��_���ک�M^P��6�<�Z���<� �;̮�<�Ne=$�"�!���Ɔ<��&=��x<1Q<q����Y#=�� =�9=eE�<�K<�dq���Y�8}�<#p<+��;�<4 �<��=�`�<�&�ٓ�<�����ͼ��Q=w�O=8�W8�<�l��:e=EI�;S��B�h��%���<�H�}�=�mI�Rռ�%�T*��B�3=?=�Y%=d6=��=m�(=*g�<d5�;��5=���;��C�U�ݼ��_"���I�����t�{;�x��,ϼ��B��Ĺ;�!�<ͤ<�,�����;�D=w�K�<+���g=��E=m�=���<�=�>��.��-O=�}�_M�
�����<��s�#�������5f=vg�T{$�~/<{����ۀ=#t�<�_@=)C�;[:�>�=��X����;rW=�P=�WH���<��: ����4=��6=ԯ,����;
���ɼ	����?)<Q:=��i��:�:9�[<6=�X��Ah��?���)�#6�;��<�qP�ε���,=e��<��D��Ѣ�0Ll<�b��.q��c&=�,�pU=Lź�����i/�^am<w�=$l$�M����`ȼ���4�����=V�*=��_=>je�3ٲ<��u<�w���6=yMƼ+$6�ޑ����J6g�S=�kӼ���9aV�;�t=XA�l�W<SF= &<�i=�P[��%��J%3�m�S=�<U-�<��=�l:����<O�<������>�?MI=s�=/�"��3��� �:�3<�$��>v�I�=�|��BJ�pͼ��$=�#=��r�9�]V�]z������<��=��D=�zO=��M���:��5���D�zF|=t�ջ��#[�=��(<ُ�;��W<aD�<���=�cx�5''�dZ
��m<�3�<-��;��`=�'Q���1����*d"�d@[=؍=r0<e�<��:��p=eY��'=�����������2t��sV�c���cA^�;fV�p��=�W =�#�<t[=���<�4� ��<�o��-yN���;GT=��i��ʼ�>S���c�І���&�;:=�E��A�<%���UU;��q=�F�ٛx��>=/v�;���<]lR��{N�c��oFS�/N�_�X=|�o<\�M=աP=��
��;�Ꮌi$n�c���|�#=5���f���{���D<�p�
�=\!Q<���y4�<F�<��I<�3C=u,�̡r��)���;ppB�2�<	\r=��n=ݫ-����=�<[��%AS=p�Z��ļLj�<"Rj�R<���ͼ�>�6��752=�[=�Q�<�l0�nkr<�����Y0=�H<gI�<�	��ad6=R���ۼ&W�� =�|U<��N��<�L?�,1��l��[�<ǦX�����~G��iǢ��x\���^��=�<�[��pJ�<8Ho<Br���Z������<x���R׻���6Y=N�Q���<_�D<o-�|��-!��ې<��H=�:��+��u��XS+��`��<i��<�4=Ɉ��&)�b����=�a?=�ޭ<�bn<�ȼw�<��<cX)�g;���a�����<�%=����8=�x����O�Β����� �;�@�rTV<Nɮ�Y�a�ɲO��^j<҂�*s��?�<k�<¹�<l��G��<�b�<Avr=��=Z	 =��4���`��<l�g<1���a�L��ciu�P���E��<gɔ;��3� �&��L<<���s=�S'�c����<������<�kh=�~R����7=�\�8(�v;�G���;	��;4;�����f������� =p_=�L���4�Ļ?��AӼl�;i�<�= �[�{�=W�����5��<�݁���l�4�U�Լ�<M�i<z?�lD=*V=��==P� <
0���(=��+=+�<>�d=��^��Y�<]��<Z���Ї�=Fb��9���B<q�����~�(��<.�0=�wm<�=��!=�*=2�I=F��<yc\��C=0��Ѱ=��=�ּ���<�O�ϑ=�['< ��<�%D=��D=�o�;��	=�4��[_��c輭��P}|=�8<[4�_�м��;D��<��G�=�N=��`���?<{�_=��D�`���0L=�+@�\�C;FI!<��<�fT�`�8�Y%x;���<�28=��;�Y����.�<���<��A<�9�Q~�;>�-��1k=|s�<
��=�f2=���<�Ѽ��ںɠp�Y�<_�Q�N#�y8�<�K�j5V=�oF9�x�<�Dɼ��<%�:=�]2��;���;m=?=�xw�	�C=����}����
;�gZ�:b�;�@�S��;~=Z	�9�]�I@��6zk�g��;}�����<L��<;u�=�UM=�@�<!�U��;=�Qp��=��<��	�<�G=Z�<`��ZP=��<�L��0��wX��ڹ��D$W�M\�����<��R��������<����w��m�*�(o=�;��Q�T�.�=�wH=pO"����9A��=/7H<��#�r4�<�ԩ<PX6=W_������<��:�'"K��'����=+�A=%�]�L�&��>�>O;mȃ;��K=�yU=7�k<�ei�-��=!�4=�4�<z ���;1�#�-�m�cy����� C����l=��P=�\-=����3��� <�*=����c=��:����-;<�C�<��!����<���<�;3=����=y�޻�_<�_}=7#޼+��<�`9���0���L�񞻼;�伆������9��<�ʂ<�E�<��=���3�\�J�=.va�ɞ�<���9?Mh�&�<�)��Vy�A1Z�V��{߼���8Z<7�
=�0��_�q��yF=l�<��"<<�;�
=`\�<?E����;� 4<�m׼�=}�;>��=X��<�}�<aI����P=��V�j0G�d���Fz=��E�uf��Ѕs�B{�cU�W�8;���<����eoV=vi =$s�W��<@!�r&p���<�aD�ӱZ<�PP�`�;��K=��M=r,��`w�<�Q7�8�� q-��ڻ�a��<�6=��ܻJ�e=�H�����w�<�B=ĢN='�N=֪�_�)��=u����	m=|�"=^�o��>=�Ӑ��M�����<�?���<�$=�_?��P<nL�A��<4)<���<u�	=�f�<��8�щ=/V�<��>�J�U=��,=S�F=��;��:�xu��W�<�\|��W3<���].=��D�j"=�S<l�;!1+=�N��>]<nZ�=C(�<;�ļ���;�a�<�IM���D<�=G<�5�v6�<J�<�a���a�<�H�ܿԼ8�<�<�6C=n�=�m�;���<�X��f��������<z?����={�μ�۫:X]�:���<�Cn���r<!X$��&;c�<�:<>f=�y��%��<f	`��fV�⮼�5B=g b<	�4�Za<�4g�<~�b���.�d�)�zE�:��<�%���:=�.�T�P<R�
<��<��:=\y@=r*Y��	<\Z�<�..=h�%�;H0�f.��K�3	W�Q��<�&;�0=�=�(��<�^N��|�-�,=�!Y=�<`�o=��#�#xԼ�	<h(H<]l��%=Y�(�{iɼ)m��HF�<�w<�z=n�?��=��޼�Ͳ��ͤ<j�<-�<��'=��<,a�&<�<����	�6���ջI= <���������u�1���=s�=�,<=;O�f=�<�=v(=���a�j��.�<���n�N=�hg�׌Ӽ@I��G��<:؅��i-��
[��J������A���YU=��<��!��������-=H�E�8CP<Q�,�켮�;��<�^v��Լ�a�<V�K<zc���Y=4,�<��g���<3���ȼ[ ¼�ﻱ�<�:=F�E= �=�ጃ<�Q`�/���U�<r}Y=�3=�y�,��}E5=��&���(=n'� ����8�ı<���?o��_���S��2��=\A=�$=l��<�e=/J��Լ����Լ���8dK�,��=��#;t<�;̙h=GK=�,�9�,=�D��e�< f=�6�	ٳ���`=a���=Ux�<��=rVG=ɼ׻a�f<�����<�b`���ڼ�Z��%x=�;�,X=�^�<�:�4�<*�ȼo�
�7<�<���;>��<H%t��;L�T��<������ۼ��8=�=�x*��4z��Q��{i�<*��<UܼL�=u�<x �<��\<�{C�P"�/�W<l����y��H��(���5�;��M=�=���<^�L����;�+=e��)]���:�����2����< 	g�?�>�!=[�����e=ϰ�A�o<��h===��%�=j��:@~�<��<�M�OO�;�7���ۻ��*��4�r`f<���C��sut=^f��ݻ�����9�y��<�!"=c!��}
=�'<��2��HF=�[=#��<*&!=��6���s�ӛM=�b�g)P:�8�=��);��E���<~��88c=�=�^\<Ϥ�<M׻��O��ő�G!<�M����;��<F�J�C��;ŦY�F������*�<��B�>����u6=�_���=f>�j�<s�+=$?B�;�C=[�\=�N�< �==���<���;��<�ڕ����=��M�"��<��:<�K��<6j�1��;I����=l8=��b=Gb=��\�Ԭ���7�;�����{��$�<�U*��|�R�ټ:4�<�)V=3�<G<�<#_�<�o�=+�`=���ͨP=E���.g+��Ǐ�L=���L��9e�S�u��<��.=&��<6�N��2l�K���e�=�
輬s���Bt���<
<&�<���;�m���=�%="��:P�;�M��L7<� (=�]�jZm��ؐ<Y]�;�D2=��e�,�D�)��G�<ܻB�ڪS=M��<�~��叼acg=E�չ�����n<�8�)�<u��D)�<$��<^~c��b��A���-�|]��H�)��+=�9h�շ:=���9��V�<?��<F�
�OY��bF=�i;=�lT�+��G�<�߻ �f����0 (����S�q=�^<5�=�$=Ѕ��V-9�N2�
F=��7�6�
��)=H=��	=��<8�4=��;��
=&ӻthA�H�V��=Wd⻛��;�j<K��:x�=o�=��;��<2K;�-;�Yk�
s!<#��<Q�L:��޼�Tg=�>t�㶓<��k�][V=��׼�sλ�X]<��F�"��S<��<$<M
t=�W=��)���-��T��� �qz����޼�(�j-s=��/�ir4���
=�*?=�cA�$�J��=�0�;�m�i��<�5����N�}I=���<��=�lx=�(�;�]��9�;.���T =��>=�W�P��<�`�<�rw=^N��a2U��R�<�D���U<әz<�Eu�^��<��<����`��%,�����7JƼ'#�����8(�ӷ�;����!5��6j�`rR�x�t<<2=y����f+���<r�<,3��f�<�H��6h<��E�����P<[=�HD=.$v<�p%����<�̳<+�=��5<4�#�cI��6�<S��= ���_;���(��G�=*�1�Is�<��Ѽ��-,��h=4�?=\F��]�4����=���<W�p��X<=�<��='.)�dK��ߎL=$9)=,4�fo%=�D�oig=X_�<�>g<n6$�$'4��2x��{���v�gհ�\!�</�<DƟ��Y8�*>=�*f=��Ǽ��<���α��D=������.�(�<
��;-.��۾��=�<���I�'�B#=�$��>"�׽=a�
���N�)�'��w-�R�{�J�Z=G�D<E��#N6��1'<H�n������`�x6k<��a=�w��`A=��<F�3��S\�������<�����l��?¼��
;qX��q�<�V��c��=��-=f�ؼB��i5�����<�}�;��=<"=����꼠|�W���p`�aE�<�_=���<K�-��,L=�:�m`�<�P���&����<B�l=l9�<���ר`���=�Q�(�<�y���H�0=��；8׼(�ռ�Zx���T=V95�a(��=�^=dv?<.;=5s�9o<�֭;w��<S�=�I��6�#=���;��ؼ������|�~'U=@��R�H�e�}=T]�<�oɼ#�V=��a�lWR�wۅ=�]�O�3�K����<�O?=I�F=��1=y�=[z�}�$�Ҽȕ�<N�B=Xۊ;A�ۼ��euC���=d�=�b=�<�k�Σټ�!<Ā�<�{!=��&�iO.<"�=w�<��a�&�=T��Ӌ������m�<l��<���<X��<}�
�*g��~�@<=������<mYл&<��;��t<eͤ<5rI=��q�=70<���$v9=��k=���;"$`=݈�!���9CD= =�<Oׄ�Ԧ�Ynw�rI���h:=�̻<6�7<ʼ=�Q<t�K=;��!أ��᛼��.��i�����k�h���9gH�;��$<����aq=T�)����ϓ\==��|�S�$* =*�*=�Xt;�|=�3!�^^��q=��; ��ye��Ƴ<'�������'�=����\'�u�	������#�>W��P�$i=��=�>���o:�R����;C�R����<�����T���<��<�*��ُ7=ݼ5����<��Q<ɀ�p�F<Y�<��{=}_��i+s=�/ؼ,O�<n�:ms~����
�O��Qb=y8�<$���"��7��L~�R屼� =�D������8�`�1!�<��@�dX��Dcz=��=�=�p!�~Hλ��=|7�eQ���x�&�伳�5�N��<[g��}=�ތ=׼s;_tۺ��c�(�Ӻ�F=H��"H&<З��P;=~Vؼ��廝U�<��[��<��g���0���R=P������:����7A�<L尼;	���q�<��0= �Ǘ<�ټ�S�Y���2�Ml�;�C����=ϲƼ���f2=I =(��<U'^<<J��TӼ|r=�4!=��<ex<(I�����3'='�<������<��A���W=�L�<+\�;aB��/T=kL=�G<P�*��< �a��r�o�<>/I=*�9���7=z��;�۫<}±�k�.<��ȼ��;9�<�#���ݼλ��P<͊`�f�=�3��t��]�S=�*$����T<�]!=A�=��=�R�2=]��C�������˷����<J�%;�Y��q =�s.������˛<��)= ���gȹ�T�m��7^=R�
�67�g6�<����D=��B=]�J�۾�<�OI<�*�<�,;� W<�QD�a�=��?=d�/��F=��e<�@���ej=؋��-=��|;��;��.�FS#��t2�� �<�3t���,;�;���ݻ�yz;p���>V��BR=018=k��<c\�=��b<��׼�	#���ٻ�u����<����j=OL�󄹻-p�Ҭ��0�N� =���"���K<=���[)=��W���$=� ������f�vH=�v�~�=͎i=�b��p�@�)�5<��S=�BT<sXU=p�[�i.�5��"����Uj=ǆ��|~�<w@�<T'X<%���#*=��s=�1)�0�)�E$)�R�E���ݻ�^=�/,�q�(��cۆ;�^�x�'�f�X=�IC=�����<�+ �E�
=��@=G=��[��S%�^,k����C�_��������n��B3=��P�����2�u=_g�;�}�<"[�<v�<��
��u<�7�<HO#<SZ�<~�!=�K=��T��)����;�u)�=.��=a,J<@ɻ<��;��.=��2���;�i���~h���R	�8 �;��e�<=�쑼�R�<δ����=���=��=�L#���
=�3��a{�<�x�6!,=9���F|�</�=����Ճ;!�.�� f�j��<x�=]6f�~������<#V����;=ɢ=��|<��)=E��<�����>=힦�ih	��hڼf%�;�L�SM�_Տ�*��<��!�wQ��U�	��<�)X�uR�<��<ʷ���.q��k4=��]=ì�:�-<�����6���/=l��<��(=fK=��u;��4���2=��
=hOR�8O�<���V�=����������4=�f<*����{=���<������-<���<��ּ@��0�/��C������V����<��F=��=��B���F��D�<�&<���<[D�<%g/=��Ҽ׃�W��#=����zԼu��<�� =V(�<<:�=������dN��Pl�`ȍ�?�5���<ѩ���<�:�:)�*;�SL�¿Z<*�5=�]�<�v�PQ���ϼ.�1IC�n_e=��K���]=��P�M�M��*=�B�/� �=/����G�<Z�<3G优_�<O�D=�B=��7=����,=�������1����j�m9O��弾����7<ғ�;�(�����s��<i�a���M��� �b^=߹/=z�i=qw�<�υ��'�<��N����R���B�ű�"H�<��Z�7�x�\���:��W=0g=��{=��3��<�U=[�Z�\F��s囻|n�<���;%Ą<�'�$�}�P4����<����͸�D5=pe[;�9��p9?=���<A�Q=�Է����<�μ�t=x9�<��)=N	]=󲃼N�<t���V=K�f=>+=��"�$m<>E��:�;�[�<X�X=+c�<��l���[<�����X3=�W=̖����><c�\=����(=_�＠m�X�<?==�T����<�����RؼV�=y�¼�˃�D�V=�"=��v<д��B���޼?���"<ꀲ��3g����<~�*=R�¼Yg��;�=����26��<�P�<݁	=7�[=��C=n����K�1�:�A�<&`H=��\=1���6=V8=��c�/�$=�	�,���l;a����<2��(9<�}F=��(=�P�(���<��˼���YӢ<��-�̨���!=��=�lq=���<�O<`�-=�W{<�֕�5�=�����.=h�v<�j	<W�M��lw��>�w�=K7�<�v�U�<3�J=�>��e�[��]��y٥��Q�<=~��=ٺ�*R��bt�-��tF|;L�<��bC�<;�0=Y��n��<룻�U�v�ǻ�;<�<L��<g�J=��C����pi?���
=+��<Af!<%�
=�(;��м⥈;�=S==G=e��<A�e��bD=8�C=�T��\<��^�����j��c���[K��%��F���Х ��,@<m=��:�)D�;6&	���5=F⃼xӹ;�=<�;;<8�E=�ُ;V!=b*T�?TL�4�м$��;{�����߄h�i��qeY=m	Y�(�ۼ+�q=�z�/�B	S=)�<2=8�@=�?�<�<�lz��V��UMC=��S=�����X=s�H;;���jd�%�h;�M�3Kz<�Q�<��c�7;.��<��=
� �����L�;���<I��<��<��a=}�
����;}�;�ԼV��<1)������&�b���3���6=I:b=%Uu=�ZQ�p��;u�7��gX=�Xm��T�;c�<�Ҭ�~!�<��0<D�W=��W���Z�`�=���j<
.5=3Q:���-�<"[��<{!$=0B�:�/;W
=[�=��?�����Z=:�)��� ���c=EGU=���I�c=^�s�Z����Ҽ/C����������=Q<�E3�Yzd=݆�O@�;���i��*�<�2<L�<Ô��RP=���;�(�;Q�&�����%P"=c�H�v�T=#K�=�d���8�7�[�Ǯ{�DE9=�Ps;��W=�P�<<5=d�<2�%<�t��O|=][��x���3(������1���|<���֠����i��%��U���C���(=��R=F�}���0<�j=\�6�W/��O<D'���<:=�z ;"e�
�>=���� ��x�ϺӾ �,̕<���YY=��f��W����M�A��@�ak�<*ƾ�>���<=�0-=] w=z�'�<�:��= ���b�!����&=Ĉ�:� �<�K�;��<q��<.�[���;Í}<��<�r��FT5=����F�jbW= sD�a��<K�B�~�V<��*=�^=/�μ��#���;J�<���<.�<#q���yq=῾����<:�żWY]�9R_;>��i����!�#9;�a=nc= ~?<�a:� VF�ؘ<�k=A��;ޜ=�H�S�x�7�v<�#.��7<��<t�-=n}=�"<D�X��E��蘼	�Q<r]	=oo[�{�l=���;�.��;����<8�<sGW�c)�G`���=��μ�g��(����MR<Q��*��  ��^��%��ˊ=ѧN����:�g<�}'<�8�;6�[<(o&�H����2�<��=R����0<�N仿���M� ��M�ۼ�
��>�<���=e�V�A=�ќ<L��-s<�Y��C��
�*�v�-��#�<��N�t��<�T��p=hh3=���;1!=E�-=�mb;���G�;r53�z����;{2`=PF!=L���dT��_���51=9=�6�X����ߞ<����W�/=*��W�]�<�==m�;��3=�yz:s\b���<04=u)=Hȼ��;e]_<= ��s�C<��<��=�sB����:/����:�Z����(��j =��=�
c=�W��;{�=g��$ƺ��[��9e�`j�� ��<
�:�/��6�&�Z�@��\��
K�dM?���� <j��;���L<�V��R^��A8��u��$ =���;D&=�f6;L��I=�!=ĺ���<���<�Fn=�S�<E=�=R=+�E�7�N�=(�=7�E�"��<��#=��f�<I�nv�kƋ<��r=���<�Rf�B�ܼ�fw��7=<�9�;������^���<=��<��?�	�st<L�A�W	�A=*=�w�;{˟�Ĝ";����&a;��/��2�����g�Ÿ�<�s�.��<�bt=���<��Q�<���Z�W=Ĉ�Bh����<�bL��V޼(�P=������̼�m=�
<��!=����7G�����^���߼fN�DT��ǫI=��m=�Y���<��<��=�p߼�|�S��<T=v��<��m�f/d<*�˼5�<�:ü g=��t�G�=y=��2<�g=�qU=��C�ˈ�<e�ۼ�3�<>w��� �[x���0�<'�o<"�Ļ_&<l�O=���<HL;v?���!=XS���<'#_�>f=�*n�O:=�i�@|ۻ�M=tռ������=���:�.��16�E�<�3�H��匼*D�;�_�[�h����g/��3H=	�*=z#==z(�����uK���R=�Q�;F���C/=��a<��2<rJ�:���;gM�;���|�<�����)=�"�;�G��D��0�O��r�N�<�E=H��<L�V<H���gp��8���k8#=!���^��l0=��w<c�G=rx��=����=��NA^=�N�=�B�<N������<�
x�Ɯ�<$p�<!�P=��<��2<���2G켳���=1��5���"#=#��<�m�<��/<u�0=c
=�����1����$[={d=M&p��1=�C�M�
;��.=�����K=5#w<�n<�P=��G=D�f=/���Y�$��}��͍�<��*=?���J����2��>+�5׼�	=I�<t>=��:=��O<�����?<�q;���㲖<⸒�X�=���q�x�J=�M�<�Jc=*P޼�S˼y�<��f� ����@��w@����<=?=�u<��<�f�Y=��@����<v�6��V;弿d0�_絼"S=����b*B��he�Z�=Uuq�M��<�W��߰G�uł�f��^�j=�;l<�s�<�š<����E��;b�=nh<xC<�Y�O�<���R��<o�,=D�c;��e�B�c��S=蝇<z�8�.X���ݼ�I�<�Iy�S3&=m]E<��1=ca=���p@�վZ<^����ﭼ?z7��B=��B=I=u�Q<�F�<Ol4<��:���J(�<���;Kk=�;����q� =;[�<Q��S*9��S������u��H�@���o0ʹ�a;�e<в%��,;W�Ի��?���<]o����v��C��W<I��w	��
S=���,�o=:>n=��l��ۉ;N0<o|E��q��I���!=)�n�<����<ư;֯h�Dץ;Γ��L�.=�+��X��k´<
���6��<�e����;�9<�3=�7�< '�<��!���l�r��>7<����%�+=df� +=x�g��=�<�=�>�n0����::�:�Oļ�v�*�A��Qj<���<��=P��,�ɼ%=�핻0����oӼ�7=��]=x���4?=�8
<	��<�
R<�u���+����=�=V�H=q��<�?2���J�Ϸ�<iA��	!��	m�ݳ2�p�;�0`=��]��<E�J�2�=W�j=m[=h0=4|��c�˼�K��g�<����)��;�W=͡�yR^=�������<�q���=�&r���=m���?���[�d���<l�0�E,\=�>�<醗������8�P" ��,y�~Vf�1y��צ�<!�<b25��,кA�:e!�ƙ<+��	�;�8�]h=<��<��1=�~� 	�;ʠ<�n�;�=�<<�+¼=�<�Ɍ=.?�;M;=���<v<�L3=�&�<��-=�ڻ�B=��z<�B=�M�֡I=mR`��VN��LC=�8�<�圼��<��0<?��M��u�<�ġ�ح����2�x�L��#=���Q�=bJ��FO)=��������N6�3S����<�q)��;H���T[=�E=�==���;?d;�?�:�6T=e����̼�<�<脬<���>�"=��b��F�����UX»v_=%P=/�<G�=t�<ԈJ=�.D=����P���|=D���O?<ߏ��Z�<Sn;S�<HE�<�Ic�2�<���{/�;�:=/��<�[=��<p��������<=\�<��VA]���>�<`?��}#8����$=�#��|R=���x�7=�s*=�#����;���;s0=Gp �*�=��P<xh�<��=�E =%�1��G�Pr4=�����<n��ݵ<Lo/=T\!��cX�wT/�y><�Y*�1�0�O9a�R���禼�hW=�?]���N��MW=�l��W=�-�6m伍̑����=���<����=�}��=�*1=y�^���g7=�a{�,,�Q�N<��d�-�<���?=mt5='o*=RQ񼡈�<`)P=�y='�Ǽn��<}C��f�o��E"�:M<�֤�셡:c�;[_U��8,=xn9�DSZ=�WN�K
R=��#�j�|<��*=���E��;%]6�Kр���=h<��u����t�;��w�gk=�Px���?�l(��ЄU��WF���-=
}�<�Z�WRj�m(���r�q/S�h�+��7;���<oX=y��<�����������X[����<�%M��3=p&k�+Z!�SV�<�a����ǘ<�+�d�,=�=q�r=b?�<��<`97=�E@<�t��|�V=[Y���=H�=�&�;��=8�ͼDu��Hf��lO�� ��'*�1�<�7/<ӝ���1�=�@>=7q׼�<�.�(�#<q|U��'.=�f=�\���ٻ�;=;��<?'K<1��;��N�O�<\�.=����8;�c�ȧ��M�C��7�:�XV=�?G=�$�:�<��7��e/�>�P���=I�j<��=P��<�v:<� ˺�(<�n'��yK=` ���eB=�YX=�7	���ҺcU=,N"=�V.���	<�P=?+���*?=�h�<Iz��,�,��<��<����X/�A�E���w�QF;t�û�K��l��<��<���l�=�*�߼��	���y<2�:=�v@�{�w���_<?F�NiZ�r��<,d=T ����n=)�7=�_<�e~�U5=�ؼ#kļ�����*=k��<ۨ]=��=�f=舅<g����:=��_�f����<O���V�e��<��X�H�%�� ����ͼ�4�o�M��h:�+?����<���<��7=�3L=�.�<�2��I�<;�,:�3�"�q�^3=��4=�,2���L=�	�%�꼪m!<qտ<L�;�Z��=��Q=�F^=e= e���0�<կ'�ӆx=��<t2����?=�
Q<r9��X���E<��h�<�&G=}�0���;<s��^�`����;�0=��{�:�{8=���<Ձ=D�>��}X�-q:=��<z�ѻ�^�P6�=�G�/�$;M�b=�Ҽ�>��,�<�
�<!�8���u��e=%|@=���>Y;�z�e�YR
��I���>���n=�k+�k��K=��
<7��<)T��Ke�* �<� �:ε�������J�;U�)=� �<n{,�$a��@i<�ü��<�����0=�3�<���<\6=��=cw4����3��<�m<��Z���:=���k��;b5e���u=�����$P;��
�C�:��A��Z=*Mf�����U<�1���G��S= -��D�<��b�i�<y�K=5���WW��_=��żvJ<���<i;��:4�=�~�<U�̼6�<��T=#sE����<�P��1�=���<���t�;V$"=ޝ�Bl�<�΍;�1,� n9�5jo=U���h�<��z=�'u�jD;�����f�׻�3�P$=��<k3���C=��O=�4C�� P<4!g�%i]=w}c=���<�gj=��Z�S��+�<S��u�<S.�<�V�b=E�^2�"!N���v<$i�<X�J<�n뼮�W<3���v��<.ז<&��<�'�<��=��p=�2����͗<��?=/�d�iOg<�J����C��e;�<��*=�R>=�1�;�̙��	Z��� =Mq=���`Y�)�?���J<��U��(=f<�A."���8=��M���9�� ���[<I�㼲
�=�2c�#S�;�=7��Ҫ��1�-=��-�M<�<��%=��.��^�;}5�2�����k�T=�Rx��c�E߱<c1�b�=v�케m��w�l��ک`;0�Q��'�;��v;�F;ۥ=��k=�
����<�>H=�(�vzҼ���e`=	�=��!� o��,��m8���<����G=��t=c=��ܼ7\�<�˼ؑL�IH�<�/��3>�c}�<��ݼ4�M�M�E�>#���oa=I�<�(M=��A��OM�H�Ӽ�
6<*k<#��<���B9R�#d�Xм?��<�i�<5�����<�#�P0(�{.� +L�55�u�:�@�p���<=�;g{C�*#�<qL��H�=�!<q���G�X:�m.�<m�<��B=�j<����i=v���}e;����{�o=�='�:�7�_�'���<�==	��<��1�f<>������<�Ҏ<5=2�,<��-=���<LVi=8&?=�'���<}����Q��s0=!g,=��?=�%=Wt�|ŕ<Ģ���E�=�+;52<b��;�s�<9^f���<S��<R=�!g�I�?=�U�L�U�����漎������<�,��E=hZ��G=o!�<;�?= [��9����<�߼����X:<>ډ��#+=��	�{�:z=�D=1�-=M�"�l��<��H=���;1���`Y:C�*�~L�<>�����W=M֛<ݿ�DE	<A=W���^��+�<�l&���j=�+�<(�ԼA@S�!�g<�b���c=�B=��!=��<�M^=���Ys���d��莼*�2:d[��
��@���0��"i=�Ya�.�	t��_�2<@�n<8�M�o.�<β�<{O=�_�9��;o;<V;^���B��#�<��&:��'�'�:�޼E�N=�=Ӊ]=�J�� ����#�B����;/[�<[w��q���R<��ż�қ<?=��^�=0;�<�;�$��<�,��2�!m��`�;QU����=���<nJN<A�K<􎤼�`�e\+=�g���u"��X <n�@=8M<��Y=�(ȼ�N*<�����<�M;�Zf<tD�<d��Ʉ=\c	; �Y<��c������y=|��N��:�ax<<RJ=�䜼gj=N�=0���ا�t�=�:=��>=H&�<����Z2���Y<X B���O=��μ0�&���=�̻�%E=k��۩c�\�<+�����/=�qF=�[�<'ۺ�"0=��G�5����F<���<	L<J�<�#��gX<AJ�<	?��7�\��{k�05���c<���<;=��J�񿾼l[=~��Ot��V=�<������1� ��q��!�<Xԕ�V'q��<)�d<]q�<r�����������F=��=^{O��O����U�/<2��x
���%=�8@=����2qR�S���뼰p�;=�<���:��<�f��6= L�<�����O,=T���ż{;J=�1�<��-��ke�C���=�*)=R ����Myͼ�;����$���<-��=遼Ҫ<	�<B�	<��g�O�t��9=��3���0��k�_`�<V0@=��U�ԟ=�����5,���(�{\����<��9=���ռ��b<��x�J���K<�\��|X=bK<	�F�V�k=��޻����0�<}M��V��E;XBe��K��Q ���H= G=��Ĺ~{.��<��!��'���Ce�9�}�H¼Å�<�t�<���;�ݳ<�ʠ;y/��0��g.��8�<�=���<#�5=Ӟ=��5�N�=d��<�X�;e�=�i�<��ͼM�*=p���F�|<X"'=�9e1.=�ȼ��:��=��:��û��L��z=����4�4<V=�q.�����4<I�ټ�%
=��<+������NA<�G=�&��wi=��j��hd<�=��O�C��;���+`m<���Zl��;�Y_��J�;��*=��ڼ�Q����;��z���`��%�<��m��Y���T=S��+�s��Ϩ<���2,=^`=D�9<�,B�X3=����=�n�9.��<��e=�K�<g�Q��tzw=�H<r�Z<Д׼�y1?;�5t=*7��b=��8��<%�r��Q�X�^�:�|=M=ZSe���;����,4��^�1&%=�uc��=��'=)��W<	�<�?�B׽�7�\=�-�[QJ=�i1<c�<�2�\�=F��.��yYs��3���m�<���<W9�<q=o<a�=}�л����L=��(���	=��L����<'鳺9���;�=f��{���v�<
��x"�<���<
�+��{�;�H=��S=i�T�a\o���J=b94<u�=+l<�*s����w��N/=��;v����m�S���n�"=��<�3Q�3C=��=MS���N��Q���X=C�[=.��<��~��	���K��g�=7�>��4GO=��"��\K�h�K���m;l��;�6p���l<�C��QU��9O=�w+���ŻPB7�w:ӻ7�8;ͩ�<y2<��2��AOO�.��u�<��i��l�<r�^��_�<Б�<s�<l舻+7=6Q�;/:����j� �
��gd��>N1�r6��(��{�<�||�c��A���3>=��n={r�D71�<�<n�[<4t����Q���`�Y&7<rG=�$�
g=�<,�Q=��-=&* �Wj<��<�B�<2�>�4@$=Ҝf��ż&��;�1��������9弇�j�~p=>Nʻ͙��F=Q�����b=��G=y�q�v�<�x����=����}�
����^��/=G4;����4;��<�ܫ;�b��d]��C�<�����^�<3(��=�=S)=/\�<��<�O=pK���`��P=�N�:B(=��D="wh=��;��c��w�<9���6< ��|�;��<�׻)B=��[���=\;=k:�\�����<�eV={�j��
	=�숼�쫼*�?���!����IFB=��u����<t�<zX=��=c�z3�;_k=6=;�
��B=\uK=��<Ce=2;�<����l�F=� ��o"�<s{*<��C�8��+���s����<�&����@�sz�:O9��B�w�|�8OT;}�<=�v=C=&�-�Z;��b��G��	�Ǽ�fR�'B�<x�t�h��<	�1=��0<�����L<L <��<�U<� �=t*���C�oD��:������ب<\�C=���;?�V��j�<�n��U�<��5;X�=<�M9=(E��gѫ<e!C=�B�:>=zϼ�s꼍����HP=�&�<%�v�:=)��<;\)=2y<=�
����μ�\�����d�<!�h�li<���<٬��z%s��=l�<�P5�l'=`$Z=��(������N��Թ��ڼ;g=o���Q==v�ż�F��ט�u��;nX=�=�1'���2<1"=��@��<�u��O�<If�<��4�P�B=X�P=�(�<Ik����<�?}<l�i=ѹ/=��0��cL=͂���r<:����<"�%�W� �g&6���<��=��4=1������=��<�*ͺz��O�<�vp�rC9=1�=G��=��߼��<=��ּǘ&=��<4b�G(S=h�K<	9�<|�!��<^����v��V=�}�^�=��=K�=T~==�6=���<���XK=!(�^�*�ۺ �d��<�����.=�x:=�~l=
br���o;�=�{�;��N��Ag<Uc弆�S=�¼Q1<h^
�Џ���5=�+�<RU���9=�Se�D��%�=���i�j=F����I�����=�ڀ<�,���9+<j�?�f�<�ݼ2R�;T�Z=��F=�G_����.�=���N<H�Ǽ�<��p;�?==AK��v���̼m��f=oW=f
s�p��=Wb=Q5W�"J(=z��:kM�b �<>9a��0�E�#�U:ֻk�C=�3��j��m;]A�;�֏��N��A@�m�w<�e<�&�<�]ļ���<�J�VS���ї<<����;a�<������0<:�C=��V��+���<<�P+=��o<�`ƼF\�=�N&=������}=���������O��=�z�<�%X���]=�BK�~�r��[�
���ZN<��-����:4v�䵄�3�D=��O�:�d����<N2�<�-��b'�<��<�b���E=�1�� ^=G��<V<�X�'5�3�q<�6~�#�c�y��&&��}���#��	��;�����5��8μZ/�gT=	�=<�A������<�D:龋:�嘻��T�W�==�t<@Y.=�;:��=��<�����><wAh��S�<qa=��<]�=K.M=���<�[�e�;Aj=0Ip�l�8k64�rW�=���aM��NR<P�3�T�<+��˦<'�C=껁=C�!<������9=��h���<�3�;H)=�h#�%�` �Ե=d�
���w���K'ܻ��+=V3<��9�c�1��Rr=b���O�,��f6��FK��MC=>Y0���<��=d0�

=[�K��!=
ٶ������=K�<?.=���<��^��7b<+�<#u�]�~��<��=l�F=6��<$_k=�4<�*�;:��;Q��<E�����W������e<�9��ƌʼ��O�Q�������R<�@+�mG#����:1b=�W=�h�,�<�Ǽ�� ��C�;,P��:i�<6�W<
�.=���Neu���<ruV<r��Y���=�A\���=����W�Y<��@��=�fm= "6��ݘ�Æ(=����<:���;'<�T�<��<4�.��>����<ۆ%=���:ߓ�<��+���ɼ J�<�:Լ�(/;� ����<��B=Q�D��<:�ü��;�b"=��;GҖ;}�I��s���߼�kY=���g�<L�j=S�=�L�<&�^�$q<�9���j;#�E�'n(=�����	Q=��;ʊ=m ]��5 �����F总������<���1�<-�C�Z=��[<���a�F=��P��W<e��<=���uc��C>=��̼6h<%B���{=�㋼b��=��<��M<_HB�[PG�����& N=�����ZD�q�=��}=��'=+�9=�U8�u�=���<�= l�<���;�K���*|<>��SH< |=y�p2@�]����_�;B�9=?�=�R�<��I��1=�q=��<����^��<� ��R;���綕;6kN=�ы��������4�}?��v�ɼ�;���<#�����	=q��<: =H� %��5/=�!��L������U��C��_e:��v˼61/��J=	s=AkL��S�Sg9<_�f=G��;����n���ͼ#E߼�������:��)���^��e�j+�EF=O����ܻV�.�Yr*�R���B=F��<6�=�$z=�hY<�tY=��;)v�ΐ��pb�e��<8�F=�:����R=��;�n�<����Q#��{$Z�����I�<۱Y���9���ܺ.��;3k=*ᶼ̖$=)_b=��T=�n�<�>�l<��-<�/��'%=�N���}��ƒ<y��;.�����:z�#�r�S;=��<��%=�G����;�6 ��*i�n�S��$���߼ǎ���ż^&�C%�>������aB0�(��<��	=2~= e���x"<�;�<VB>��j�`=��!=��p=��t=�u�8�p<�&t=v��<^M뻣<_�r�n=\M<ÕW=�.�M�&�b�<�>�<�F�&f7��¼�"��&	�eӺ<!x��z��O?`��^=0�(;��*W=��N=U
=��U� ���Q=�*=�8�<63��	�f��}�-jN� "�<W`�<8}�J�8��X7=�	/�z�o�`��l	ռ6Zl��!�:^M=�G�|%��=\^�<4 ��a��<�<PC2=���<��0��k<�>#<�=2�K�{���G�4=�,�n�����>=�-d:�+��Y�<p2��R�=�=\�s<ܗF�8�Y=
d�;dD�=�=.�:�-�l�<�C�<�$�<-��<��=�l�<#�X=��ɼ�!��(m1=�:AɎ=vt<�q �	���oH�7K��N=U�"=��;,��<*7�<[g�<����UV�o��<b=�;=Y��hު�J�/=��U<�޴<z�'<T������դ��j�<��»��;4=�mE=�k���I�g�8<���zb=v�4��S�=���1�H<ٕ';�1=�%��P`<���<G�6�"Q=%*::���M`��G�<kw�G]a��;�� =d�=�A=��޼�6��H(.��P���ߺ.-=��\�+޼�g4��Ϝ����<p*��5��8�9e;5u_�%@���I=R���d<�'��T�������=Վ4=��<C�=�:S���=�S��+���A<Fx���I:P詻>��;���=~���"��;��:=��\=�E=��ϯS�o���U<RЯ���#�<D09=�ȓ�Nॼ'>>���w��, �h�<^D=�f�<���" �;o���*>��=Ŗ�̶`��� �.�<瀜<"4��=v�<%� =H�=�7k<�U7���=��a���C�b=��=�z�A���|
=Bi^=B4�<����T��?)�<tt������<)5=oS:�f?E��@(<��/=�6<�Ӂ;�
I=�N&=��<4�N���0��/J��3=�F!�-F�OPu;�-=�2�;մ=��M=�=,R�:�U=�;�<�)=Oʗ;w���*<!��<��Լ�VO<h�<��0<Hb�-*=�S�<狸<�g+=�g&�^<�h���!]�=�8=D�8=�j3���l=A{�<ʵ<P�;AȂ�H\�=�=O�6<��<�A����7=��X;%�"=��7=���`ŵ<�=��=J��;EMz��tU��+� u�����{��+�'=��'��kS��B=˗U<�J~�+Ѡ<�/��ؼ��<�4u=�.=�61=kB�<����0�w;z�<hQu�.�I=�1R�,��8��Y0�Ǡ���Χ�f�(�>�=v�0���<QiC=`�;���<Fh�A=��^:��,�#]Y�[jA�]_�<�U<���<}p<@�
=
(�<��=�K�K+T=�?�<7��=����<T.~=�G��f4=���<�yS=����^T�NFc��H��p���<�s�;�?���a<��Q�.V(<�r�;v.�<~(W=B����k�qvp������=N��=W��j��z===ar="��>5�<QK5��z=O�!=:G=+D�J�N=C7�<�=��-��ޣ<r�)�	"!��5;�{<�=,��g==�μ:użA��D[ڼL��<�k~���<
�����Y=-]q�����^=9x<���<�ĺ�(����ɺFX6=ߎ<��8=���<ȼmf�<��K�>���g��J"��?\a��#�(^<�I�<��;@=<ܼo.���j��~ּ�a��C�<��#=��H�<�)�Bni�<m;�RxY<�)������v�6(<x��<_c�<p�*����<߳���9���b=��*��"��i�<kf7<kK��jڻľ0�ң;��;�.=ۛ<#R��Oԙ���<���ܰt=b�]���,���"=�&)=
�v��F�9�SܼM�o������<U�����GӢ���λ��޼��[��Va�'8l<*�.���7��*+<N
<͗=� E=UK=Z��GE=�=�-�i����� ��D�;q�f�^����<��iY�<F==3���͔��zM���%<������:�L����:=k����<�<	=X3=<$<!6%<��"=Dq'<���L�b<}�1�N=~s�<�5<�W��hn;�y.=}z�h�)�+OB<� 9=�e���#=8�G���~��B�<�NU;�U���=\�j�[����Bq�*f׻�R=�ɪ��8E��=��C����;VY�<���<GK=��s=����ҷ<�h�<@"0�q�缡<顬<�<3o}<�Q=�5\�Z�V=�������I=s[g�:1	=د�<�@>=��V��&<c��<�87;]Ӷ��"�	�\�Jϫ<�<�se�0��=V=��[�<��<�,<�wn�Y��	��80���a�jl=np��eBL=�G5=�~1��e"=��C����0z�:}W��rLg���Q������@�Ƕ����=�);��n
=Wx=�{�m��k@�^r��"⼨�e��w�;9��;�.N=����=4�=��?=]�$���$=M�=rA�;P���W�dF��;��bJ=�tg�)N�<޼�<ל�W�p�\�D�Tg��|��^�<��x=��(��>K=�:V=�4>=��=^��<�����N=0�=`�=q®<T�T=�-l=d�_�:����/=2������C<e#D��j$=Ɍ?=uf<x���S��I�6A�<�I�~&��ք0=]@�<���������Ļ��l=,�(=���:�]���<ûI�Q������<x��Zv�^^�]�	�H�+��5&�1�<Nm����s�>�Y<fV�<t��D�4=��i=K�2����� J=��Y;Ɯ��R�<Z��;O�9���M=�7��\=�_f7��Q��g<�$S<]@�&B� {=UW�<�ڼ��G;U$y=����E�[*��S�<���<�ۭ����=/�W���==�k���D��g���ݻ�G������)���b�=�;�{B�<���޳<�/��r��<� ���C=k=,|`��	�;"�1:��E�5̀��� =��{�Dr ��Z��볼�-=�Sd<�酽J0���
<x₈<�����-��{=��<���<D_>=���<w�K�|=�3��ޥ;���9��t��`�<���� �f���(H�<�2$�x�z9s��L2�<P�?�q��;��1�W�ϼ���<��=�@�D�8=��L<�.��p?c=��߼<�λ���;uE��@U=K��Z�s�p�c=�������j5<�X��.�9*!=�&O���=��'��!'=�0����J�w�<��Y��� =��={K�<M~=Tٮ��H=@a�<s���Zj�n^�b��I�<����@�;3Zܼ��̼]�<ˏ��P���M�;�p9�R��^$=���<���a,���r��%���1<�!�^k���_��W�<Ǻ5=��\��&ݼ��=�Yd=m��w
���S=�g��*=�ј�[�<��ּ	�P=���<�y"=�L�7=1N�{�F�4�
���=DQּ���<�'���׼��O;���<Ǻ�;�S�<�i;?}�:"�C�G��:�<=�=��|<�φ<^�8��K#�bD��8=f���<�,=��<�@���m�9mV��'�<ߟ��3�3�$�����=��ؼo�E<�&6=@��<Xżj|��W��?�8Y=W�i=�{��G=M�����,=/�Ⱥ��<t:��0Q=���歺�+�<]"Z��.��'w�<�E��%#=nK�2%e��?��ao;^�'=�u=&�,��J� 1j<L�0;�����c���8�;ʇ����<}�+��\6=U� =�vy<��M<�y�0�-=Ȕb����$<=��%=-��<p��< �n� AZ=C<=�; �M5=9<i=��A;<�<J@��߻�ܻ��a;�2˼�5{�<�==��3=�F=a�ܼ����5+���|�̘~�I��bv��if<mdy=�d=��\��a<=�<^nѻ��U�	��=�ջ)�I�Y�
��U��<p)���L�O	 �>�<��[<7��;�,�<>O8�k|=�/z=B!f=Σ�;<�`=����#=�hR=]rT�����F==ε��|�P�ͻ�XU=�>=��P���Z�f)k=}��T�U�[�	=�_Q�zsJ=c`�Ұ�<%����祻���_�Լ�&6=�pC��MT=��ễ	s<��μ0U�<�KQ����<��;e{�lLh=&I���	=���e}�= B/=y���#"K=&1/�[��_.�g��<�5=�X*�8�D�Y*=�쉺5���I�>,�R:V�h>�<�5�NT
=p��=��<>i��.�H=V�=2�K�s�/�X��<�gh��I���̛;CKʻ�,Ϻ�y�����hA=88n�.&,==�=	�%��zE�����YkB��K=E���[I��B=<>�N=��!=��̼2l�\缇���̼~�=������ü

��7<�yＵ�R=i�m�����3�":��=YG='乹J�/�^C=?���^�J�c="#���=�bQ�%��j<_�F<�����>�]�=�9���	=3�˺ѻ-��|< ;��\$i<J��iW�v�.����U1�<̝�<�<�
=/�;ںE=�+ԼE�����໖f��8K�<��O:�4����R=%��<*s]�Q�C=+��s���}�}��=�
�(o0��i<���<
JI��S=Հ2=i>J=�1t=~�=ޮ˻7��c$���;=��+����;=]=Gr�<��p=�U/�ҩ<��_�SQ�5�	�e�<=rN;7��2n��˟9�z<���E<)w,���4=~����<ž+<���<fQ��_E��5�=Ò�<��{<SO�<� ���X=_�:c#�;`7��l���1�܆��Ǽ��7=�cJ=.wY=o!�%l�<�][���{��N=K��\�@="ټ����T߼���$�$=�ͼg�� �J/��d:��^MS�B�v��6�Z߻�V���=�߻��!�@=޿=R:"`�;,=z.~<Yi�<p��ST�!�1�#=��吼��=.�ڼs=K��!�<ş�D���"�����W:�{��Κ��oW<f�=Ǔ����C�;R��<A��<��t��k ��D�ps5=⬺q�e< ��Er#�zw�<ĦO��=�G9��(U�ݧj=�,�=�WO=�<[�)N/�=�X=�~<��=�e�<�(��\=����<~�x)	=��r����<��dRG<�c޼�aU�� ;��8<��C���;u%:��U��ʻ'�4=`i#�����.��<�<� �<�t;�7.='cѼ9s<>�"��&�<��/=Sx��/�>��ؐ�<�����;R�h<����7
�¤;=�j�=�o0<(�+�A�<�ԉ�EST=�V�8N�^�ռԝV�OO���1n=��[<N�ؼ4��<n=%V��:�;a��<?�����$�A��x=n��9j�<0�|;OW��͖�U8S���J�j�5|Q=�I=ww��J<dhm���b�����<�P=N ��)���/�<oѼ��;�4�� 1�)�<���k��Ǽ1���	��M)����p1��K{<�Q��P/4����<�Q=�e=̏���/=�O`=�U:Ӣr�5r�<�2<�34���=��C=>"=��;����=��<�}�3߼azv<he=`n	=��<��Ƀ=O��<�{;��;��=�B�~u��f�<��9"��<�^�;���;g��;cx]�>k=P����<�SG�Q-Ǽ��&=��;F�@��il�CE=���= R=�#�����<ϸ�<x�A�vn�<�6��`e�᳂�i�[<hn0�~�=������2��D�<��=c�<�m ;Mw����9=��{=ԩ��Fs;^��;�n!���Z=��<�-o<C��<���; ">��=S�<�0=�YN���z<x�@���%=&W= H�UҎ:��?�<���;ߊ��m��6
�<�QH<݁<M�@^8�����8���<~)=
�R=}T�=[>]=�'a�
�<ެ���n<]���= �ơY<0�1�q8��x�r��.O<B^�;��M᳼o>��6?=S�d<ь�<��=��Q��C<�=E��ڼ���0�P�	8o=x�d=�
���,<5�Z=��m=�Z=���<�н<NF<�67=Ʊ���$����Y��j��`R(��%�L_�:3=�4=�ņ=��%�NUJ=�鐼ë��tkX;R�"= ��zY���%=���P,=$�=�^3�&5��v�+=<d�ޭ#<��[��\���ӼV�����b=&�<��v��	j=þe=��]��Zu=��Y=��&=�=�Q�<�+�<�=.Vc�2�<=jy�<�N�<��<�,	�Т=���������'�=e�n=�G��Ȍ*�6rj��9�<?���v=HΩ�	Ý<Ć��4]=xu^<�-;rE�<�ݚ:��,=��8iʼ'5,�z�<�- =�|Ƽr49��}<�lt=�z�<��!��Y�͘=����<7����°�9������<����1$���=5%�����6��\�<�ہ<�x=C!���J;IT��|F�ͫ�<�T�w��<$Z��h�<s��<`�M��[~��rлj;��� aF��C�c��`�c�J�m��z��<��%=z�t�H��<�y��?����3��$ݻ2<��J��<p�ǻ%�=g��L��<<[=��μ��<et���L=�\'��C���1&<XK#=f?1<i9��}<��U=�'�~�<��<ݥ��mi�=׭�<��<��[�)�<�==��߻�M�<� ]=�4+=��=ѣ��Ƽ���8�xZ=6�����<g�0=F�˼��<��-���=�[~=fb=�U_<��<aY=��:�R�M=�ί������T�5h��=8P�=��ļ����/T���^=f��:�:=�2��r�#�H�"=����l�<��<�/3<�S>���R�45c���;P�~;􍕼+͒�H�9�{!����y���o�=�8hR=o���?=ы��eW��v�9vz���V��y$�e>ϼZM
=�iI���F���_=�$�ջ{<ɱ;��b�<���<^U=�K,��>����<@���=��;�L"��=\�
IV��U"�D���XT$=!Q�j�4�M�<�䞖��V;ύ���F=���1n�ӻ�: �<�t[�n�y< �<B�P=��#=����N�?=;@!;��<�2�<����y�G<��O=�Q=��=���<�g�	?�;��S�~܃<&]^�C�T=:�;"�у��˽�*�3=Z��<S��<]=�S<��9�42h=a�==X,<E���*��5=2�#�^I=2��4P���[=���b�X���Ӽ�+l�v����_�4,=�C0�򥾼�a<��H���,=��<^!��+o���<>�<��r�1����
<��X�F��<�s�<5}�2��0"ʻ��==D+�_��<II2=N
=4c='�;;2S�;9�A=�=�=T��<if=�AV��&<��C�<��5;���<\��9zq���l���{��Q#<?͂=!eż��;=��'=��r=o!+��A0=S���,`7=��}<�� Pr<}6�H5G<&�C�ȻQ��� �RbQ=�*6�x.4=�������\���]7���<:T�ԓ�����<Z_<hڿ�EW�L������nZ=�yk;����=u>E��=�<�N�<��Ƽ��<�1�Ñ�<�G==K���=��E=�
(��M =�`=�[� E�Te���2n�	��O=ݡȼ�'D�����.=�%A���?��=��n�=a��g�9�h�SJa�<{X=�nU=�	�p��%�]�M!+<s�K�ńͻ/=�a=��%=�n =�4<iE���(�޽��tSu�j�*=��P�k���e�<��8� �B�q�i��4�,����k��L��#�=#=2�F�D;�MX<����R�:qz�<w8+�0��<��<s]��P�<`O�;6����:�=»�C�<�S����z����h�C=��<���<ZG�M���)=8<dg���K<��Y<�f�<b	���0P=��v�lt6�Gk<���f�U�<����B�="�<�`��0m=���a��<[�=w�D�`�ڼ�x=L���c<�h�<����L� =�����3��v�L=��A;z���4e�<12=��2�~�ؼH�Z=�݇�O=���1G�<K3�<�U=ݲU=�z�ۅ^�R����E��63=;I<�79=}C�;ȯʼ_���z~�9�U=��;xZ����<н�<Җ�����<����=�~�<ƚ0=��f:�Um��,=G�4�:^��"=s�=�M�� ��<s,��(�pt"�g� =��!�%Z=�����:�fd��aT=�WP��^r<w�;�4�< ��<p9'<Ӑ�:ڹ�;'_]��G�<�w=���<�H=6�=��f/�<Z=R.���9���a�m�S=�l��"�{<3; �~r���U��\&<(�»�[���l��S-����)����<#=�q�<Q�ȼu�8=σF=��H<	�:��qP�p?8=��;#���p$��wἬ&f;�ٽ�;*<2�<=����+=����a�u�+#9�� =/؅<��_=��4=��q�7���.���v=��U!=��Z�^%)=|�4-=�yu=}��<x<.����u��<.���ퟂ�[���o��G��<�V��ӺG,����Z=�n==p��;�C,�B�9=��=���<[�=�={FB�<
==p
<&FҼ��Y=�>��r1=v.=ȁ0�4��3F �k<u��<?��<6���Y�Q���=k�,=z���C�����<�k*�">^;$�b=1�@�����'���l=&�D�@�<�կ�A�<qk=AV^<�]e��AI=<RC=,����;����U�=�(q����K�uo��}=����(������p�k�E=�̋<��C=�f��ɸ��z9��=?Z��/�v=��=��6=��8�q�R�,��v�C=��E=����e=�����=��;�,;��:��8,�ԛ��0= W��S�d��W=�� < x�|_m=��	�7��=���<o�a��u<�mϻ}�=�eN=6���)����wp�G�<��=��U=��3���#=U��;|i����;�ʕ�.$L��0a��K�<�Π��N�^��U���M�Ҽ
w����<"�l���=�L�#�`�d=/�<B�(��4<Sʢ�E�iՋ<zQ����P=�y%<
�b=��<���i��<7��<*�t�+i��.�J=�Cr=d(�<b0=c]��&��C?�uj=�׼�:6s-��P3��伃?�<��'��)��ʀ=�==3=Cl=�<*`�=9�;== �X���:n<�=I�<
��qG1=�����?=%�<υH�.8�Y_����gNj����P��<�q=`��<7�;B���h�CɃ�@]ϼS�N=�Q���ȼ$�::��:�')���|<�����#}���.��X���T�<#(=�#�}�Z=��<Z�=�t<����Z��=��X=j=�������T�X"��L=	�<�.���H���ɻ����%_�Ւ0�lp/����W<	��X=%'=�H =��z<��H����<)�y;��g<A����O��]\��[9���� �"===o�Փ��h���d%=q%<�m�<�%=Z�=����<��=��<�Y���G���5=~�ϼn�<�r�<��
=������<�UL����21=�j�<ֵs�B�<�2����;Lr=����F�H�ϼ.�<��=�d����=�(�9�X<�uQ�ť<�2��<`���U=��,=��0=r��;��=B�<�&]��!L�y1^=�=9X=�,=���-����;�ך<0DB=�`�K뻞��<]�(=	+n=��[<�����N<'i�<�X��f4R<�=�=q�-=��ؼ0�=&�H����x�%=���(M�x�����W=�:=rf�<�Q=����+<93�;9��<H�5��{��-�G��2m=0j�1M<����0%�<J�,=�&�@���0�����<�Z �6:2=�3������ZA����e�n=�7&=|�j<A���V�)�=%�@=�)j��Z�� 躰`7=#�e�H��;��.�p/%��~=#o(=q=X
=��<t�=HֻW1q=��<b����V=����������Q��E�	���<ϴ����%�lv.�׻�K���=Iu�"�=�{��iK<@ŉ<żX=q���z<;�c<�G�<D_�1wA<[�s=�'<oP==-�<Bz=_+��^�Ἢ>�L�h=�+_���>�%:V=)0)���,�\i����T��yU=Ȥ}<$
�<Ϸ�����<����"9���i=r�ǰ<�����C�<�O ��+���'<L*M�/��4z_����<`�л���<p�¼��R���2�<�8<b�B=`i(=1]:�=�`=��	^W=�+w9C�
�Ǽ�&���=��=�Lļ)9=%���=<�1��;����S=�����-=����g��eռ��H���ϼR7S�"`�<�,�9���-�<�7����=��=�C�:<���<�i�প�6�9���f<��"= �=<,�������<?�So�<��S=͸<��'�7�j��2�=4]�<ho�<Hr=��=\Ӡ;�R�<Ej���Vɕ��E�<��<���<�Pb�z�C<�a�R]�`1v;G6S���Q=nR�:�B7=JU�+����L;=�f(<�8����ٖ���m;:7���Z�<f�=�;��<�����
��+.�.��<xJ4=8<U��<��N=3E�����<��ټ���;V!m<� ּ[�=�zC���+=d��	�t���<�B�����4�=�fe=[�P���=SsT�,*.�� �=>�K=d�i�k��<�һ��ɼ��o�X��iS=���;(=?=��޼�1=�y�<Z��;XIY���:�������=>(v���5=g�=d�7�h�Y<Ā�=��=%Z�:�Y)<uaT�������<�I��;'Y��xe�gK%�o�n;�7���̼ywc=�}</�o�<�Z'=�D=�N=��>�C�]_��e�<��מ����+�<�?˼ȴ��K�]5=�_�=Y��o伱�t:*���8��v�:�y�;�.�<�*��5�.���9ߢ<��Ժ��<oRW�y���^�<���<@����D=tD8=�"=ގ�<�w<웬�W<8��귺i���X��?��, ���ɼ���<G!P��~�<�_^=�n�<��������/?��V�^d<�;��X<%�m�'ue��z�g�7�$kV<J�<��̼>'6=/�����o�B3��6�6�ݷ=H-Y;@���<:=�[�q;"=�B;|��Aw�J���
7��z�<�����<�j���7:�������|��i�<�-=�`.=�qS=Fλ;�]��86><�	`� �=��!�d8�fCE��t���b�<�Y[��u�;�D�<v'^=��'<.�=;>�=� L<�fǼ�����-=���4`�;7I�<�H=�n�<�ӭ�+�<t�=��=г�;8B2��N@=p��s�=��|�سI���¼s��<>!<�oս���@<��L=6�X�ԓ�����<
�X=C`��la��8Ud=����%��=����<N��V�,�K�<V�=:�=�V�<{F��h ��e;��.�߀�;AԠ<CW�<0+"=p�l=��`=�/3=n]�<x��<<W�<������-����8_(F�V�G�lO�ŤD<GX������=���K�G�� };_	�<�w¼�C	���<8�b��'�哘�IN�;���<�S���\�&��s�<��뼿��<��C��O�;��������<~�ɻ�r2=~|�;ƨb�G]=�`_�q� ��P�<��+9��`����<�n��"x�_S�?�~%���Yj=uw���f�<�1� �	�H��q�<Jz�;����K$�<#*�;�(4==�I=���U����W��=e�a�Q�R<v�q��H�<r�ܻ|V=%�L�>��<�=��ܼZ��<��=Lh�<�N=]sg;�����h<�|�f:J�r�.��r#<�+=[X�<i��<T�<_��<N�'=��<1D���w�����z�a<��d=��Ƽ��񼥔<<*�;w	���ռ���;Bْ;j�{:����Q�<�,=XZ��ۼ���;�{�<�{�Ŵ7<��ļv:[�";�|�����p�<>Q��0�ט�<��x���K=U�&=��<��=�v��v=�A�oM#=��]<��H��r=Dl�?�=X&��QI�v#�<�/<���<rU�<�S<M����w�s�=�©<o����O7��ڻ��i=�2<黺<-�<uQ˼Ɔ<�tj=E���k(=J�=�<<�μ������ �}���&�<��d��܆��[��B5<bUq<���<>+����-R =�\/=�T���!��' =�Kf�`Z�<�ı�◊=]F����=�=�+���<��^<r���(��<�N�<�b��N"�R��Z��<{�-�q6ڹf=ᰭ<şk<�.��rf�/��<�=r=�S+�dJ��$(=�z��Q�Y�<vPǼ����7��<�	K=\�9=���<S5�;;��<z��<V��m�(��B�<A����[<�3�'j��	��<�W"=��h=E�=��O=���;�3=��=i�F�j�=�O��Ǽ �'<�"�;f��<j�z=z)���X=�)t���<W��<���;���;��)=Ra�{aB�
�1:�un����;���<JH`=jg�<(����=�+=�s:��c<;��5=m&���=�u��`��鏼���<�r=;3= ��;Ĝ?��<U)�;^��Y���t8+;V�U<�;b=���<H=ޱN="��k�=E�����;��ļ���a=N�t<�&��v=;��<��H�F�X���x=2@��+(=���<�|�:�/�9�=Q�$=��E��Sy��	<������<$^v=�
=&��<I�1��-=��ռw�=�Z4=��=�qa=-˰��
�Ez,��u��۷^�[ɟ<v����@=\o�h�!���4��؊<V�b�؞�Q��<�%=<>�a��=����佋�V=$�����<J����2�C嵼��9��
%��8=m¼<�����_���^f<	fz�*ԇ<�������|�<ռ�^'�Y�<���<6�$=�y�}�R=�� =���}#�<�	;���<L!�=�
��K�<��|=Ͽ�<��;і��4� ��<�^���=9���<;P�I<�w<�J=�@/<�Zk�D�<��*��P$��&��EE�<�NA������=�M��/���M��&{<�^��l�-���A=xy��{=0�p�=�Y�	�R<���;B�+=@H�?#(=���B�����'������6�=C� =��=��5�X]8=a�VX7�W1=��ü(3�;c��<�A	=�l�<���=�}��� �l����P=HƻE���)������C=�'<��ػN9���/�E;�A0="�L<&���(><P�C��j���V� ��:7��ߖ��ーK�N=��<A����h��1;=��V���3���=�cs�ۈ<����m��7��G��<d.==�}=*ѝ�����Ե<���<�;�����$<J��c�"=���0�B<T�=T��4y;�<G�߼UD0<��e�ɼ�bW��l���p��~G�L��;�L�sh= ����s��;��^��Vw�<���;�/<<��<��9^�<�=7<=lb+=�v;=�N>:+&;c�<=�ռ�P�<�i)��H�<I<��]b=4�</�y9إ,����2[<�;��v/a=?WA�bz�<��I<Z+輅��<�߹��;,_"=�a���C;,�;0������9��|��F�>{=Od6����<�#�<|�
�v*B=2\��zBw<�/+<Rj ��'=�n�ӆA=m}���yʺ�m�<�+����<<b�9�0=�r��r4_=�ש��3�<0`5<!��;z؂;B����<��<�I=7iI=A2=
,<�-����<h[m�|
.�Ť�>"=�<w��p�=\��뇽����<J��<m�}< ��0��ތ9�m���n7��Q��f.�N[<��<w��U��{f� F�
?��i*�6�<E\�<�5�:�+��	�<{n<b�<�s
=I����䯼��	_�<�:ܼ�Ҽ
�8�Q�ܼ�F�=���YBԻ
�*����<�s�<��<S�|<d�K=AX=��#�R�<v�����v��@A=�I�<�=h�ڼt�*�(�1:�:�<:Q�<��-�D������;&�n�V�;$�����{��Q��X�j�5鏼��=3��<ɢV�'�%=�`�����4_=� ��e�Ӽ ��<29��<�o<��|Q�<�:3����Lv��X=/ =��P�T�!=X�q=��T�j���C�J;n���g<5�K<�b��p�2=]=c����.�M�(�PE)=/-�m�`=��;��;�<'&�;(ܡ�!PW�ϣf�1���{"=[Jݼr��<��G<ܹC���G;� ���N�L=���E��;gm��	��3�<����ܘ�<ĩ��=�i=�yE=UC缍B�"���d�=*C�}9[=���P���xh=uUZ=]2p��C!=����#fI��Q0=�4=dx�s�f��Q=��D�K?�&��<1��<��=�F<M��<�O�J�a=��Ӽ�&�_i׻���<���<�N�v�y=1
6=&-O<�Q���;=Ȋ�<���;ޑv�s]λ񰔻A+���Z=����=�QU�+{�������,=Z�F�Rʋ��<�;n�v�,�e<NM=���<�*�<J�;5f��0�s;I���;-<�
u�o
�-h(�-�F=2������<G�C=�N= ��<�W<.Z5=*9��[=<Xc�<��]<GD̼��<��5�;4���u=�l<X�J��j�:��<=�{�<�l��a�����=6q̼�yX<�6|����
<G��Z����=,����=������= 6��)#-=�[D��6=^6�<���<���;��˼w�F�
�!��* ���;9¬�R��<��^=Q�<@j�����<8w�<0�T��J��@=����%r=ǔ�����<�Ƽ�9*�с��`6�:Z��񕵼��R�w�o��4�;@�ʼ%%�����n�	�.����}4F�P�j=Q�q��ѯ;ɧ�f,<'j<�="���*=_b ���_=��<;��;%,
���u��2=Z��<��4�&����&0�.9��G="���oiּz�B=�u��L'==JN�:xM=�c�<Du���4=5�X<#~<Dn=��P�_�<�<���L�<��C���J<��2=#�K�2�;p�?��A=�~�<���
�=���<w�
<Yǆ�k��E;[��^�$��a.'��;TZT�9F��N�:��ޣ0���l�cHW<��l��kr=��<�ܼ�>�<X�0�
=d�<��M<��-=�&��~�^���=����N�932���<�v����;���</�^<�{�<,sS�s�[��y'=���<=F
=V`c=�G<?����x�<�W�:f�����ļ�ik���&=\�=�ڦ<�r=z����Q=�QQ��#���;=�b�<�V�<|�U�<	<=�V<rQ.=7�L�/=<�=�5,��pڼ��8���<�.���� =��<�2��c��t ����s=Q.��\�ށ=W��<K�(���`<~{u<S�;k[k�{}E�c�=��!��p��v�w<�� 4=�E��m. =X�~<m5
:-�^�H�<��3��=J�d=�N`�ژ�<��=<$`=��3V�sqk���<��̼���Z;�)�r=��<_lo�!�X=l�<��9��T��1=�aC��_�<�<�<X�=¾<��"��V�툐<�:<&ʸ<����r߼[X>=?G��.=�����h�*&�;�,���d��2�;a���0D<��A�Ƣɼ��^;�
�<����Y� �<�=/#�m��Ev='t<��֭���6/���z�x=@���Xǖ��F��-=�7=�#{= ���l�<v�!�ﳃ<N�M=H�5�@=5�)<U�=�=�7=v��x4
;h�j=Hj��k=�7���<]����g=�V�:�����H�*�/=h�M<)%$=��û_ǆ<0�E=p�I�!���Е=��<h�t��Ҋ�Dz�5.0���?��=��1��I�ۘ=�[��_Q=�e=���=]]`�lծ<�r��&��1���J�c6Q�����<�4�<��&�p���M��0�`�~=��H�AӔ��w6���������z]*=�=��;��A��+=j�<��<%�>���c=y����A=7j4�H�0�I�
��=j���_��3�@᥼<5������fB==l�dq���T���N=U���34��?C���<E�%=���P�3�	��M������ӷ}���	�܍�<v?\=q�H�{[o=k�༿�N��F���= �Ӽ��L�+�7��AJ�����]�<��߼�e��p�<f\��*�<�8��x2K��]�G�>��5�� �����<v�:Q�A��|];' �;�6n=��;�D�3tV=�=U�[�F�=��< ��<��=h���1NU=�h�<.>�;U�<5;�<.��<��x��o|<2ƍ<��ż��<fc�����Ee�:�a��;�?=$i<��h��F<lE�,�j=M�?P�<>�<���;6M����;��:<;;*�;<���dY<��"=޵�� k�[����H���|<���~���S���Ow<�(=�L{�DW �յ��_ʼ��&�?�|���e�*%=~�(���<��H�o�D=׽�<��3�e�=�*��x%��P�<�����<7�w�t�S=K=���������;��<y!����<q��;̶�<���7�r�t�F���6=^I<_��<X|��f��<���;�������<j�`=��5=���<R�=�1�<��=��=�r���]+<YW�;8J��:>%=��A<1�&=���=�*c�?�m���X��c��
X�<f�+�]�<b�<�&�<���z��65=|y=�B��<��;�-��  �������%<g���+(�^+�����j�����^3<�Z=u�J<j�r��\�\q�� 9=GO��-����K= K=uBj��<��N�K<*�L<�K�<
,���"f�����q�;��&	T=�B3���'=�'�<��=��=aC[=�>!=JSO���?=��-=��= 0k�'�;��<#)�o�$=:�[��D='�G=8ӼT+q<oF�<dK�sof=5�T��x�<|�L=�μȼ�l=H��<#�@d<���Gx�����b7F��J�ۺ"���<����⑻/���s3�
:�6ѼB�=/E=6�H=U��1�<q;p�y�g=?�N��V�c��<�`N=��P=�;1��%e=�Tp��V(�jc�<7B����i���e��eZ�f�~��"Z�x�j�ɼ�pl�2�C��ͻ���º><%�<=R����1�E
�<4�j�%��<���;�V�������fp�}��<�L�������3<i��:��s��X���{=l�Q;𖒽����������=�;�=�.[={M�T������<���� �<�B�eF5�WZ�=�9�����<�.�<JxU���=��t<�O=ۡ�=J�����-�"�<Dˢ<U	j����k==�������='��<V�y=���ƌ�<��==(Ʒ�-�<<�󇼒��֞`=T=�q;�w�<v{;��=�
=q��<J��[�<Oװ;8V@=�W��:�>����<]$j=��<^:����<l)�;4=���c=��*<���;\Q��n��V ��J;e��;��I��c6��4=�^~��0�<�=���<!�<�R;=׸�<�P���=��мO
k��P=C��!�;d!���S»�2=�w�;(�*�&P�=l���?R�=v�Ǽ�0Z�����s�F�6����"E=%�Y��Շ<Kz���z<�&5;��:H����ȟ��T<�|C<��w=AO�<����(���P��Yg4�!��Ͻ����@=�9�<���:X�� �V<���<[b<�D����'=Sr��� =K������<��\=�7�<�|�<J|u<�j<�&�<��l���Z��A;=�i��'=��q���l�Wр�ќ�<��@<m�S=�?�j��<���;v[��=�R=��<\�^�z׻��)��������Q�U�
[=~}b=��D�����Z�X;�%�<�Z��F+�4��pި<	����!=u��9`�<�1�T�c�k@�<և=�|���=�(4=��m9�<���������)=hHH����<��_=���t��;�LN=p�A=da=SQ���i<��7�Xw��~0��{[=�X<*v(=��>��=4o	��`����w=��O=^��<e�<RC=}�>����<�� ��FD����)C�<�O����t�fH�ސ�<m�J="^=)�<<8��*���[0��J/<���<�<��k]�<{��pL�/~�<2v�r�;��e�����&:��+�6<١�<KtE= ��<P��<:L%=��F�.����*g����<م�<�����n� ,3�i3�G�#=<�F�Z�_=,3[=�-/��
=@,<u��<u�=���9�<��׼w���K�<l�໑����t��!�����.U�je	=�� =�&���<��=�+��M&)=���Q}�6]=�W=��k;V�<+�[=�N=:�\=c��<��������<�7�<�~����<+��:�_�<'���F=����G�@<eUu���<��$�}�<jD<������<.�=54�<��=�Q��p���Y��!�S=�y缐�Q=�v���������&��kL�<�餼A[4=A1=p��<��J=���:=S!=�2G���J�q"�<c"=�H�=!:�[�S���mZ�r��1�u�N�;ȶ�<h�I=U��	6^=i7�R)<	�8<a=<�!�<���<�t,=��<��w����8=�{<v*)�WAK�����Yɵ��(=bM����;ї�<��7缓	�;��t���B=�G��@��;O`��Д���=q���G��;��༐��9���;�=S<=u��;��1=��3���Q=��!:��,=Lq,�:��<�7~=�T���o=_ �<�6I=cD=t(<\_�<�!V��Id�I S��SܻZ�]�����;�4O��j=�|+<p�Q�S���VY����Z<�B�<����+���L�|����d�<; �a��̸����<�&=�F[�1�F=�G_��M��G=ޛI�^�j=��׼�Ɵ=Lz���T���导�.$�u <�c:2	ļ8E�9�<=	9=ѿ�Bzr��4=[�-<������T<.�.��Z=<��</��=N���@m1���@=X`��1=�(�t���O������ɒP�bw=:��,d�s啼D>X��-ü׹��ȸv�`T��0�^=XU=�f�{)�;Y7̼�l��`E)<�5�<@�2��1;��ʼK���Vo�Dd��JK='�<n��5�X�v}����<sD��ڧ=��O�#�<~G�<��=SP=H���=8�7��=�ɡ��0=y��8���n=�0��;=��b���<�Q,=�`h�6�I<�{��)��:��<� �b�<���cm =)��;�|�:�Y=�Q'=C
= �g=�"�<���1P=M�����;�$�����c$=]��*VR��^[=(l���s����)��4�����
O��C���<�@<h$=���e�<@9O=$�ͻ>sS<N�2�SM�<�=a8�Xt*=?=�~�;���<��;p��<��=Ϊ!��/���ƼRR=9�����<T���<�9���$;�1�<R��<�KW=��D=���<�U=]̭<ޕ�-©��꘺�&F=�����H <[w���<�!!=ٷF<ăҼF�=϶M�Q�<�Ǐ�B2=�;�Η<���H[Q��I=���<�PI;�M*=�%=�%�;��;E��R�<a
<�F?=3�<
,4=�h	�a{<X0��R{�jƼY5��f5�<�#�<M�2�	�༘Y8�qF��oM��κ�����x<���<��7���F�I�<��	�����_0<񗵼��𼐆3=?m ��9��Ak ��2�<�Vs������W�z��<�̀<�=/�<S,�H���A& �_a=9^�L�c=Gc��5�����cWG��}޼�+Y��;�lD�Cƞ<��"=��Y=S�yF�<zU��x'�<��==���<�(2�?�.<����:=\�V=�@�<���I�;��.I�����=O�ެ=���4����u���H=��z=�9<�]���h=ݙ=���-=Ms�<�.=���<�Z=���X�2�&6����z��P=2�8��E/�l��<G5k���!<n�V��>K<CF�hq=ȉ;=��*�=r<ǉ��$<�T���+�<�+��,=��<��K=ۏh���<�d=0�=D�X=ؾ�m��q���R��O��?�@��'=�7=񙼚_һYu=.�<����P2�K5�<����b�2j=O����e�<ˡ<�'3�O��<Ί��»��=��W�y�'=��;N��<��Z<�U=5�<"M�Ք=</�>=7X��H_A�M�� ���3�����*#=�k��=u<`-O=�.���hs��g��A�D=��K=@*>�q�P�D���
V={�R<*� =�i;X�T=��^<
��<w3=��T=�x�o��<n]=]M�<�U�<��^=5�j� =MnѼ��<Q�8=��2=&�8=e�-�����C��8\=C:�&ʐ���N=\<��<�f&=y�3�@n<NЉ;�$������v
8=տH=��<���<;�ݼ�����.=���N��lOG��cG�� ,�' m;��F���@�d�0=B?�<U���y(<J�3=��M��y=et��5=�W�0=w��&�}��Ւ���;<��<@�E�,+-��܊��D4<F�9<	��<+M�:�c�� ���R��U)�^�Z�z�b=,pٻL�-=^�=ُ�<��\�⢯�w&���<��.<�j��d �$��=�ϼ,�Z=t@���d���!��b<�=�<T��<�������)�6�Zt0:��V=�C=��I��-=H*��l=s<~藼`�"��
<U�<�-��O�h8�����b���V!=�4<�K3=����ļmc6;#�u="��<�#_=w����Q=��1=�J:�6ܼ��o<����V�����4=���x�$����<��k�K|�<+��a��<hj����I���)=j��<��@�0��<@R�:h�'=�=P��:N��<l��<��1<��L=�<�:��	�!�r4#;�ZE�q��:�=q�����<�W=I'<��P<�=��F=Wi��sW�~��<����z<��<{�1�hL��i�U=5p<�-=3m����;6�<=�#���/��|=P*<��<�a<�y6�F?n�&Uʼ�ڀ����s�;�>�3s�'�+=��e=4߀<��R={�A�W�Iv?=�p��J��L�;i-��a?���4=���H�!=��=���;�5V=�H�<{�G�t����˼9���A�<�����6�@�#���6=**���ɼ.�D=f����@-<�����U<H0D��.=V����<���<e�ټ��V=�Eb�Q���[��<�;=*����/=�2 ����ݴļ�a;.B=N�:�[�<�K�<�u�eɠ�]j<���y��9�E=xl=��8��<9O$=m3�<�*��|�Q���n=�}^;k�=D�=�ņ�
eG=tn=:�C=@�l��<�	=&�;�k�=��=�9�=��Ҽ/���伸 [��X�<v-�<`�,���<�a=�(3=\=l�޻6��;ퟜ��u'=�_5=�=�,��J:,=��A�!lJ��3P=O 2���M����ddS�9`�<�,"=��һ}��}t�;��y��=𨁼�Թ�Wz�s`P���-=�q�-�S���4��<�"�<H�&��Fd=9OK=7X=LS�<`��<�v=@
�<�Lx;T'�T��<W=��\=�E=���<B����"/�������d0�֎��Z��{�2��M;������<1�=�e=�� =��I=�]:=I�+�;�s<%�uk �1����n�9%<H�ּ�T�<nN�;\�;>����-�<q�!�-N�<��%=[`=��:�b)��9E<ݴ=����t�=������;���v�xi,=
�<Ι��v�= Π=�ۻr��K��|��<m�ɠ�<�y��fX���+B�"��Ne=^䥼��Y���t4=D�мm�����\
�<�u�<���Y2�!`_=2w�:��U;�����(����r�W=����e@=�8K�C����=��N�Kcn�F���)=9�#=GW�<��C=��<��@=�P\�Z0<����d�q=��f�WV�B���Ǽ�<M��D2=��<犮���B=�t~����:�d�����b<��~t	�6b��������;X��<{�<ms)=�A��S=�(Ҽ���<�oO�9�̼Y,�<�=��g�#� <0�r=O�<��Q�`�<�5�<ޑ^�g�=�Mֻ_sr��.��a=�ϻ^��B�<@Ȇ<�/�]ꀽ��J=�F<L�ȼ�4��Ǎ��9�?�6=��I����=��5���8�8�R��~=���<vI��8�3������"���H1�M�(=�PD�kb=M��d�.;^T�� �0=9>=���<.�9����uZ��ё�;�=_4�FIl<�EX=$dR=��ϼD`	��T����<i��<q=lG�<>�q���N=yCL=*yE;[C���z����Dl�<�\��8eE��~N=Óc���=d���b'��&��<]
=}�"�[�ﺖ*�����-�E=�ܼ�}%�ㅜ�rB< ��j+E=]�1=��T=q/=��B� q\<��^��$�z�dx�8�r==�>�)�<�a�&�]=��(=L���
�����<u&=�%��=L�� Y;�k^��M���?���1<0���U���	-(<|K=�B�<�[�<�D<��;��<��<�qU�a�<�Rݼ�3���5� `�p�	=_E;I��zrW�l�����<4�x�3��#��;�H�����<�yb8R:y=xB㼡s��Z�ڹ;=u�7=n�&<Psa��(=g�O��?<�0=}��<�D��:|�;�B�<w1�;���<ٲr<X�S�J���� Zy���<@_����&=�@�<�����/2=�n�<��!��������ɵn=gq���=�hQ��j=N��<�UX=y�=p��<�<��;��E �J����<�ok��g�*�*�9�)��ԼI��=��;����$�r�S�<�B�r�;ub��9�	�d���a�<T�EV�/��p*K�;��=	�!=!���Nh^���<҈B���9<�b�.=E���:�C��t��%�<1 =H8R=.�=t27;Y�v�CM�����.��$������<T5��x`�<��/=�==�;���Bļ4Q�<��=e�<.�d=������c=[�*�H��<��<Z�%������<�w����:����A� �*����[�;�� �̫ �k�;~� �M=��t0<�<�<��G��u��0d=!=<��A=P�;��=V��BO�;��	=)<!-�=C*7�Q�y<z"����B�iC������^5��N��)-����;ͮ=a�ǻ��=71Q��~:iNj;��w���T������<��w��(׸�C<6GW�U�G;�v�<�IJ<Im=K��E�<>h�����=��t���_�Z�����*��r�e;��*����:���<�j�U=���9~/
��_�R�<�����Z�<�d;��:�W�%=e\�<����\$=�r��5=�i����;�n��_�<=t8v���6
8�^i=�~c�&=����nq�9|<@$�6x��d�;���<�h�<�G�:���<�<�<=��w=��4H�d%�;�9�<Po<�D=A��<��.=-\�;\2	�˔;���ۼ��4=!�@=>fi�.>��Zļ
Fh�o==��=��Q=�g�J���cF����"�:;��z�@�9*	=ʤ<�Ϋ�>H�;WZ�:z�b|:�%�}��C)=~��J��ĺ:n��<�'�<�,�����7�n>�G�`��4�<N��<h�!�͹�<�ª<.`��x<�A��K�=�㐽bU=��g��-3�Ml
����<N9ռ{�E��ٞ�������=G�)=v�C�
UE=[�c<�G;=G6=�?=��*��M=܄���j=��=<�AP��F�=�uм��=m��J`�52�M��9Y�<QD�2����F�=LD������UfX=�( ��|,�3�=Z�>�+\��h��E�=?f�<����X�r;b��$Q�Lf�'�ӻ� (�6{Z;�jS�P�g�Ұ��X+Q=��b��$<�ά�Ppj��S�9}�S=�&��XA=�^=��ܼb�� �%=��k<d�b������g��{�2�fCA=���&�<�(����<�j;�Nb =5꼊�:�#�|��ٜ��@�<<���d��M��z��� =�k�"9м��+=�;�q	����1�=yr=ѷ<��[����Kj0=Q�"��
\=�1=�_]=IX,�����Ei�eܾ��9=��[&P���l:Br=��\;^�O=1lY��4z�7�/����.��!;�b���y�<z�2,��w�?������#C�����=�#���2�l�	��c=���<�3����/M(=�6;�dR���<F��=vcF=V�=�T�<�����Jc�O�ڼ�~(��@�w7��mN�M�<���<�#k�p<=0�D=��~�ם4=�!=2�h<D�5�$�;�ƻ�Z���U=��^=(�B�;2;<�<��{Լ�==�	)�䲈<< <��V=��b�r��;M�=����ż����<{*����=X�+�a�I<]�m=�E�;*��<	�{��Z%��.=��N�����<������<�{q=ļ"�#�ė��.B����<+���<�C5=/V=�v���Xm=ĭ>��L=�<�j<����k߼�L=�C_<���:��4�
�L=�A=��<@h=�;����< �
����J=2x�/�X=N�%��~�<H�H=C(d��`=>�
�Z��<�su=��(� ��<ؤ;�1���T=.�h=z_'��U���<l���;����.3�;��B�L<��û��ݻE��<���K=��*�O�B��K?=T��<�\}<�=�]V=Mz޻����55V=�+����7<-�i=�2�ʤd���ּL�<6ZлƓ�<h�;>z�k;R=�?����=$�<�S<�B,��V-���F=�U�<��,<c��=��˺�t ����AX=�2�<�?I���"<*�<e�(=��h���U =1�:�GS�����L�=�t��O=y��M{��~e=��Ѽ,�:=�\�z�6�ŝ3=��<�5�;��<���<� `=�#�5��<x'=f�<�μ��V<�D�Âf��5X;�j�`��7����=�di�{=z�<A[	=�@�<5T���=�(N<�.v��,4����<�2=��*;�<q�)=�d=���<&�1����
<��p�>�<�]��K&�[�,=�R�<=f���@�<蕧<��D=�	<YH�������G��9㻃�D<ۢ�<�Cɼ�A&=m_�$��\��<_N=���z�X=�Q<���"�"=`�@�=�F=��z�C��<-��<�i�<��6���u�Pٷ�즎���H�_?��P �p\�<e�<��B��UJ=T�\=��[�ԝ1=پ�<�h����Z4��}?�qh	=L=�<�J2=�N�Tݚ<S�I=��T�-�=�0��^��|�b"�g6O='�Q=�/���S=�<wl�<�4�<HB�<�3�<ʢ ��e$=a��<��>�&�(�|�=�Y���s!�Q�h=�A�<c�=��`=á��d��k=��9�h��I�<6z#�.��<�AA:O0T�]/�N�E�����YW����+�&�/=��	=B�м�`w=��<�<"=�7���<����h�<]᲼��&���I=����S2��� =s�5=D+��ż��X=�������}��I�I�<�ͻR6༲�b=zhm=�WJ<RhJ=e)��B+�0�=�xO�Ѕ���%==�<O�Q=Rw�`�W��_��I����<�0�%�;t�m;_�m�eF�*��<�e�<��S=�^��%o=V�;_�J=�J{�m�Ѽē������ ��%3=�O={�G=�J��'��<�F�jHK=�ͺ<��V�xH߼�1<=lZ�:ϨW<�&6��&����=U�-��_���<��<G_=��	=��ϼﻴ�=��<�p<����Q�@���a��u�m=T=A|j�P\غ�Ke���<�H�<�_6<RG%<�u�Bɼ8���Y=��<�?=5��<���<��^=;M�7�6��>#=����<�<���< �1��;i{U<c�x��PL= s=����<���%ڼg�� i�b�8�'~�<�o��;����;���<��컈�<R$7=&5�<js0���==j��<�{�=�#=YU�=�2��z�
�-}�={�@=�0�:�-b=@m�<��=�Y8����?:��G=��(�����-�w<md�<�֥<j== =�e�=!��<^��:Z�W==|��N��<�M�S#�<4蘼-��<U� ��3��.5�=�m�#0��Z�<�s�<��=��p=�J��wU=��.��	��Uύ9�&�����A(=T�ڻk��s�K�/��#=������e����_��;��<$I���{���Ƽ#4ü<lX�����l=_��<�8��_�T=�c�<*^=10z��=dv�<dK��"=�Ms<g�D������'=�V<�x=��TI��}��]6Ҽ٤Ǽ� `� ?�~=:��;X<�=��=˰<��?��(�<���<�I�;��<Q��;wE*���>�t�@�}�Y���"��r��7=��6���E=?u�;= �o��;&�^����;p��z2�s�<�
k�(r\���;VN�:�G��~��=Y��<�D���V�D��<bq=��:��=������<=+$�<c�F=���<�����S�y���r]Z<T�h=�\I�4={p$=�{���L�%���0'=�f���0�R��<�:�<���vHC��H����`��	��l7��h�r�x�K<�i�$,M=�g=�뉼�mW�A���P45��?�A�_<M�ϓ=<��"�(k̻��<�"A�;�K���"�~�=�]\=ݪ;��mż�,%<N��<�R�#�����һ����(��$^��G1��d�<�/���`�"�,=�=㍳;ϸ/��~R=�(`<����=�{<� �#*=*�`=�� �I�=WF��B=�� =� R�ܹ��g=x�z�ܺ�<�)����<
Z�
i�<�'�c�M=�?
��VE�K.�(�8����<�V��I/��c<Ov*=��f=A�Լ��к�����1�<1�=�ɋ<!T<ݡ<�Q~��8�<�<��N�s�fzŻ�Ȃ�,)4��6=E��<�e�-J=%�;YF��p��<Suf��=o�1=}��$��/�<��]=pof�Q�,���#<�B�ʑ�;�w��4���5ׯ���=�:=�ܼn_(=�T��_==Ґ�<��5=Vn�����;`q޻e���c��6;�Q@<Bv����<�Z�:� �<�}=bFB���K��b��<���\�<c-�<��<�s<�<?��<�����9<�[�<I{���f=-��<�"=6�=����<�Ӽa)��8:=lہ�#�v=�J	;BP�;�P�;"�v���V��=9=jOX=��=�>�<��#=�#=��x=��5�lK3=��<��V=Ki�����</�"=�vg=���<ϰ����,�����(F=oP<���;�|麂VO���<��޼%�Q=�u<��J=�!z��#=��T<*M=�l!=�H;4=%��<m��<!d3=��~=Ev��F_=���:H�$�ո<	-�:άF;�G���������<��f�b��Ď�ԑ	�H=&�>=��<�����<��iN�;��	���V=2��oN��1=��=*�<���H=S�C=��=k�¼d(=�T���VY=��y�D�q�@��<d�I<�B<��>=�?K=ۮg<�.�;\���2;V�;��������<������z<���<��E;�!�s&h��V���=�S�<�A��f��~�;?I�<���*=FU`�O��<�q�4;�;�`�<R;=� =l;=�6C�>r5=Ɏ�t�9<h8=�/�Ѵ5����<����9=�Uk�u�S�k�N=���9��<K�<5��u=*��;þ�<��0=&1�<Dg��������;�}<�F�:�Y_=b�P��-��o�<t^=�đ��&�<�7�kһ���<��ͼ����m�=C.<J�'<�O�<��<�/���`��̼/O:=��z<_?����<��;�i+=�Ӽ3�[=���z�:�@�<��<����u�<%��������a��C�P�9;N�<���<�_V<�@�<���:{��j�;g�G��?<-
�<
*��],�%��;�����=�/^=���%�/)=�=�1��@�gF�<$y���K���9!=%B�;�-
=R�����I��ZG��7���=����=)�"�xPG=}��L�="=E�9=��Z<ւ�<�%<Q����B������<�Z��m=S�����̼!�n���'<J/#<PyB��'=(4��,==fH<��<ep��6�"��=�Y��5=c�E=�N���ǁ<�4w=�(C�E3�F,���$@=�6J;ض-<t{�;o{��D��G�j�����<��f�}Ƙ<�����Qy=KY��m������s�%��;��U��Y���%I=��%=�����p�`j༻�>�E��<�{	=fBм�0D=S��<���(By�u��/`�&Ѻ��@kE��+�9� ��
c��#=�E�9�T=��); ^ =�ڗ���|��=1-F�`�/=x��</(;=�v1=��v��ed=iU@��G�Ƒ���+�Su�<V5<�V�=�Q��=I��<i�O=t��<��n=�qݻ�
�;�Y=E�=�y	=�ۋ<d�X�v�t���=�]m��E �J�=�/�sS���y"�9#���<�@��K�g=�GJ= �F��=�´��f��^=YX���������N�D�^�=��C<.yJ=���<���;�
�L䃼鋃�3!\�.�8=b�4<:�:�߯[�u&<Fܖ��sS<P
<��<~t]�m>̼X{�;�m�<m����F�=Jg=Q�[�I�<d�O=]���f3���u<L��^�<�s�<k�<�eH�����������<m�<PT�<~:M=Pk=���Pw߼�؀<k���=M�<t���O�;�?=k��;�Ư<��b��u=x�a;BF�<�{)=ߪh=g�	<�BD�|�<P�#=��<ȡ0=�D���=�3i��=&���ӭY��%�<���G[�ρ�;U1=�jټյw;�i<}/�<D�
=e�];I$r<� !=1]���ߺڼ��<��==E�N=.=L�!��y�ke�;L�<r83=Ph=V*Լ��y��#��W=Ɓ<Jh�;�]~��ؼ�4�$j�<��鼢�Q<���:ϸĻ�����B=b:8<�Rn<U��Q��A�;�2�<um�<�.��=�)���*ea��A��Qo�+�Y�)e^��A�<�h
�&<�ۻy�k�=�˼�ځ=�[�<�at=#�2/��^����n=ȕ?=�q���`=���<��F���	�}'���;v/Y��6=2�S�~�=�����;=&c�X�uɄ=L�*����:�,��aC=�Y����Y����Q�(�V���A;<���<�-==
Ǽ��
�<�Լ�`޺8�<�B��n8`�hA��<h�:Z=�
T=�"��;�=T��<��+=G��;�8=k���6輕�/=��(<���<�o:=�W��^Ow���׼��N=�P����n�]�ֻ[@��=��N���J,<����#G��T<='�~<��{����<�_�<�Y��V��;M|�<\Q�<Kn=`Y'=�6n<��(=!h*�8����Y=A�:�M��;��f<����<.}�;Rʡ�*3׼g�H=�/=F|�<��J!{��=![(��[<�>��"Z<W=6�<�
=N2=���<%�U=^�q=7�Q�o�׼�D�<�.=��D<9r)��&��:n�}m<�#\�K�<�/�T�΢��Ab=��"=2��<h�.���=ks]�w�(<h[��F���wC=n���AH=�,P<"�ʼH�;��a�G=��a=���{�<�6i�����]v=�"��ag��<����`D�2�$�+k����0��x�<�를9h���P0��X̼�x];�ct�oB=o[;vz�<H��cw;<�M^=�L:��<�<�.=�^3=&Mv<�<�<���:�8����1�6�'<<Pb<j�<{p���8�X<�"4��E�;��M=7�r�ٓ��CU2=k)=b��<eD'�]P���=�u�<!���:�6=������Լ̦�L9��t=�$G��I����U=�W��{g=Hh��47?=�=+�Ɍ#��X<�Z&=O�Q<F�;��0=��b��<("<���<#��twY=R����E�&u������rǼ|�<�2=Rdq���;N�<��=u5�:����Y�Ƽ��X���&��٘;�|�;�*�;h��-�׻�B�V��6���6J���1�}�;8�E=v�H�>�R��z2���<��S=���<��N��l=�+� �a/Y��|p�ݍ[�N��_�<��<��<��[=��4=�͝<4���K":��.=_�@��D&=�v?=00==]���{���;�;���h�g>=-]�<C��4 �nV<���jp��1�<B=N�<kX�<"�=۸�<004=�Pd<��'=�I&=��<��M<�?K�ڝQ=���8��"=�=fZ<�O�,<"W"<�*����l��CE���<5�3���I=̳s���;]�=�pl��	������w�I: =��3=��<�j�̹�<`5�a��m�<V��<$R�z�A��5�<-�<9�+=&�<<�`�VRd�y�Y�ģ=q�<<�a=,ȹ<@~�<�#)=J�����<�x ��S޼"��<Ҭ!���@=(;=�+�=�@=��߼���<���<�|���D;=_�(��["�XU�<�ǅ<H��<(o9��=��@=Sδ<�
�<�����K���_��U|<r<;�R=W�.="�+��f�]�¼{��;�;�T(<��=��<�~N=>	��|��<���<+�S=Cc�<�ڻ�.���I�!��<�=�6=l�= ������"�����_=NK`=�S ���=>��<8�+=s}��h�=�x�;	~ȼ��O=�C=d�D=��8=eA��<�d<���<g�<��^=��X�~��f���K$��U5��¥<TQ���-�P���]���,�<���;O��M�2=L�;<�ûɽ<D6�;Y8�l�K=�"/�$��������}S={2=�Q����u)����<΁�����<���S=]=�i�=�)�FH�;���;�Qv�ka;<U+��8�<�	H��Y��>�\<X<r=)�5=��_��\=��H�#x�<����%¼���<%�W�DW��XG����=�I���9D=YR=@��<S�=��;��O�o)=S�*�憆���;�6O=�r=��<��D���R�8u�<��;=�D�<���<�����<\�/�m�;Ig=AUE�}x<��]=��<q5u�����)�<�ؑ<Q�� �i�R� �:-0=*=Ȯ�Oe�<�������C�~��S�#�!���<�F�<�
(=��g��^>�m�ż<Ő��qѼ����=b�u<Rs�V����;�<����.G=�*�=O2=0i�<�<��2��=%�
=;hB��v�<W�b=�=� A=S�$=�i[�y,����+�K�w�e�b��(��=�O�X�����h|���L=̗'�y�>=��;y�u=�亦�=�h���p�h��0=7���<�<S=,�=�o<t$�;�1b�S_�!8Y=Et�^�F��d6<A���=�*=�UH��$@������<��׻q�=]rH9��>={��<p'�;ԅX<�o̼�1�C�Q=��<Aj��(8�<Y�����M=��:XF�6M?=b;K���<r�=��W<���;�e��%
=�j��2'X�	d�<�{"��Z����}F=�e���O=MՓ��0�<�&=�@�<(�+��&���b����<�V.�z��<r�@=����n���F�A��t�W��:.,8��;ɼkE����;^ <�YZ= ]o�Ҁ�=@��<&�;#h׼��`��$�I��X��Ջ�<�������x�<�l�;��=�&K��O�;z�e="As���)��<%S<Ar==�!x=�<�0@=N(==3�~�]� <
���h=k*=��A�oF�<�����M�=j�:(y=!s����ҼV����O�<j����2��#5�4(n:v��^�G=��1=�<�<�O�<Y�û�06����9l
r�P5h< �u�=d�ȼ�r�;$#"=et���!=���;I��;���ԋ�<�>=�I�<&�=2�=�~=��޼{��<*�P<v����0��`��L�P=����<s#���B=����N�y�K�a=_�=6��<ZC�<`�j:��}���P���?=��1=�v��n���,<��¼��P3a�;�Y��gݻ'�>�]+*=_���=�H�� ��jE;^�q<��<�p�<��i<܊<��y��,�;3�к`FD�۰)�!'�<���z�N�$M�<  2=�TB���M<��%���Y=���j���"�)���f��W ��9=w�:c�!�,;ީj=�~(=�L�������=�{P���=��N��j���=�j�<��~<B�=��=��?=��H=-ޛ�x�|�@���R9��I��0��ҍ����]��y����R<o6<�C&�����<*9=��<	��<`�4���Ȼ��8�.6������xi���;!�[1�<��=��<Zp��$�=E�|<�8���ɻ��̼d�º�^�m�c;���<kP='�Q�
�5;�<p�N=	6=D���� =�#[��)3�x�=.KS�`_==�C�<d��=��<�"J<B9:��<jf==�B="�P= @��I����==��J�Jy����ɻ�w�<4K�}�C<0=��xFf���W��F��9�T�Ok�<�� =[Ė���="l<{5���s=Y��Z�#����K���-S�hs=�E�<�Gi��h=�TW��l�;��ɼ�ڴ���7���*=���傱��D�����B��;O�X�=�4�<�sK�k�/�=$(2=��Q=agN��s<sR�<6�:�ʫ�<�#(��H��>Q<�p� &M=�g]�ܻ�R=��Vd���|= o�<$�;����Ƽ[n;�N=�NP�f�<�1U��b�;����'�%�b�����h����"9=~�e�RRe=����<�"=����@޻�B�EU�<�^=�b껦�:�C=&�d�3����_=�I�<�j=e/�;7�G����yջ]B�<��;=�>�<D�#�&�B���h��_"=I�ɨ�<����n��:�K*�@w�����;�'�<e�ϼ�a�r���I�;.ز<�D�OI5�%a9;xc�
L;��(�$��<�>�<�����}�Z^�H3=BbQ���4��_�S ��%E=Y+�<��7=�q%=�)R�)�;�<��%�=UF�;w8������j��0=��/=�L9*'�<y���gE�\��	�5=Q�E���G���<�@<(N=�l���D���h��'R����:�=m�?���?�Db
�}��a��������Z=��0��GA<�i����EI=l��<����.=Y�H='�=Ӥ1�o0�<��<��7/^=�1+=�ؒ<8 E��E:=�6e��K2=�H(��['�1#�<��<��;oO�<m��<SY�<P��-=E'��s x<�}����@���K=�]G=ש�<D�<U�p=Lk��s�<�o=���;�>=|�=������a�s �T�N����< b=������k=������<�#��y����n8=�޻�,K��wF�p�ڻ>��� �Bc���=�=g����;�Ƽe�3<�f�S���#���:=Kg=b#�0h���,�j���u�7
<�<�2o;�
%��!��u�<��6=����\D=p�-=��;0'=.�7=w$=�_���=/'d<Ev�<�LP=����0h=%��z:&�Bt=�P<�r���)�<0i�<ƄO���'=�T<�＝�2�@�e=�X=O�:<�t}<埍��{R��r~�V����x��N=E���d=��c=Wv���<�t�;3�#��)^=��@�[����=��M=v�E��[��U,f;w�=����<{:=��k�i<m�<=��<\���'�u�F���˼��L�{�$�Q/Y=ߺY�tIo<�6����<�OL=����K;�-=�9?��=�B=`1U=�IQ�~;�<���V���|��l;��G���#���<L'��/¼��-�o� =ghF=��9���-=5�#� ���B3=�4Ļzy�1�<6L���=@����
&���2����<='X=y5=�����24=��u=�a�;u�������1<���<z���M��R=��_��5��?�|;�!<��<hS�<�~�؛��vf�?�Ƽ�_=�Gn;�v'<ʪ�;�;���<�`�Zg���=j��<�H�q�<�:U=d�H 	<���d���H8=��B=k'=���<�36� <�\�<+��<@X3��o�;J-滓� ;~�J=,	�} ��[��^K��8�򼙕"=�c��?�i�<�q�<[���o�.�=J���s�=��ڼ%?=��
=��<)6��h?<Nb�V0h�]���N=��+=�N����;��(={�E<K��[��<w�D=����z||<��$=#���V�����<���<�R��L�-<��6=��μ�<x�<<�����倽
��:<�p�VZ=�����������9۔W����<J�_:r��<_Ln��I=(B�;.=U1�=!�7=i�Q+n�ŀ�<ltK=rD5<��%=�*'�)�-=��s=�=�h=9y=��0�e�M;@D=mĕ���4=��6:Ր-���|��F�:�.&�˅�<��D=hx'�������=�Y<"�=��`<�����=�����F=4�^�1=������<��<��5��	��?B��b�\�J��h=(�;��0�H����=�<C���Y=�.=�y�<��,=���<�&�<d��<�$�<�ּC�D=���<�O=��͹�IB�yw�<ܗ���\���t;��Y=��<���K,�<�@�5�a�*=Ц]���Q��[=R�
��_8��(㼪� p�f�=�G�<��V<�x=Gs��+�a�c���A=�]���!��%=� u�pm=�k�<W	e=��ѼJ�?���%={���C̼�����<G|�ɤ=@�O�����=<9<z8F=G;�Y��;��d�qH����W/̼�!=�O�@��<_��7�	=0���O*=.&<�@L�FN=T^,<H��:*m.=�Ŷ<L]3<�}=��Լ��<,��<-�6��과��2��:��Ӽ��V=�go�j�<(�[��
;=��<f_ּK⻼�]=@=�悼d�,��N=\f�[����9Z<�<��<օ|�9��9-2����U�#�Py�1��U�eT=U�;a}?=���Ӭ!<+����M=�\^�fkO��0!=���<��t<B �<�r<��<�������<F�!ͼZ�ټAie��F���l����<:���Y�'�[��~ܼ�����	����<��?<�l=٤�<H���I���z�>���X�w� ��"=�]='٥��V#�j^�:�m�:�p�fW!��ML= X�_�	�lg=72=R�;���;
Fd�4�w����<vP���2<�M�|)W����"��<]�;7@�L�;-�M�R=9�E=��1���2=3�X��>F=�k���7��/=�<5~¼�᰻���9���=C�UQ<=ˎ�<^�:��<,. <ng�<m�`�(�;��g�
��/=�2�N�I�ɼ3�u�6v�:7v�<?]B=��<2���|?�2NƼѭa���ܼ��8��[%='S¼|B=�4=@Gd9ą<�v"=�e�<:���s�7<�J�<�lG<z�<�P�<D���J�<1V%=�q��o[�<����[=~C�<7�=��ּ�������J�%o=&�i�-�v��9�����];ʬ��y�<���<X�i�g}<�&���6=�e
��>#=���<p�J�+wӼ��O��T����,=L�`�=��:U��W㷼31R�c�3<Z�;ÏP=����T(���Q��CW=w���g�<���=l�C�{�G=+VE���U��3S=��d��]M=���<)�a;���J�>���=ј��з�<�a�J���4����^�����A��hk�i��7�6W=�@=��=�|��׾�<��';ķm�A�I^ümT�4��<��/��'�JON�-�G=��B�`����E�<<�K)����;�E'�x��a��<�M���*=͓_<���:}�)��<������X�A4�<ӊ<���iA�s}<�,>=�JZ;�[�~�6<2�����b��Rj���X�%�;�SL<�3ȼo=�_"�ֶ8=�8��G3� �<d�=�'���F=S/<�$F��@-=0��<a�<��%=B�;��6�(��6X�;�h=zwg=R��q8=9���{;2�5=U�>�w�����K����<��<>��h�e���C�Tm���:=ڦ=��<݃�PT弹h�<I�G=�?Ҽ#0s=jTi���P��o�<р=�5e=}����:��yT�̺�<s�H��PV;m�[�~=y<�<G��<�9=<�|K=k��=�<�����I�"�=;��<�\<ե�<I�c=r�`;7�����<�&Z��&C���M<W񁽷�:NM4��>��1OS��a+��K����<�6˼S�'�B&0��1W��2p_��)Q�'3�<n=��'�k���"�D
�;z@ļ�=��`=�M����:��=1h=�)��ED���<=3��@�d��;PE�S�=��y�@=��Y��M<��=�1E==y<*�=ɠ"=҉�<�M:=˧��I�$=r^��O3�==x�u���=��(�81(;�:�<�;/=�=t�$�lt�*֔<(=+�\=�d�<�m�9�I�'�5=�/���s=G#���<�7������~�> �:�W�̶�<d�!�rdG;=}G�|����1��
�m=�N�<�:=_q=y$ =������=0�QI
=�ى���<�j<�L�W~�1$a�o  =�⠼ҶO=QX=�;=�棺�u�:��h������S=�� <8X��qO=�ڦ��@���a�>�ʸ^�<���<�-��O�<"f�<���}�����=<,!���,B=U,=W�:=�Y@�Ѷʼ��^���<�R�<
~ۼ(��<��<���<^Oq;_�;$吼8F=;�9����97�V,=��<�x��Ͳ<��<i�z#=�ؼl@=�����h����<p=�=P���3r���H���]��Ms=B�=~8= "�<��<�~X�<Ҭ�|�)�s�<VP/=���<� C��n���>��㍼��t<{M��s�+�ĺ��!;�R�;	ɼ���< �<�ه;JI��� �3o��6��`<w?#;�� ��؀�D�;�4[�o�<E@����6<�'t=R
2<�9������<��=_z�9$w��"�=��<�G4�����Y�h�O�D�D�+���V=������<��<���;����K[6=�z��;��!��ޕe�|�;Mo=�2=	=�ݼy=��<=���<+dm=K�J=���<�>=v� ��~�;.`(=���V�E��<�}�Ǽ<0J=��h�C߸���<�X=�馻��<0<�Ì<�<��D��m=����;�甽���< D����<BR�AB3<r����]=�����:SQ�����m�<\i�<�(=���������=����;���+=R��;�q�=3���G=K#5�!�*H$����C)=�\=uF���ż�ͼ��<����׼m��������;z�Zr=m(=
	.=��s<k缁c=�{Y�%�7=��<;���D*�������B�(�
�a���<�)<ׯk���:3.;��Qo��I;7&=O[��Ќ;��J=t3<<.����;=�ٚ;�VF=���O��P9:�j=�t���[���)=ή�GG��1�����}��<��y=��<v{<r���3<��㚽�? �V�<�]��<�>(���㼑
B=ΐ==TN<�}ۻQh�]��<�	�#�<n^��aѼ�x)<��U<��;�f�<�K7�(ڂ=%�<[��<�$��#��<���;Z�x<6zm=�?Ｓ��qφ�f<9;�<y�g��������|�i �/���_�<�j%��#�<ёr=愵��#伭߼���<�A�;�,�Q�_�3蟼|j1��8ں��ܡؼC��<�a���Db��Cp=��z<w�<��<D�=��:J�1��˹<�.<=��`8:]���׈<�=�^�<��μ���s��<�X=�N/����<L��;G=f�i�|~�	H�e'=�ez=�)=�xB�;��<� =8�!=U�����<�
=8	=%�*���A�Yxh����@=x�Z��y*�,�<��F�Ex�:0�<VuP=��¾�+C	<r�r��<Z0`�L��`ּA|;�3=&�<s{�S��%��;����=Y��<:S���<�OW<|�{=[Q�<�P�Êy=��*��=��q���=��2��ܺty<�o�}=�����S��]��^��7;#=�
=\�C<_K�����'#=1t(=rM=��=$[X��)ڻ�V'����=�誼�f��"¼�2�<�N=�lg��j=���<�]���<4�	���=	�=b C=
-=�?[� >�<5;: )���&�S,��du=����F(e=g�4=�!=��/=Dc�<�|��P�2a �V�a=���(<w�����:����.�<ڼQSH�Ί�<�P2�p&=b�s=d=�.T��gF�>���}�;B F�tv;��d=��a�:t=<�}!��G�א���:<gT=�)G=�ɼ�5��ͼ	b<���;#�u7�ռ�?[;)�j���;�K&�{PA=Ɗ;���K��<�����9��k���;8.�<���;7�=�׻E=��\=J�j=��)�K���ݰ���(��=��ѻxH=�	=X$�|#7;w�%��E�<Sڦ�Z��<��0���H���U=U�2����<��.��oN�}�2d�<[T�;|�<3΁="��>��;����K2л�=g�������:��;Clػ�o<�R�<��/�|sz�A�c5��G�<�\��r�:M�<���-�$��=x؆;�=�m <{mڻ���<��y������G=۠?��IY=�5<c{S;i5�<�7���w� ĝ8��d=�T�E!=�JW�L�=#�\�$�<��$��_*���=ja��S�H=p��p�=&�Y=��;���<���,xE��H��		�����cܼ\�%=߄%=K�=W�T=Y�E;ݜ��BI���[��N����E=��=Ȝ��Ѿ�<��G<����vܼ%��8�<�S!�UB �0��U���(�=�[�=�ほ�:Y=V��<��<��5N=�X;��s<D$�<�V>��N/=vw鼁Y�<FԱ<7�f�'���$�:�Bc�H���f�G�<��L�	���8�е6<�:�<�);�����<�^�9cD�d����UM�l����2��D��<��,=���<�辻�d��h{������5���W<�~����<5^��h�w<�t$��M=+;8�7:=/F4<�z�<(�<d�7��E�<�)�</��<�d�<�p=-#<C�˼y���Wq<�H���=̌�<�X=�X�.rH�RlW���7��K,=�hw�S3����:�5��#y-=��#�G���6�����c�;5#h;�v=�$%�Cu�<^:=���<.�<�2�<	I�=o�;<�<b\=�"=�c;CUO=ES׼�L-��-=��F�W�%=[|U=L��,Q=X��=��<�!����ޭ<L��7"�ά���=��R���M=e6��0=�s�<�����<��:����|��c�c=~\�H����t�<��=bF����[%���|=�@h;i�<lO軛���B5=dk����F��������$=kjL=�hT���~�ŝ���~���L��������������2�����e'j�n��<�D��U���<�W�<Z;���7��;7:�G�1=�`�;=Aw7�0�B;]�y<:��r,=�-C<�O׻�֗��T2��󼷨=��=���<����O=��<�k�<p{=��(=i6�ʡ����JBr=�{�;���<u3�=*�+��Kc=4��x	i�[�h=�����p7==�<L@f�d��<ܮ]=�t=�(���/Q=a"�/=A�'=%,=����;<h�"�<�;�>!ӻ�P�:%{/����Я%=Ȅm���<�a8= <(<��q<>MY:/��<�A:�c�̼�=�:��M���;�474�A䆽�&N�U���+i�;�eP=,�;=D`�Z��I��<qU;�J�=zE��Z��O��M敻Cͬ���I��:�<�l�9�;1=7m�Q�R�1��jѺT\J<MJ˼0�;<<�<���<뀔��W�;��<�� =�Ĵ;�W
�Mt<=�y�<=���(�Q=98L�E���;K�t�d�X���μ�@��G�y���
�^2�C�L=\q5<�e���,�Q()��;�!�<���:���<��B��<;�C;�aռ�q�<j�=ϯ�e�b<��+< c#�$��<���;SՇ�3D_=<�6��m���䄽�F��N��0�=�&�0�����:��<g�θM=&9=ڸ ����Nm�<߁����h�h�&�*U�;<f5�Ϩ�<-�.��,���!=D#f<=�<}�A<�q;�4
?=���<���R@=�Us�W�8���� �=�L�<�Y��j�F���%��1��=�=��G��QR�a�K������n;�2�<q�g��)=�J =:W�;j!=��H����<g�=���<��8�F�B=�F�Y\���}����<������=�W!=���<��[�GY�=P#ȼ�ws=��<U�$�Д�*^�l��<���ѐ9=qB����4�<�ɼ�qi<�D=�9<g�5=&�a�d!�=�bi��Aʼ0d-����<�Z�<�g<m�H���S=l��RKE=��=�������=��=h�,=�ͼ[�=�9���.�<�C=�b<7`���<=�^h=r�6�LQ=��=	/D=��2���D;I��D3�<�v\��[�س-���8u4=I2&=F�90� =J�};=Ă;�SƼ"�7=^���1����I��t�<t���h^���;�I=o&
��:뺮ꌼ�B�<��<��.=��&<�~�;��=���<�	8�j�G�I%~=�É=��,�$�e�NU2<IT����;��=O=��= )=p�L�:{���=��'=c7� ��H�<�<Ƽs�.���<b C< �d=���<3}ܻ��X�)i�6.k;�Ե<�;<'[��%g��1�==�d��� .�C�'=3�I=̬W=!�)<(:d=f:=;=$�U���<р=/�4w�<��X=��h=]뼫��<��<D�C=r�Q=���h̼~�"=M�A;�?=~l�:��˼|+�<��I�w#�߁�=����7#�;�����lb��
ټq��=�<c��;�2ɼ�C� '
�^�=
O�<�i���(��[�I�����h�=�o"��2����D�k��M�{0��6�;��0<~�=xZ8�;�M=��3�?�݁���+�;��?�|:=)��c����� <x�ͼӃ,=��_�����»���=R;�����X�6�݀�<����V<=�r4</U<�3=]X�zG����<H�W�KX��3�̼�5��)�D=��ټå�D�);���;�)n=��z�z�;�l[�4�=�Yk=l��+)	=�T�<[�c=�0N<�6�O#��I=�)��4�h��Yl<L+�<A�_<)��<ͅ ���&=n�.�GC�����;��<N�L=��w���<�o��V=HҰ�z7�<�Dd<���<�=�;���##�;(�<@��<h����6+��S@=��2����f^�<k-=�z��N�j�<�j�<�v���WK��5=
���%U:�b�-=)��}�j�HP3��x��;5�6���2<Y�_�ςO=�����$=o����N��N=��=�[���2�;��9ʺG=:�;�żcnɼ��;�J�<Z�R�<g�����<d�<=G�t=�˜:�/=�P=��3�;[Z<Yz?��}W='H�ƞY���I=�p&��4=s3^=F"��B�<=(�a��z`�z0=3���Zٻ:�={Z��#�j��	�<Co<��2�7��;n�\���<�-�Fj�����+�;�W���=tE�<�e��^�=�TS=fz.��Pc=�/���bϼ&�<r�3���<�;��<��,=�Ë�Gy�<�&�=�CD���<���<��%<n�h����;��(�=%R�����gs׺�-x=<������Gd�<�8,=�I���v=C-�6Y=�<�>n=m�T=,�;;Pg=���;�<V��/��L����2�csP��I��O!���;��a��*Լ��M�x�;��e���"�t�6=2��)Q�<�E=�S���=e�%<6�s�O0�<�Q=YEԻ��\=�?�#�d=��1<g;<��4=��"��:3�ۼ�/�:ͩ�<��<2�ż��%=AxS��˫<�t=���<����{X��lH�L�<��!�]�=4Ӂ=��Ӽ�Ơ���G=�Am�!R��A����a=�c/�K���Q���;=hӃ�2rz���Y��	��8���ƙ<g�e�3�]=AN�<�M<D)6�,6��jKE�
��s~4=��=on�;݀E<��2<�W!<c�(<Ds)=v�u����<��(=MM2��q��j�廫<Ｑ��;�u_�WO �r]��1g�<�>���=�-&=�)����[���=aP��D,�����鼭�K�8v;R�L��LU���;o���R+=ȷ�<9r����:��Ӽd5�<��[<ɔ����r��%���E�޽��S���0!\=2 ��ńD�g���<:҂�᤺�Xx��n���R=DYK=L���^J=D\&�F�;{�=�s�;;lo��au���4�O{�r�<HcԼC��<��<p`I=,l�����"<������=CL�:��ɼ�WҼ�O�RK����<+IZ���;3+S=��=aC����;x��b'�;-/=�MN��2�#�⺶%=�q4;�W#=�O��<Ҧ<����{	=���<O���;�<��;��꺚(c=L�]=��ȼ��{�!�;�&*�O���4�;��M<�/��w0=��Ѽ��<�i=9V5�Q�	����;�	���fL=��C��kl�*p��*�[�i�<(d������<�|<u��;�Z��b`[<^�=S=(���z%��9q�y�b���D�0=$�=28���D=��@<�8��₷��,�;̌i=n�<�	�a�e���<����2�;K�C�;�T�^��<�yJ=��;<xu=][�<��=u&_=Z*��d��.��|/=�Zp=�U=���<��=�!����<�ء�������#�CT2<Vk,���<��	=���<)�ݻ~��X���Kp=AC=F#=�-o��޼�0¼,q=%�$<(G��_
=Tlü�C��Q�=�Vx�PN��}}8��,�<��<>H=��~�%�B=�=Q׼����1���<$�z���8=E�Y�4,]�H<�=;G4<�==�[0=���9�'U�]F�sH�M��<Z��$�+�{�=Xb,���S=�������4� =݅
���L�r�\=�}g���a<�������Rf=.߼�F�<c	+�t$��
�<)�!��<�%����s=2��:�������$?P=$����X=�Y��1�N<4�=��<���k�<�f���L<#��̃�:�H������۴��&v�<H��PN�<���<B=�u�<��P�'�=+�=�Ë����<I<�O�Ԏ{�IG���߼���s��^m=ɪ=Jx�;�K�-~8��[���<w;�#*=����».�<�%�RWE�;$<�x;��߼5����d=Z/�s�:���)���;�ߪ<�t�<��=TB��m�<E-���Y���<�zd=�5N=n&������=�}<�d�<�˼e?u<R�<Pq�<�= d< T�;HKT�lǡ��	|:0)u��jb��E��`��*[$��p;G�T�C�y���U=4�O=[��<">��4�L=�b< 8a=N';o���7�����<e�	;&2\<J';���|n�;��b��;�r�<.�D
=��L���X<�:G=�,��<�}<��<���<
n<�c=Q��<�g=��d=�E�=z�c=��V��殼
$6���j<~�A=�p��.�%�9ݩ<J಻�2A=�O/<�z<���<�����$<�^�W��;�t�~!�����9��C��9=�y�;q� =g��W%<,?a=d�iTg��\���}����<x`�.���й�]�=X��B����=�S��!=��<�%�E�.�eH�<���'��U?�"�;�h��*<��M��Ɵ�*sY=�>��&E=)����<��#=��]�<��E<=����5�<}A�<I]7;6&a�1,�<Ћb=�b=""�Ⱥ7=q���ӹ�:�l��ٹ��Rͼ��F<�p^=��u�h�)� ��tA=��黩�=�Zi=��<<�А�꙼��b1=�"t�C�Q=�b:��?B<�����=�Z%�{�%=�=���:FnH��`��9����Ｑ:м�O�G��NO_���=��<����<�%���<n]��;���<}��:>�ؼ�~��� �ZIQ�)�8�y@�':=��=�l�f�����#��P&�w�C���b=���"�|�U<�ei=�<�Bؼ6*ּ%��;�g�F�WDS�Ƀ�<G3׼�D�;*�<�ik�5}�;��%=x�^<�)O���P�Nؼk�<�g�������$��K	�TwF��T"=�`��E1=��ڕ|<eλ�8"���<��<��>�Tݝ�3���"���Z#��9ȼ�[!=�!������\ȼ&�;�Cq�>�9�:<5��<fQ=v-�<\��҄<��h=�+�<M�!�}��X=��U�=��y���<U�
H�<�
���<�z[=�Uv=�O��:��=�2���Y���<�bu<��㻊E=��������d=s���J���=$�d�6pj=��m=���;zW����;;�f=���������<E��<�e�S����� Rռ�\ <��=UI"=���<7���B	��<ii@��=C�0=��B=0ҵ<������j<>T�!��<5$#=c�,=[��<�h=�j��Od����'=�Ci�M�><$���
�ۀͻY�)��(�˼̻V\<�P��ȟ��x�X�;�==S���=渉=�*=��!u�;V0ۼ[�<��==wC�:�rмt��	�=`#~=ҵ�<���~�m�!2�;��R����;�i=�y�<��N[|��Kg=������b=s+�,�j�u|==�"=�����Y�<A���b�k<�T�<�4y�=�y=ՄQ��/�<4x�<��A=�ƻ橻����S�<������M�<���;"[G�N��0�M=`P=�<�c={)�}z��xJ=��<��5���y=��1<�����<~6M=�L��ڿ��̌ڻ󑜼�+A��Y�<;W�<�����<��d�"i)�:�@�}
P�E�
=�|B<PPA���';0߄����S�h��t\<O=���@^m=��$��![�U	�f�@<JB ����<�R�֖�;FL<�+d;��������%|H��X��(9�|I=N��C�ڼ�2�cG$�gt<Y��DF�<Ks��U�c�T��`2=Q�μ���<�=Ϋ=�G��`7���"�H���=�c�<��)<%|�<,E=�K2��&j;��V=�{@����<�\e�A)W���0=�A*<sqJ����<�^�<�V���4E;���;�A
��H{<*�<�=~	=k��:�e3�N��i�f=�0={H�:A^4��H��Q:�EOܼ�3˼�y�<z�<>4�<b���\c=�#��z
˻�,�ۯ�<�"=���<�ӂ�j�7�±E=*��1=K<�X=�1e=��j<3�2=?fú�O��Z:��U=u4'�;]�<r =]�>=�S]���-���+=��<�pE�YV`�L��<��^en=���4�F=/��k�z��<�3=�P=�k�</�ἤ��<�1B=ٜ�='�1�q��9ʹ�<81��/��K+�<7S`��3ٸ��<P�<U�j=V� =�="���:��"��<Zj�<g��;���<W' �Ǒ�2�<��<%dR=��u=���"X��L�S=�a =<�<�;����^=? e=cR�;�9=�=1=�^a=1;:�׼�$)=t��;�}v��<?=�ώ�"A^=!�R�,��T=��`�l�j��V7<�z�;n	=G����m$�����w<0v9�˦�<�S��[�Zf�}�'�h���:ML[<���<�;���{I`=��K=j�=F�==�.R�I���Q�=T*	���ՃE��k�:Pn<=)�_�,I6=⊽��1�<��r��-=��%��C�1<�<��e��<�KQ=q�<=8,�Y��<tn<3 ����*�
=n��<�Վ����-,8�������b�zE��4M
�`�F<�LB=��,=�^�;��8<��	=(�<=ħ��߳/�!@=o/�@�<��n��~�< �2�==�gA=�:ɼ�#="o����=�y��F�����p��<���9*&�<�S=?�N<�U|<$p�:n^<�E��ց��0�=��<%�=�H	=0K�݄	��Wg��M.�]T-=�wC<D�j��0��c���6�<8-��[=)4�<{�<==���	��.�<�z�;��;�N���P���<���<���qW�J7� y�<�%�<N�=�h�׎;�y�:��B��Ǽ/8�q�\�	E*��]K=ɂE=��t�����Q=`�~=�;=c��e�AS�:��;�$$�k�C�����`��;�2 �}u;?����1��J׻���>X<����9��Ӽ�)�$�?=eiD�,e<�8H���U=���T�_�eSʼ��%=�r�<�^.=�9��$�;�k"�mc=��c=g�r�-�<�^�*��<��j���⻝ż)�<�)�����;�#���;Ս=��;�9�<u��<%D��W{�G�<�>��V
<�
�����;��\=G �}�<0v�K��H�G=:�_��"j�\h�<��O��d5��It=L��:�wV<�"=���<��9���(=YD�A����ɼ*�D=#`�<�
������r�N=u��2�;R�<��a=������;:#=ūټ�X=Y$=;=E�<: �<
�#=kx>����</��<��!�`	:�?M<Cf�<l0W���
����]�"=�#S=LN�:L�V���d=���4!�<qN=;3�<b�����C�
�?�"���/�tqh�z���9=A�h=ʢp;�KA� wW��<��g��ز�"]�4�=FS��м�	���U�<�rm���<��4��=�u��鰺�9�;l�m���$׼E�W�a-=_��~��5�Q=�9n=�?��߼]�6�����5�=���<�>`�(W=���<t�2=��a=�+�(=�&�<�)�<�1�<ӧ�3tM�u&�i|�=�%=�e
��e�;�RV��ӿ�iaܼ�(�<f��<�(ۻ'�I�7��<i�»�w9=����k3=r��&�����:C�:P����Ns���O�*=y�I�7�<�0U���I:��=�W=��=�h��1<L�#��;���}<��{<Az<zl<�݀����r=H�3*2���j=F���o�-=��~=?��<�]��V=�i9=�����,=;��<��=(B�<�KZ=�t#=�l�=$&�<)�=����Qm�8G��@��RU�PF�<���<��3��K�kd����0=Nv�<�y�<
Q=����};
��� ��<~�=�X�<�'0���<<Ҭ�'�A��P�:��l���<����D��/�d=�u����= I=A[=i�����R=M��e1h=��H�&WO=��;������~��<~"f���)=�d�<B�i=��:ۼn<����n=�/=G:n<�2W��6��@�<n�Q�St�<C�G=�3s��D�SN��PO=u��<�G,=��ِ<��M���<5r,=RQ�<P��=/�/=$�-[��D���;G�u.?��¯��Dt<��B=��伊D�{P=*�l�G�<ϩq��:���=���<R���#=�ɂ=R=X�;Y�+�=V��C�<�r����A��V���</��<g*1���-�P�U�%�+�?$%�a�c��KH�p=��^�ς��-��`=1RC=�>3=يV��%C=�O�<��6<Ѡ^�r�Լi�m<��7�$�����;�-4���<�#���l�M#}��MX<��i�:����o9=��μ�<-��1=����k�d��ʃ;�켳�^���O=�i;�� =�p�:�~ �k39�D`��)�5����<�S=��=v��<�\׻x�P=- �<m<^'�<Q��<�$===M(=ʳ+= �)=��<�8�C��<����Ȃ<�M�����.<9�� D�23F=8�	<�c=����x�ٺ=����:�.f#�[�f�~1e<_��&�<�h4���P��:�<?g�<�
�q=[�<��G=�=R��-��3�� ?�&���ۉ6��Ā<�� �2�=��<؆�<H����s�J��5��<�R6����=��o�P �<��r=�|�<%������<-�$�Au!=+�����л`c�<8��]�;^%T;��O=��~�a
d�k����"<��;�U�ğK�����;.V=!Lb=s�(�|`=`i�����vH=�H�U;O ,=��[;&~=/��;��?=�� <�f=�kn=�n��;#=���;�S�����~�;=�*�<��o<2 �>�����=X�����7<��<�b#���J=�e<�,n�<�S0���(�[����]��k;V�.�ͣ:<{��<�w=����VR=�8�=}E`��R<v�C�g�=!�<"�ռG�ϼJ�J��i=i=�≻���<�~�;�vW����H0��$E��,�u*�<L�a���J��iE�(�g=��s{=��<�4V=ϝg=:�C�6��]=�a�¦Z���
�֎�`�٪���^�<D2D<�Z��ż�=�Q�<�=]=4�-��;�<�3һG�A����<Є�q���P�R���bf<��G6���x��w�;�鷼w՝�H�6���<zy[�wƼa�0��S=kH��<�SA���<E�R=�9��1��������<��D=�\P��F�(�<� p<7ZY��4�s3�&���DJ<,�r=�KX��?6�<��;��Ҽ�t,�b��<v;�@�?J�<Bw�l	����r�p<�4<@W�;	=(=���<�e�<��=�v�<`t9qG�<��ؼސ�<�M`�_�ܼ�t�:UWY<���%J+=v��;�<=LG��J�;�S	��v��q�;��3;�<�μ�.q<����F]$=ލx;|]���9���ʺg�x��봼z^�<�s��P0�Tɭ:A�q���q�I��< ��<�mT=��}�;�C�e璽k[4=eJv=�v�<�x>�p_�<Y!�t��<���<&TN=x==Y�弇�<m�����E=5�E=��<��̼3��<]�<X�:=ll=<�6̼��S�h��<�u=X�=�|i=�1'�'{:�*����=���<�k�"6=���fh&=�t�<�Ӧ<��1���,=��;8*P��	q���{�����м�瘻�s��i�X<K���.2!=x���x�
=�0e=��<�=J޼'=��L�������g=���ӧ='A�<:�>�f��<r��<��u䗻_�=�
��=���<u��< w�<Kݵ;b�ټ�������e�_���O=�7̼N=G��S==�s׼��<-K�;K���|��<�ϵ��%Ļ�	'��D<���<ҙ��A���eE�~Z�{?4���=�^L���p=��<�,3��B=kJ׼�l�;�e=E�@�?�ޤ4�Q��X=�w<<�4�;~sC=�\�<[ջ̦=���<nD����q��y�;xS>=c^�D�:�<J���.�}�=��1=￡����`�<��<ҼN���,$P<y����<�;(<?K��	z�;y)P��=MAB=<U�e*�Qm*���C!D�M4=�ּI��-����r�<)�m���K���ϱ<�N<�����E=�4=y�1��H;�)�Ȕ����9=�M�����G=�j�O+=�9T�"k��p��H�<�^<�~Ǽ*f����<)����~;[=�꽺-=R��T1)���;=�����,�&����<��D=s7J=�H=���<z�"��]���=�;�&LL=�r�<8����_��L����oj=Y%�h�3=9�1Z��͆0�n�<�B��������<w�=�c�<�AD=�=�>��)H��;�j���5<��<F=�p��vM�;Q�O�J��<�=0��<�1���=��]<����O�� u���`-=V�
�*%�K�{��_��MҲ�$b,=]�\��<��I;����P=y���4[뻃K�:��<Y� =�V�<=��<�(輢��<M��d�=}��<�]�:�7�z2,����<m�=�`<���<���<� =��:��i;i�c=oD�<~i"�q��;�(D=�4<�=b���(��:�͵:�+żf\k=Ɖ
���h��p=���%�G\==R�1</�6�N�=a�Ӽ)�_�����A�<�(�>Wż�S���A+=���<���<�p�������-=9�(��;<ļk� =��<�K�ڑ=>�=%��<�M{<cxm���D�� �i`��=l�x=}��yX<�A�B>=��I=r;�ᔂ=e�;`'C�`� =����y����/<��7�^�2=¶o�[PU=��#����<����e�;x\S;e[�����C=����n;��IJ<y��^Nm<�ټ<�2�
nI�'m}<��T�����.O�b�m���6=��;��t�y�ȼ�ռѡA��i�;���<:�h����.@=;o�:N�6=$!=�[&=U��(� =~0=m=��o��9���:��j�=��=7�Y=QxI���o��9=���Yn[=���<���=��,��o�;V�^���L��ǂ�v-�<�9�<j�Y��=A ���YS�!�c�=Y�����<<�>=vᔻY-V���=��ոǳ��ʥw�DG=�������_����D��ݕ<�{T=f.�<8�<�1<�$�4�j�;��N=h�!e�:�-=O��I�,�S?��
=�0=Pʎ�!Z)=_�I=D�V=#��<,����=�N����5=�<T���L<=!=��U=b�!��e�:mG���?���]=�WF<��N���)�]�@=ÿ��rk���C=8lͻl]`���n�$�Y��� <�N)=�\�z0y��T\=�A=�gB=q�L�dI����V=.�<��6<�74=��H�Di=��_��4A=W�����a=ai�;G'b=�9)<��=��^-*=��<+��<?~&��^P�~�u<�DJ��uc�?c/��<�����8i�;N�s=��=�L��~�<\�6�a�)�7*=�V�>�<�H�:�b =Zf�_���H��T��р��a�}���b����У>��2'=-�q��B�;��E�3s�#74=��N=X����=��h�<�	O=�j=���ֳ�<�P�;�� <q��S=�[�<w�<�������9}��x)���<�	%��/(���g=�F �*�[=��/=��:=h�'��� =/.=����]X�<�A:=T\I=��7�	�<7�g����<�`=��V����<u����+���*=:V��0�6;���<�=��I����E9��= ������g3=9�?��!�dr�S�<�R =���<���;3FI=�T�:ķ��j@�ޒ<�r�<e�V����:��@<��\���;�a=�4�<�MU=ݻ'=ws��5:�<��+=s����+!<��t;5���:�t��b����<F�`��sN��`%=�~#=.�����$��<�<���<`><9ϼ��v����;qޙ<��\�j�4��\M�ֶ}�G���*=��;���_���<���<�=;D\�;��j��)�<��U<�=��Q�^:��<x�,�C������ �C0��W߀�("��xh��Z1=��&=:�<$�;�:=�+:97P��R<=LF�<kԻTY��=�2<Y�<� =��G=�Ǳ���;��=�P=���y�<-\�'�����i=�7�����g	����/<�����\��P<Bk==�p<YL�����r)= �@<�	`=�e&=*�ռ�g=$<<������x;��<�'�'G=:�f=vZ=a�%<��</Q���IM�P�=�N��Dk=eף<h�<}�R=1s��>=���<]<�<{5!�*�=�k��N<
�����yV=Er���.=*�<�
2=%�<�/��w�$rX��=,�V���<�$幺/˼��"�(���4<�=��=���p}�h�<�5=A��<m79��U =�|���Ǽ҇V<9�L��n���:_���;��r����߼� �gB �u�{��� ������?%=���<������-F�k2=�6g�B�� Ko= ��?����<g�k��3��2��/�R(<r�H��-�����?�=!<=1&I=��='�<9�=����r
=)ɒ<��;�DV�>�8���Ό=!��ۨ��*�s�Z��<4�=��<�GI=���
��;���KG=��G�լ���=	� =�Z���0���"�<_��<�"��sE=����� �<�q����]�����=�/��&X<^����E��g<�M�:��Q�MN =L��<�D=tQڻ��5<�`><Bj�<�FP<�?��k����<J�;JGi�Nl<(;��iRV�5A=� )=Pg.=y�<4�Y�M޻����.t�=I�=r`)<��=�C<Տ!<�q�<��h�<�\M�3s�<�v=_�5��Zռ�/N���9��̳����<�ʙ;rMv��8���0=������VX�]�*=T�	=�ջ�ɔ���ǻ:��<jM|����`�ڼ0W==��ü��	<�6<޼�<HK���9��j#��d<�̛==�x�0W=�u<�(=^���:�m���$��!7=U0=z�+�Z���!�C�V;�
=.v�'��o��<���;윖<�$�1�T��5�>�O���<�5=��D���o7�jFE�����_�|<���;f�#Gb=^u==��M:ܼ�}�<�N3<����tC����!W��`i��ng=J4���;��D�<X?��J=�E���0�T3k���m<=�n�@�@<�󖼙����N�y�<1f �˷�<�i�H�{���;U(Y��Q���<C<�>�B:"=���<���<Q�x;{k�<�)&����ȉ���1�7�U���[|G��E�<��=[����-�ݼ�mX���`<��<�a���\�ٸ�<��l�J��<��6=�2[=AGI���z`=�_=�_Z=	M�;b��<\d,<��+=I��7ŻwiO=�n|���2��`v���N���<=v
�<ȟ)=�]=���<͊n=0��;�$�i�-��TG�˻���<���]n�qx<�$=>Z<�m=��<g�>=ܐ=��W=4L�!�_���[=�<��2=d�����༳%=9/ �����}l=��s����<�]<�]-=A��z�u�w���zۼ��\��~L=� �#�<�
�<�>=8p;�+\=�z=���<*�b�!P=�W�<����S���Ļ�
�<|���;e<���R�f��<�����<�T%�����'�}mX=�(!�ް<<<�C=�rp=<e�鼦Zj=s�i��A@9�bu=3���ͪ=:J�	���>��.��<w��=r��<�u^=븠���=���{��U�5=��q=�w�}�%=PtW<�9=&ּ�k$=�0��8��<�����;���<��=WR)=�Ӽ9�a�.�|�$��ü&"=Q�=(�<��ȼCNQ�q�K�@�;&,=|Xj=�6�<
8�ޔH="V� xĻ�ђ��uE<�ݾ<=�r�yU=��Z��9t�P= h=�(�;܌�<��'<|G��xb��S����:==`�+�Z=�ی�u���� �=��"<h:B=�'M=!�����<���c�n����{�<�_1=^8R=S�;"m�M>=0�"=��p;aH=��K=�xS�ආ�0��)�et =\*
�oD�<�l��L`&�\Ul=��<#"4=9]��0��;�I����<
-<�=;I�:_�;����Xo��qp:=���P�3e�:z��-5=�[C=���8�xh��
!��\B=0*�<2+��q��`|M=O:+=�2�;CM���X�Ӝ�;��Y�� �<{9��	S='#��Inu��*<U�:xp
=dҥ<>8�J�^ A�x�<}�\��=��+�$H��]=;X==�`w�CFH;��ȼ��<�+W=�c�<����uG=Xf� �<�5e9<^i�<��=8��<}�<�-�;�ۂ=���{мK�:�6R���<=�À<�{9���D����<Wf�<t��tN�<�"m���#=�4e=��:WeT�YO��;WS�;�N<���#=J�	=�U)��x�<s�R=�3E��z<��&�o-���O=�V�<e�k��6J<��f<Ǘļ%G�<7œ=0�<��=������{k=K5��� �<���<6L���u`<�h`�̷	��'�a�8<r�=p3�(׼g#׼����s^�P�=���Y�q�vuI���L=�q0;>�<W=�꺙3��%��<�#=e �RI�����<S�=����wǼ�+�;i��:.��;�:=�==E�:=&�<���<|Zc��;�V�K=d���=~<q��S��$�;��<j?�<kҼ���"������:K�'��m��/�=H�A��z?�0�X<��ɼ�~=h}=y!<1Zj�
h�<�d�[u��J8�F�b�z�~;��k=_��<#7��"W#���":���؛(���������ZEB�ȸ%�J5};����oԼ�Z���T�?8B=���0 �8�Ἱ
麅�L�ם;e? =_�;������C<6�=L��<fd!=��-��J�A'Q<K��<c)����<�ɺ<O�H=����Qm<:�<���<ta:;Daj=�e�y�=�(�S�i=\�ۼ�=^G=�̣;vD�<Jo���\ռW=ބ<��.=��C�b�<B�=����Ć;�&����<D�<���K�=�@�Q�I�&�}=y8ؼ1�n��==�Kj�C�k<^rX��/�<ݡE=�5��5�׸/�ļ�1�<(��؝�<��<B���QK=NmU�SD<i�[��7��;��o=}�/<r��<c��=g�=n�3<E��<!f='�1=��l=��5=%��(�=�ȼo�#��.h<Ջ����<N�
<��<�<���:�T=��;��<�b�7��@J���Op�Ib����O�4m~=��<�:�I�U��d=��!�m.@����<�듼Ȑ�����R�<y�^;�'�<'.1=��_=ofD<�|;��#�<��=eK�<�:<��5#=c�����N�Ml=�lh=�t@�n�r�V���5Z�d�l�cR/= g<�;�;�m=2F���^�<�ﰻZ��<	�����U=R�;Myۻ�	�jӁ��q1=y��<�=R��������j��$���6=I'���>�������>�<�+=<�o#<�g���¼ꄫ<KJ�=q�;@��f�0=��<qû��<gU=i�}=��=�Yf<�W6=7Q@=�`[�9�<?�V=*�Q=,�d=a��/�]��C��^��;^�:U���7�I� ��:c�"=d#=[��090<�gw�f򙻂W%=�"�=��=,�R����\<��*�x]=��=�M�l��o��<�N�;��;
�p�{=�C�<�^P�v��;4�<��=�#(=�Q���*�<���;=�߱<�'���~;�>=��<�@9=7�<�Y�W��s��
��J�����<j^��Ӹ�DB,=r@�;L�<�F��\�z�i=
Wo� (���S�'�0��=�(=�_�<MPA�9N����<u�A=�q<��6=��)=/+;11=�"	=\`�� @o�}!�<@����Q��"=�	C����;X�t<�kL�Ku����;e��?<�����RQ��M� XC�.����0=�\/=��B=��_i��P�<��=�k=�O>=�u7<<KY��ص��$�<Z�i=���<ܨb=ԛ\<Y���dI=�:-���0��m�<.#��I��\�����=�]<����;`���3<[��u�<�7������`�C<�9p���1���� 	{����Z%;@�S�L����B)=Ĕk=���;���;	���uFp<�x=
� <���< D2��p;~�w=L|��U�;+L�xxr�+2=>g��o�<��a��[�~�֚+�z�K=3�W��*�;@Wo��==�o��u���=z�|<#���X=y)=1/ɼ3Ƥ�?�0=��=l@�<q��<�l=H�ƺKB�N>
=7g�-em<��<E%�C�����żB��<偉���5=����]�?�R=�;MC=.�=�쵼 ���̼j8��gnC�?�<���<�Q���&=j�\y�����<�=h&��q߼�!�8���־��S'=-=������*��N=p��OsA=�w��=�B3<�I�H�@�,<{�����e<���9��v=�]b=+W�;�5�<G<?S!=�œ���4=F�<=��9��̼�y���En3=������<�H�@*={�=���<������Jn;�2�9`����=�߼�.���^�=HȼSE�&b���in=�ؼ�9�7;�:�]<�ɾ<�,���v���=gN�O��	=�N���<�!=���<��������D=pm4;a�T��g=٭��GO����<ȋ��sA=s�&�`[=o?�j���)�U=�u��L��<є=&d�<q;_�R ��r=0�?=r�=�6)=IC~<E��(2�� �<�	G=A�R��]R��h=-Z����]=�=B�t�5��;�Q��
=�~)=��[�T
;�;8l�<,E���==�n�<t�<�_==��[<-O = H=#̼��e���2�Į5��<ѻD�W<B}���&=�? ���1<�A�<l6=��0�\������
=�vF<��!=��[=���B�k<Ce.<;-����<o�@�P��<��=�)�UL=��=�D����B=�V0;r�<��m�g��;;<C=	�3+�߹鼇�b��~�<c�6�xM=m �8��!�<�<�啽<~v�P�*=󆠼Kވ</=�<%=�߃�L?��]��<M��:���n/�V�_:*�9!X=L��<�S�;5����N=�@��	�!��yK�`9;����&��w�;O�+�����<�'/��?�u��5�X��̌=nÊ=O9 =<�"&��<̼P�<U�`�8�=����gTY���]��<�_��)�<�a,��;h<c]�<�B�A�����<G��.�<N���'v�t���C�ռ�~�e+B���W�T-2<��5<��ȼ��ؼm�Ѽ�U�<�k<R^p=�u��<��t=N?g��ӧ�L'����=��><�!V=�L=�<O���S�7=��;gu����=��ù��	=㦃�Beȼ��<���<>虼
]�<9�E��B�<��j����<�m��A*� 3��w
��B�<W	l�g�h<>�a����<A�ټ�.��Hͻ2<�W=,��lT==Rk~=�*8�2$=s>=���<������,=|bW=K�g�>y��v�5�Z�ż�G=N��⒏<����p��=4B���<zR(=ԜD=q�<vSͼڼD�_�7��y�v�4<������S=.C�#Dڼ�(=`�<�(/=X�\=�I=m^�< �'=��;z���o��:�߱<(o�x(��̳=\+�'	=1�0=W�*<3l���d���<v�ڼ�OT�]m�<�@M����<@0='W�9�H�U��;ւ]�� ��9�=:{�;tO=9L<������=�g�;/7��;LJ<d�r=a�Z�í�=����ʦ��O�Ӳ��{����.�C��i�x�������9=�����g;�aJ<���h��zT=�$#���ʼ=,�,!I=<I�<96N�Pǟ:Ӆ３k�<d��;���<!sg=g�c=�W=�)=^�C��o<	&��I�e=�.!�J��<5#V�v�<����B���s�=�X���<���)���F�-�=�n�<B�=�NT=a�q<�K��=� =lc����w�_�<[�'=Y��<,v��=�sJ=S�$=J���\�=ć)��*�<��8=V9��$)�*�<��ݻ��=G�=ѻ=�d=n�!��y�i�p�'"<=F��m*���,=M�:��N�<5k�_.=*~�<��"� ���]i�s,ɺ��)��Z v<�$��b7=�&=���<Vw�9=�>�<i�l�9#ݼگ<�!%������V<�B9=R�;Q�`Ɣ<w�w��ݤ;��=<��<گP��2�����<;�E<Dͩ<�L�<�T��E���*F=�Bt��Z=�`Լ�L��ps�<�Q==9~�<�l)��p��#���-���O=��N<8�P<��:<y/=�'�<|Ի�e8=�M=�="U�<�M\='����B�<��D=�-n�ʽF� `׻�&���p< �>�هM���߼!:+<�����2<����<�����Am���<����?����;?�=�X�<9l�#s?<�$4;��������x;�8�\g=suu=$H=��\=aq�S�[=ʔo<���<|���|?��'�G=�����.=I�$=/>v��I=��|=YZ;�`y=A�=��@�g�B���B=�r�<%u���X��++=H�x<�)ļMȻ��n<�Eq��_�;�����E�E��Ck��W,=��B<{:�<Q��<��^������	=b�<�.h<�ֆ=�V���Z��M<~��E�;_��<<����yT�Ks1��n)�Z� =#=�9@�ҼŲE<CQ<E����AW���=��(=��S=/�>=ު.<�TZ=c
@=|,
�"�v<��)����ż?�R=ҍ�̰����'��q<���<ļ#�Z]���e=�+��5����켞��<��-=�(��u=�W�8���J�<����D,��?=��
<5�<$<�:~@�Bz}���ּ�Q,�I>M=��?��DĚ<���;m��;%��<n�s�F�C<8<���%<5><�QE=&ㄽ��<��:=��D=�>��@w�-��<ݹ���$�<T!��)�ӻ��X=搽���<���<�樹��x��}>�N^���=D�<B�����$0����=w�<>�	�?+Y;���n#��D�<]j0=H!ϻ#��<K&{=�μZ}ļf��<��)�S-;;����k<a<�-=N�=;Am���F��G�$=���ݱ���R�Q�=�@Z=w�K�BY�<<F���R<N����<���;@O���a=g �;��=�l+��J=�|=�? 9d0=w�7=�AB�3y=ud��2�@)¼[׼G�c<v���V#�¤'<��=/^Լ:�<U,��c	缑�J=���!`��Q�漀jz;��3�04׼�K.<zqa�s�c=O*+��]�9?8=��e�$�B���&��<�Ŀ������0=hb�2�="��<!P���< R��#���<��<JFL;8�Z;L���y���}�&�£=�o�<��+'<.T;���<�u�-�W�G �<���<�M)<ρ�<����-��=��^�<�'��N����o��H+=��;1�Q���<#u���<���]QQ=$��<fNi=�>=�T輫! =r�4�"i�;eB=�F���%��e=<K�<2���b�{�=�qj��8��e#t��:}�YH=*-=�*��m2=�<�ܬ<a_��;F���V���=F�޺m0�TL=�`�B�q�"=���<����˺.F=�E�;��`<n���'�	�b����<�"=X��<��@<���M�;-����>�%
�<�&0;�<ŻP<��e����<h�_=�2�<��k<��I�x�_�^��5�R=�P=k�߼T6��-!<��`9"�N=Z4���W�|&�9MgC=C4\��C ��1��#=3�<~[b���<�xK=��=[J�<e�<\�=+�}�߲�=4+=��e������ڼ�F��CV=�%5��-�<�)��i� �X���=;��
=�-L=-><f���@	�<+ɬ:YT�<��5==�ԼY�f�1@2=��k=�V�<G�U=�C�<��W��L;<|��ʖ0=^ؼ.��<���Lb�t�<`�p~�L7K=�*�"v=�����<��0=���<d�׼�E;�Ҳ�yc���E=I�޻܅�<��.=O1=��=u�%�:%=��Ϻ;ߚ;�AS����U������d<
"��ʢ��<=a#�<��ļ�"�<�7i=8��N0=,�p=>��<4"�ɳ'�l|���m����<�<@�	���(�3�<̶;<j��<���:3�=�N�� ��aY�</=a�]�=�%�<ղ�<<����G��E�<���<��.���޻c"�<
�-=f��<ǫ<��-�K�=R��=�I���<F�=��]�]%�:�3� ޷��/��N�<o��<'�<�G <B��?�(<|�=`�E<m]=qO��H?=�x���n�<JM=�=K��ya=�5=k�\=��<õ���2�7 �<'/���P�<!�'��{h�<Ş\=��\���+�5��\b=<,�:�ze<$������,=[>O�p�@�F�d<����~>:DS�=b%�I�P=�_��O+��;v=q�ct,�yȼ͝A=JW=y��t��<K���0�=V�1=_�b=�#D��ݻ~�r]<�ѻ��'��U	=�>�<KE��� <Q9��G'�<��p���К&��i��b�<x{�TA	<d�=63==ϰk=ȁb<�W<]Ը��im<MH��}N��$=�#���s<M|%<�:��#*=������</���P'�ry<=��!�k5�<��-�=D [�%��<�Y���e*=�<��;�'���|=�1=�!�<�\+=ǚ@���ż����n��<��b�R�"=�M�<�?8=	=�g���],���<�Nv��]�<�͐<Q�=��\�Ѵ�9���<l�_���C�7��<�`@=1�<M�Ӽ+�J���D�M �<-¢�aK<�׀���=ki-�����6=#V�<�0"��<t T=>R=�����=j炼�5���=ˬ�<61?=�V��ּ߽2 ʼ�T��p��PX;�,��N�Q�.3�:���A����]==�<H0�tzP���k=�=F�F=w��ժ@<�g���;=�o��6�<`3N=��=���<�;�J��6.l��E��7ռ$�=�xk��F�6�Z�=�=�A<��l���7=J�,<HF��� �<�'a=�#<8} ��&i<?�����+=��6</un<W�3����<~�c=�X:�=e�4=�.�>�/=0�<G��t߼G���=��F��g=ᓚ��)w<O@<��=�(мL*6�u$=�E�<٦c��\U=�= ip=�?뻪�<!J=��E="1�;�[�;=��;݈r�ş`<�_X�-`�=y_:=�/����;��_=[�_�S3�Jϐ��y=��D=d)�U�j��G=|N�Z�&<l
�\X=�JG=
�"�I=���9�������
=��&�=
��<��A��=n� =�L3=D=~=��)�*[��E���b<���<q��mp����;-�=��<2K�<	�x<�M�8��<�2;��5�j_�;��!=K6���7�=���;��=Ͷ=�D="��< ��<o�O���ؼ�^u�a"
<�մ���z����\`=��>��+���:���<�<�'m��n�:b�8=��=�U���	=-z_=�?(=��s=O�R���!<U*J=vBM������A�j٦��cS<��;ж�;J<C�<�t�;�-�=�p~<QO�3j�<z ;�r|�=�R�F�.=��7=L�����@=�T=
�=X8�<4�<��,���<�C��dGO=�0=�&z<�%/����<�;D��eN=���<�i�<�-<�N�[v�:�h�<�tj��?ﺣ�u=W�/��f����!��K�<xr=���:�D�n^<�cW��O=�j=�=;���=$=� =��=4�S=֮���K�<��\<$`�<N>>=B΀<����N=�����(=Q<U�_�}7���=�T=�'�<�V����;$�<�N��aR\=�������oz��y ؼo�<�81=%M�>��<XAQ�Y]<�&7=R�:<����M��J費��F��O=���;��L=��-=1*B���m��4�<@"���:�S<<�����;ە�<�V"=2$��1�":[�+=�р<W�M=|E���;cc���n�=�:ü�&
=Gy�=��3=�׼��~�h���᝼��\���"=s}���F�[������<�,��P��=��q<������=T�E=�'=�?$��C7=�O���@�����<��̻�<��.��<*�<�K=-���Xz�;��=�5&��4�1��<��:�礜��Zϼ�"=G���ۅQ��y;�/�����~Q+�����L�ni�;>G"=�9 =/S>���6=t	�<���=@��/8=�W$��NL��Il�Ą;�˝A��y��Ϸ�<���<{�=Q�o�uc�<��7=R�=Y��<�zO��)=�KD=�`����j�L�=|�C=#v���^�����|w\�z�<,����(��G�ݪ��j'=�yW=s�E<�6=!��<��H��qI��=_��<�+��v<�O��?Ͽ<%a7���=]�*�-�/�����r��Z�/�D<��0=��
<ܥ�<*$���0�D�/=��ټ�\=�@J=�㼼u8��n=��Q=ח�='�<�r�P=�D=iq�G.����<'݊����N�üum"=�N�@��<�!�O)�592=/�;��<�?U=~PI=M�J:�c�<�&��5���=��"=���C��� h��t�_�F=��8�v��:=���9�U=iJ���U���(1�p�]<}
c��d9���<e�;��%��	U;�L)��N<��W�=��J<S��<1}T�|�û��\='�>���[�E<�P̼۔n=��g��E;��;y�8��?=d/�!P^���;�h=�]Y�^-�<劏<��N�VcG�:�b��Z=�M=����J]E=���<�Q2=�!���;<��<���k,I=���<��摟���E��Ɖ�&�'=��+=7=��?���ύ��̾�V%]����:F�	=7�N��������D��4=^(���7�;�
��;� =��ɼ�#�P�޼;��#=W�=>=�f=/�R;6+�����<�8�Ã������{A=V�'�{�K<V<?<�m��&�9�fu-;�y�_���/�R��91�8��CN�_����3�`�<~yi�jop��$�<8Ϭ��rͼ~i���yu=�c=��c��Ɂ��(;���E�?�f�G�<w�<����~Gq;�ռ��<9�<���<
�m<Q��J�=��;��Ƽ�l=|wU=p�_=�nY���=@żu׺<kߢ<�H޼k��<}��%��;�'$=�?Ȼ������2�k��kBA=/�%����ռ�2����=��;%�M[���μ���<UJ��4q�;�g�<�_����?�Q� �C�!=}x���O�HC�<�GU<���:�O��1�<+c�@'=�g�&-=N�f=�O=��8<�+�XܻY�z=� �+�n=}y'���C���=�˻��N; �û~����Z<¨޼��B��j(��N=J^D=� ���8<R���;�zt��-޼G͜��U{=¯<�Ƽy������<%�u��-`=ӄa�f�=�	=�M=���em<i�X��'�~vZ=-UD��:��K8#��)��7=�}G=N=7=��L=_�O��SD��WJ=f3O�?#=�c��(��\�B<:���<lj��P=���;����?<u�H�w�<��0=��k����]W<�6<?&<�ܗ=�y=�|���U�R���`���tt�<�1�;��Q����pKͼ�_�+T�v�<Ĝ����L�4�*�=��
=�j�i�ż�w���ή<A��=��?=mI�:�R=;��F�2�!��<�]M=�$C���`�*�ü��#�H�=*ż\񈼿E��vo����;'%�@�=�[�;�d��*-�;\��?e=B�T��N�|�V�A�t�KB�F=�8���=5���U�h�ȼ	���ݡ
�g�<��$=#��<��v���$=(b=��*=��	=!g�<*�d<��[�rr=���w�<-�`<-��E=�Oy<���<=\����;w��:�I����3=�"r�:�=�.��k= ��;B ��-�<.�=%xY���v�F��~P��&5�M ������f<�`����<'�s��,A=];мA�K��༚�׻��}�H�s<�<���<<�=���GC�<�д���F�@��{=��и=5Hv�M@~=��������<i*�[8k��"=R<=��T=_N�;�ho�Pm��薮�'�ͼ)�������j<��Y�}=�S�<���<Xe :@�M=�a=�l\�F�:��-��b�=���<:��<Ϭ�<�#e=���<��=V���� =4H5<)��<��k=�����<5Լ�l*�0sU<��h�P:��
'�١%=�𼿢D=��7B ��+3�ᦻ2:�:�ⅻ@N3=�>����<��W�YX[�;����=P���m7<g����»Z��Z�����W�Iѩ<`'5�r�5s$׼�I����5=9ճ;�2=/�:=Zݜ��]<HM���8=�F��+e��S!�R#����*<��-�?�D=K���0=MXH<pۼs`
�t�P�Tc=�=��ܼPz���l����e���s= A=VE=���<W&���6�<��<��=
�+=��ٻ��Q����;Q8;O�D���)���UC��L9!=�-	=���<�sż�F<tx`��_=��$��Q=��=xJ�OE=����=�=�>�;]��<s�i��Φ<�FF=�­;8N=8�p=%=s&�����<؊��L�G�P= �<"
<K�)�d\���Y��(�<L6=��]�c,��@,��!�;HR�<��U=�X <�CM��t=��:U=�pF�)��<D�;3Z�<Ĕ�;�=8]��b�<ϧl=�P,=e��9�?5<�E=��c=��W=�`����k����<�WS�F�R=���:����"�*����,/�<�fB��?=S D�u�=�u�㯇���)=���<�A�����L@���5=�(�ゎ�K=�E�R9=1*=H鼄A��LV=��<="�<rW=Rٱ;���:)Q�S�=�C��f/�	f��#?=p��<��#�ix�����<U�ں��M�+�#j��[hP����q�R=��?=zé��#F<�0o�����0T�<3v?��b���+ =��=� =B�a=�&q<긼��[=�r=��ؼ�=�%+�<$�<�A<R����<K6�<��`i=��l�<R��H���)>���=R�-��/��7:_��T{�S��O���S�<���`������<SL��&�<%Q[����<�1=���<G���7��<7)P=�f�����;p���)H���'=kI_;\��<T�K��vf=i�=3�������=�@ἕۼhC=ν�<��7���<k��5�<P�N�%���𬼳h&=��Q���<��<^X="1:rS<�z4:N�Q:%O#=0��ۑp<�<C���.=.HU<;a�;�!�����;����;�+��dW���=��5�-q�<�#=�	�<<�><�ɼ�9=4�^��K���=�Ev�[�L<?�;&ct;KK=�J=RH7=ȥ�E�\��nF<�Jټat��G��`��#�=}��<��<&_�<(��"��<5��2>=l��õR���/����;�e�ҳ�ˊu<��>�,���;x��<��<�Sc���aN�.a��N<�"=�=�\��<�$����"�<P�<�yy���o�v��Q�<�j�<C�*���2�fX�;C��f�x![��4���_=����k9W=�b&�;%��� ̼���<	����1�p?_=�3?����<.�
��L�,(=q*#=��=�eM=�#��6F= �M=<�;���<MK=��j<��{:K�;Lq=<��`���D=��O��(=�#A���<�N<_J���l��(���	�[U��D�}Gg����l�<��U=Q=򬃼�,=��+����<��+=��<H]���D��˼�q�;D�`<��<H�	�>�2=�>��ܸ�ů6=����.�<��<95ڻ�b�R���08��ڼ`�9�E*�<9Yv��C=��4=�nμ������
�<�G��z9�*M�o?μ�C����G��+B�M+B��Yh�H�y��w�<~si<��"�,�����&=��'�I~i���N�	E��H*���=��̼7b�l�ڼ{�p�wK2���;�������=.��<#�F�U�8f�P)=�N=Ox��~;=hX���'�7�<E��<�0=�Pg=�@�ɒ<�w+ۼ�_��/���F��6�9��
=$��c�-��`��<!��<��Q=na��hc���^B�M�Ҁ��������r=F[=�,=-�.=i��;�z��j"=��м&�ռu	����Ʉ=�)*����;��ҼP9μ�+'<hs�<��<������;Qk'��峻5�T��ĵ�P�X=���<$rJ��X;��l�,���=W��:-nS���I=],�;,2<��b�2�f��c=�62��Y��sǼ�,C=�01=	��!�W�<��;��W����<��̼�[���p=f��0�;��b��d�<v댽l+
�.��<0�ޖ/=:0�<�S��d=OY0;��o�ɓg=1�0=gd��Jz;��+�&$6=5]\���"=��:�D%=�ha��}9=����2u�<���<U��b�5XJ�3D6��+��=�����_�O*=Q���O�<����y=1=�JȔ<\a��[=y�'=R����"�[�<�vf��'<(ͨ�dn8={~�ks�<�K���<azc<�v=�5=o9=m��Ҽ�~0=o�=�&1=��<��6���;J����=��&=���<q��;e�̻%6ֻ?�s��ϭ�dvf����������<�<=Ѕ<�}=��<�A=J/�:�3=�Z]=����+<�Ա;4��(����A�<���D�8�n��<��m��>�����C�[�v�<�{=2j+�&=?����<U��z�ȻY�<��ʼ��W�5C����=X�d<s��;*=�;`�=95Ѽ��?(�;�ӣ<=�7<��=���Un�B������<Z��;��<k=%�6�<��=#OM����rh5���=�>��.�$<�c7<���
�7
T���t�H�������wǓ���J=��'��9<��=td�Mۼ#�+=�t=�7=}��;�{ż�a:��>����<|�p<$.O<a�<�=���-���E!:=�V><� �IF��l[�fu0<.;.��<�4���W;Um�;�$9�
J�;�a���2/=l��<��q#�zb=�*��.:=����t`=�Ƽԥ�|�=e�#=�d�b1�<jl�Bj�< �n={]=t'�;(���03=�rR�Oڃ���;b3�l9�<LdF=cz$=�;�'=.�ɼN �6=���3=�$=�e8<�b��씼i�2��;W�< �Q=�ځ=�K8�������R�=��	<wʁ�&P�,�b�
�R<�ᄺ�²;x�ټ۠E�ِ�<��B=��O=�!��lj�=cN=�P<l�)���G����<�l������$;x�H�rQy<�N-�b�t=�0.=�ț���"<a��<#�<���^=%=ՁK��'�7��<~ �O���D	=)W=�mH����<�@���D��>_=�=�����H<nD�<����v%�8T��p�A���p=�<y�i���37�;U��� ��0�)~�9����� a<5?��v�=�&=yo�<0�<��$���<�sD;ͼ6=�- �#˅<i�I<o&�0Q���D�<���;�>="O����C=P&���}="��<�	���<v�<0��ϖ<�����<�Y���(<g=�q=iS#��&=iJ�z��Р�<���<���1BZ=z>��4��I��>�:=�
=��<q�=K&ּ�1��D>��V�^�o=Xb"=L i��m3��E�G�_=U����(�W[@�xű;�V�<o=�o�;ʶ�<Dj=�Zu�<1��*�*�yP=T=+t��T��rC����, =�;��
=���]h�<��绋!c<�:�9X!n=�*�f�׼��m=۝��ϪӼz��<�p<=��uj��D��)��FI�d��<|��<�a,��;�<k�#�h�3�|@B=)~�<;a�NX!��	�*�?=�nU�����ټ+7����S=c%<���j2�<6���Ǽ��f������v��6ݻ9�=�Z�<��c�ȹ�ڍ?�����K��	�<���:���:���<Wv��b�<�Y&=��C=�=��h<�2����<�;xʩ�`��<��&==҃�V�\=�`:�%_�P�p�"�T��y@�
�����ʻ���� =hrw=Jq8=����ڼ��;��j<��;��T���K���x���ܡ��7�;W)T�+����ּ��=�μ+V�W}ּe�0��%���1�<���.I���<�k���_=G����ѹ{��<�l��e�<S�L=��
=s�h=��6��m��F�=�{�����<�Z��*7��<��T�h=iÔ<Ix���<�O�<(VR=j/�<(nP�GD�;/<���<n�U�I�=#�J��9N�7@��!���~=��=�D�<J����f��<��t����<�k2��=8�ŻZ2��T缮j^=�I�3�=�:��r='�����1��n=)Z4={2<��;���;��=�ɀ<�Tۼi�'��'��M~亚nP=��)=��=Fg����-=��(= =*>3=��¼+�-�~�<e.��B�����Y���J=���;�) ���r=��<��ҼaDv�kߖ<&K=��ü�bC=^(���P�<���#��;��B=8�c=!{Ǽ�h�<	��9"�¼�h<��,<q$����<}Ao=8Q����V�<.��<��Y�`Sl<�<"���<��R�Ԯ�Ȃ�;�35=�5�9h��V�
�V�l<�&��@�V<0��='=��b�ϡ伜�s�8=��N=�c=E��B���&�<���<\�U=�ټ���<��
�JI�B=�⼧�<1���F/�����K�)���?� �<|�������\@�9�=䓞<��?=��n��޼h�(<��p=(9t�:���!!��r,=��м��X=�C2���%��7=9�B=�j���� =K#=�B&<M��݋3�ND�<G�c��=RJڼ:�X=�s�<n�<9o����=���<�~�X��� =�ao���s�����Z�<}(B��3�s�<ƽH��v��z}��m=5�'={��<��Ⱥ��A��;�~,=A�=$�4��E6=�P<�9C=�!�<�<_�%=�Aa=��;T�=��żP/P�
��<�_�e�غ��Y=%|�?��;��=S]C=|fs=}�9^3=�0�H.p=�2�<�$=DH=��/�jd�;l��=��K��VQ��`=�C)=���<�a<�3�-�=��=X%=��W<83g�!���*��gϼ?8=x5=ݫ���:Z"Ի�0��R�KX����= ����5;��<zh[<5�W�DE =��;����<��+YX���&=����ao�&4�T�<{V�<��<}�3��@�;�:�� =�E0�d�T��f��Kg��{<.�ۼc�Ag��]�</�"��4D=_pC=y�u�~�,�ք���g=~V1=��~�` Y=x�ռ�V�;׎��Kּ&jz��oS=m�fU=����\�3=�5g<D G� 7�<{8�Y4��o6��t����<J�X��jw=��	<��L=ǙB=�u<�yJ�P��H_��>=�C�Ȼ�6|0=�)=��<����@��<hغgO=�=����R�;G��=O��Zk���v���=�'<L�e:�̼M�&<��<~� }����6<�JM�T<y���II������<+ܙ:�4=��J<׺E=|�ѼG2s����<�=�޼_}�;I1]�L�|��(,<�ag=]�����j�����ʼ��`=���tد<�i<4�W�t�(�PC=e�3=�!�;��N����<_�<:���݀���	�y�?�U<�^C��[<$�<���;-�m�b�m=�#:����<�fE=�|,=�"�9+N�=~!=`l=�jg=�T�q�P<_�ּ϶:&:=5�;=�"ؼ��K2�K2�;��
��4K��e<�,Q���<�7[=y$=R��<�ػ�)0��?"����<"� =�=-�^=�A$=�=�sv<�����|�R�u���
=�'�<Hu�<s&=,œ<���/�=̻S�8��<D��ܓ�H =���=&�]���6=������\�|)��>}1=L�="+=%�B=�^뼁��U�2�b:<�a�]3��pݻ;���ͼژ�q�	��(
�	<_�����=��o=Y�=�$a�O�<#�P��;&=~�<87=���?�i=���<��=W��<��ƼhVB��h�R��;@=�J)=�Ȳ<�I��p����<;{0�;3!�X�<�L<T�=�V=M�==&3�<��ּ�LH<6��L:�n����g�<V�ռ�Q=(�ۻjX<��R��	��=����J�=l�<gp��Q=ii�<���I�������nM��E��
�D=;q|=���<JC����h���څ<A�;��p�2���R;@� =)8=����`/N����!�f��?%=�=�if�|j=iO�:���:�<�R�U՟<���;e�<ͳj�.�<4�i=*���	=���_<I�=��<�˼?ƶ< �ļ�mT�[�;e%0�[7ż�@;˨��&i�f��<QY<�f;,@��.i�<�>�.�B��pĺŀ�$w��)"=l�<��-X=4��;�$v����fK��b=;4�<�h�<�B���|	�T�<ԇ弼��#=��R?<e$���^I��I��[������=)�<j����;��<�ő��n�;��!=@���O���F����T*��^@��M����!=��5���&<����TS<�X,���=�	<�K=-Y2<��,�<�,L=-����=���:>lQ�sex�B�=�cJ���7=�]6=e�3��N�bCμʻam���_��Zi��9�<4=��=�	��&h�1���"-�3	�<>A+��O�����"ߑ���<���s�o>\�����I�	�KX:�?O;r�?�QG��Ɠ-=}�����=e�	=n:r��+=���<@k'=d/�<��@=rba��-ƼJ#m=8\5��u��i=뉦���Z=d�)�=o���~k=G�t��fT��FG=9`��9���X��5<լ�<3H =B�_�nk�(�d=�K�CM ��A�^z2=P<���?=�H�S�B�mzʼ𕟼���<�1;�э=�=�Yb<�s��3��d��;P�d=&���De=BB<GӼ��x�L㍼��l=���;Oa���U煻9,��e;�[{=`=6����;�f5=0�@����=�V�͉��pF�<��;P%I;0�u<��ԼN�;=^�<W�w�����b���;�0L=��W<O-=�N֥<0D;e�f��"=���;�¼�t=V�'<�l,�;=�;wD&=T�<�}�;8x���F<��0;�f��<k�����;!Ė<d(�@4<�}y�r?'��z<l�+<�jR�t%y<�}5<��)�E�$�<:*&<e���-k�=g�q���<���<���=k�e=mP�y2B����������U���p=\�\<Т��`�X�qN=�8�;#=>�3<��o���<B�_��LK=��=��e=��F<�	J��r��������[<�r���	Y��8�<̒#=ԯV=�q����O=la@�>��;��<l̅<�v���}\=#+F�Ǻ*�~�~�>�;�3�wr=��<��C��	0<��|�^靺Q��<�Zq;7�J�2GS��5��Z̹�Ô�NF�;P��<�q��K=�t���#�L�<{�.=�^�<�D];�{<����d=]���b�<��G=����W��� ��<߁��멼���
�Ӽ�N�<��B7��μuQ����O�>=8O=臻;��3���;(���+~�P�<G��<���T�D�T� <oo[�H0ȼ��E�ǻZ��q)=�-=p|"=��a�Rļ�.��0Ҽ�==�-�'�>��Gm�33o<8&��M��<BX���(��^ݼ���1�<��5=jA@;� �<:��z�<\��;49��4�޼�<��V�2",<�L�</_\=ō����<�ü>�;؏�<�N �W]=��縼��?��)J=��N��,?����<�h��6�x���=;�S�Ι=y<y^��b�:8�ݼ;+u�����N=�E=~��<)K;��`���h�eQl��K*<^�m=f/�T�4ux<�LF�p�<�q=칎:bi�5����E�<����ϥ�0�%�����NS�
�мc�B=�]�q��<�61�b��7=���g��f�Z=��n���;��<o\�����e����<��<A�_<t�==qT�E����<��&=B�|������=M�)�p��b+�<V=�l�r�8�0������甼�d���[��w׼��G/=�=�z���(S���Q��G1=ו�<үx<��n��6=ڷ��&-���2�Pq=��C��&"=�I��uP��E@<�ǉ���)�h|��x=r&d���Q���h=�nX=�佺���B=��7�;�=�VI=�VM<���<��;/E =���<��+<N���1<��<j�H��,#=�;#S=%d^=��Y<�A0�����⩒;-�q<�헼�(��7�����~��Tϼ���U�=��Z�� H=���J�t�!<�3ټ�Z�K��HhQ�o*Ӽ�g7=|��J���VR���;�T9�_�$����<ྯ��0�P����=�w2=��`��qW;��~��=H�<^�l<�U`=S��Lx��d��i\��(#=�k`����� �5M~;<)2�ʸ'�J�&=v=�U�<yf=�X4=;�1p<��<=e�<A�<��=�>�W�<�8=���=̲�{"��.�<)��������)=>�ü��a��R=J?=*J�:�<�<�S/=�6p��^»�}�<z�3�a�;�����&=?�ϼl���[�e�F�έJ=g�}�: �d<w�<�<���s�<ѽ<O땼�Z߼e��T��<{l�<C�Ѽ�/W�o-ټp/b���M=dU==�YU=IH�<��?���q�6La=�tY=�E��-1)=�V�:V�<=(��/��D>��~��z�P���<<]�;}�<�h��x�O�P@�/΁�pU;<����4�f�<
��<��?=@����.�A�<��w=�����u���e�$�=��9��ӆ<=v%=���0��!�=Yn�=Q���i|���=�%�<Y�C=�k��О=��S=NF=%�	=��I�L�9�����
�<��<�38=̄��U=��=�>�<�
���2��'��b�<�1��#F=��E=��P��Rȹ��;K��>�v��N�v�U<[у=Nbh�����6t;� �NW��0z<]xt<��="=d�</Ys�4e8<b�i�<�<Bj���c=�L�:�LD���Ig�;����1&�Nλ}j��c<�L�5�м+�<�����=���f��<"%�;i��<7D��f��L<5� �E�<C��<�	�cź�������s[C�� �NK=��F�����$�<`�i����L�:���@=��Ǽ����G���H��SX�<�gF=H*t��6�����< w��w8�����B�Q"=V�.<W�K����<�W����ʊ[���W�d�[T=�p��*�<zc��j�9@���g�:�ϼ��N=`п;t/����Հv=���<]�M�I>��Z�μn����(�+��3�j=�Ŋ<+6�W'#�98����'=�𼯊E=���;F@<�=p�ͼ�,C�!Zϼ�`c<�H��s�=�F:�=���<l���*��6={�]<|�#=Jwc����;
&�<�tͼ��<��^=B��<�(�<m�!�Y�~=��F�o�6��׊<��b=@޼3!��5���+=��N�m.��I=���B��<ٚ7<֨=��G����;e��a)O=�|(��T�<*wi=d�Y=	(e=-�X���Q=�=�=�*K��l�Ѽ�UM�PҌ��7=C��<�=|3�<*��\��!<�^<m��ԯ.<�&�0)t=};6=u<gv6=�W����<=���<�5���P��j<��）=�r����W��Lk��=H�<�fY5=�0<`�����i�d�=�!��;���i����
=�3=���Q�<Db�$:���Ѽ�<��@��uT�Q�=��<�s=w�>�r�<ڑ�/�w��n��C =��V=�bb=G�;~M�<�� =1�=M�7=��0���<�z=q� <�+F=��<�<1��[���x�#1�p�<�ؼ%�.=<�7��	�|�U=�T��W���زi�+�<Z�;4�����<�zW���<� =�=�)fU<�<��I;T�!=����*���_`���y�*Ӧ��:%=�+&=t��qh�<�7�<΂9�3%�;G���k=�=v,=�pM=��w����PF����=�g �82x��b�O�;<��=�&n�B�;E; =&IO�����<�6�� �	��t��������<c|{��;�V����2=4`�c(z<3�r����+��ż�����<��G:��Z��2h�uY(=�*�~X<�	=���<�2M��x��@0K=��p�(�<��%=&�4�a��"d�����<�Z	�Qs=��d�6�c��>�k	�<S�L�NQ
=O��<���PD����;�$)�n������<�F
=v�<��=�A��_�=l�#�iž��DL�|#�Y㼼}Z���<dh=,K==�yi=�R ���R�=(����T�Κ<x=Je=��A=��:=�Sż5�=Z�_�0����<=i? =��˼=��?= :6�*=\�[=�Z=^�;B�����{G��.�����<���(���9�<>2M��M=��j2�t�ż��d=��A����<Z0 =�b=θ=,�P��*�<K��L7 �J�C�U�:C@="r=��%�Z:N�4�=)�i=mI�;X26<������ =��:�ˎ;}��"�V=DW��V�$2��
�{���l=H]2=�T<��<���<��;�䊼|ST��{�<�&<��;������*��nM=�NP�}����<���<ݶ"=Զ����%<���;-�;0�=�z޼�W������<\5˻�'�<x,<ݎ_=Ȥ�</$��'
����_��s�L=�g>=�O=@�1�B��*�a=ȷ<ה�X��,�%=s *�$t����\�O5�<��<��u=��Q�C��<�[C�24q:���;�8<�@7�i�/=�[�;��%�����Q$��
�:��*���<���~���n�l�f�@��<hkj<Y�T=@�o��I:;^�Ի�=̖Ǽ��=!��B�L=0�<=ߦ����~r�<
�.=���<�z����'�y!�<݁�=a=���#�;�w���6����F����<��~��h���;�-U<U�)�	�)���-<fv����K=�z�z)L<�=Z�
�f�=c��K��\�8���<|�6=�^��ط���J=4=B׼�d�<V��5���F=�7=T��08�<�[�r�_��g5��Q=d&i�4�=,�=:���M?��������d�;D��̙��f��А���<�ü{k=��=��<Pk�U���RXۼE6�<]!ռR�c�)�H��K%<1��<�Oݼ�t<��8E=a����Ó�t2�;�9��=�9-��W�Ogj=~3*��²;t$<2�2<��#�{B=$�]��x��$��<&J7=�~J=��2=/�Ѽ��K=��<sF=�Z��Lܻ�*4=,�Z��	0�L�=(���
=�w����<vY=�ْ=SDL�"���%�
�n5�;�R��$=��=='��It;<��<�4����<������<���Fb-���g=�<ԹD%6�>V.���~��P)��e=�{A=4������=�M���U��z�e��-�<(h<�i���vd����<������ҼS�Ѽ���P=1=%�=f�=�o��a�<%]��l��<	酼[=��G=�^:�7u��ț4=QJ�BZH<Nn(=��=e�	�+y���������}�ػ�D�<C�?�X��A�H�ؖR��3 = 1S��mD���O���e=`*�C k�5%��S/.��:� �;�܇�Q���B�\���������<���:"�<N@	����=��W=�#=�B��k:?�R�=��*=��=�o�:��J<V�D=t��ļ_�_==�P��WI=}%�<u==�
E�P�<�\�a�����<��=�T�<F����P��~F=����R�5���=�b��[� A=	���<ܕ=U���z����?4��J0j��͝��X=�G�<�NU�� �;��=���<�U�=^R��*��%*:� =^�<P!=P^5=���w����Y��a��U'B=�,`���<z�;J
<�ۺ�� I=���;�@���I:���<4�d=Ai�ơ�<wH���)����=�6�<ٗ=2���m��J�{= U.���_��xJ�c��<U��w����s]�؋߼�D�:E:\�����	*=,��O塻w���}Pn<���<�7�������19Z�;p��<�����;(�<=˘�;~],=L���n�w(5<�j=<}��P3=�_:�(tm<��򼱁==\�:<��r�͵j��^�?0�-�.=@rc=���<��E=�<�wȼg�����,��:����^��3=gh'��q��#G���V<��,=U�м|�=��Q,�;}�S<��+<#=��L=�M�:��u��>(�<p��<ᇐ=
��;�x���1=�l�}�<ɽ�<��C=�E=�ŋ:����r��^�A{��3�q=|XI�� ��z�B����<�n=��V�jRv<h����߼��i=�A�<+�=ax<E�)��CI���K=r/=�U��=���<zD;��lo=_�Z��~D�ihX�=3Z���<	=�)<K=��6=ԊL<Gy+�U����=��: ��<�ټ[���༪>=Od<����s=�8<Λ/��!=6��;��b�H9���o=}�<�=EP��< �``}��!E<l�n���*�=�C�js="�|==J�.�;
-=�l�<Z��<��%�|WX�x�=�y�<�}=��h=il]=��_��-�<Sa�vc�<Թ�<@J=$z|���'=�^=���;�p��Yi0=�i���4�ݴn���.�Xu��P*�BUg��Rx;uv���r��`�<Q\��D���&���J�x! 9qź^��<ٍ<�R=+�<Ŕ�#����l[<�ޝ<|O<�Hջ� 4=����r�b�1F�</E������;���<�5?<���<6u��q�<��@���$��Q�<g�_�,=n�1=Dͧ< ��<m�=�l�<�Ѽ̐^�'$=�b�<��E�lS��[F��0=$yT��?0=E3���9%A�;�<,P�<&�==[e�<ق�z�t=�f=�"���K�qֻ�P%�_�9�W|Q<ҾK�Q!<�U���7=�r<��<Q�=��}=��+���?<�!:�<�8��G���r�<���=�܄<��<��>�c�Z�>�R�b���n�e=AN�<$=z\x��־�L�j;c�s��9X�*'�<�/<sL���6=�M=$-F=�ȼRo<����ǥ<�\=�:[��O
=J:";cM�����������;S�j�fy�=p�P=�g�9^V=�#�5�N=�$=�(B��ie<m�<R�.=J��o�<P<=��i���L=�I<���;> �<�u��+�v��:';���=�<`z��wJ�Ѽ�i<��O,=���<5���-��a.��t��`�<�5��\T=��=@�W��+=��9=!+�<r�˼��=b�L���z�X�<����#;��7��2�qW���)=��<&A�<�m$�mM�<�f����;t^Q�έG=B���i|":�<�H=�0<H"o���+;y*ǼNVH=���Zf=�?=�<G�H=�O���Ax���F:?�@=1�_=3�^<� �:�e�;Y_y<�25=k��<��;�Y1��3L��-;�6�<�nټߔ`���d=� ռ��,=�ܼRn�<^�H=z���[?`�j@�i2�<<`�;�,=��I{.<�|���\=n=�5��E�<��M;�{s����;ȭu<��7<G�<O���{<�����B��I�*<έ��n��5��q����Y=����h!���	<🻮�<�t={���������ش����g�Ά˼6��<y�=�刼��G=���D]��ǟ=Tv�<�2�R�9�Tb7<҅j�}"�;��g=W]=y���ّ��O�3��lJ=n�=5`J<�PZ=��<�,6�mͼ1��<�s���*�9��IF=.�;�Ӻ���p�e�5��qy<�&2=ӧ�<��8�Dq�W"�<+H9S�N��� =N$�=�5=|ܗ<"�;!�=���$��<EsB�a�m=��^�oVC=4sQ;��5���U=�}	=��L=��G=�W�:��ż<W=��E�K�<�X=�g=�P�#�	;�3�����<Sg=����34<��ۼ돰<̺��<��-;Hh<�G=7��<'4T=�!��ϑ�kw�<��C=�*����;�!�<Y���lp<5$�<��
���'=M��<�����/==(�2�K�J��.=�^Ƽ��	�L�-�!Z!=���M�ͼ�w�<�R=�����6�~G��5��}�Y\�<��=� �<��ۯ���Jk=�m�<��(����>�O= ��<f��<�7C��nҼ�[f���U=WﻼR�-�K^�Cc�;���;@2=~_��NF����Ah��5Փ<��C�6�>=z�+����������2�QMW���ɼ`0�<W�!�4;���j��;L���G=��9��ȼ{�*A6���`=g1�O//�G-�;#K=�Il�S)3<P�S=������d�u��Έ<�C@���:�H�<�,J={�6=O����=	4<xN����%���#���;Q7��oY���l#�Ld�<��=�J=���<ph��YƼ����}><_<��A��ƨ-=o5�ɔ����������<�4�����;������&���e=0���T).=߰3=>+�;V�����j���v�ج<�l��l�L�|�7=d�V��7 ���ռ���<i�P���;�j=��C+=K� ��:=�;�=���VB=�4����b.=fl׼H��;��.�ǐ�<DE�=��:m���p޼�6=�@�-�9:1Rü�(���υ���m�I�z���<��{<ڗl=�M�<A[)��c&=O��=�m@:k=�F#=�b��\��rz<ZM�<��=K�ؼ��:�gp�|�<�"�<�Z��Hf�a=���x#=KA=R�=�9'� �Q�D�G�L���|;HB�]�����BM��'��_=x#��J�<��|���4=�x<�x�-�a=,Q�<��N�Խ�<V��t�=�6����Q=B=�}{;p়���r�ͼ��N=����9I=�����<�B�7�;��8����%΀;�;�W�9=3L%<D�N�"7=H�V<�;�<+�����8�(=T�K�dt�<=��<fXD�˨|���V����<] <��Z=���eH�<,%=��\=��9=��8�#O�;"��)��ż)��<'=b���6=�WR���<��V�p�<����$<��ݼuk���gD��e=�ͼ,�_9<��<�Y�Lf&;6��k�4���RE=�����j=q#>=e�2=��<���-�=�k&=��A=
㮼�H��P�Z�<��<�\�?�>�t=���<9=��<֬=2�;�-ûTl��'U=�=�\Y=�ʝ��Wa���=����ZNQ�xS�<'��<m��g��<k̷���Z�+��<�����:��<y<D�L=���2�<���R��<�`���m����<��=w�l=��'���z<���ea
=���9��Ȼ�~<O�<,�b=��л/R���*���3=FV="b\=L��<b��<�1D<=n�<pg<]ѻ��ü�b�<�:�<q�� x =^�<	�ʼ�y#��=�:'�K=E�!����<�>����i�S=:��<��[=�Q���8=�鼡|%=4�R={m@=X�^�z�=�]ؼIA(=囡<0SҼ�H����K�W<���<�oG=�G�������<��'��'���<���<1o=@R�<	��;��<F8m=�;F��<����.���<�V>��!=����
��<)��<ej=Дm;�v=�8n�^���,X��ʼ�y����O=�~�;%(���9��@�3�����mf;=�1�Íּ�=�<̲��G���[����9��<�E}<��
=0�<����J=��<bL�<b���A8��d&=ʏ�<�����<QL�<�=��%������;_h����=l�<�k�;�Ћ;Q�Y=@4J�V��<Lr�և�;�!��>��<ۼ.�A=��=�Y�������<53��
"�K������<��3�!��sF=�o>=C����h�;$3�QR�:��T=�ú�����p�7=9�G=�G��K	�]�"=�h@<Ë�� =E�5�,���Ҽ���<9�<��<����<a޼��;=4ٲ<�g;��'�Q�(�Hy)=SN2=�����<Ϊ��ь�>�<Ӳ@=:O�<����A��A���7��<���=i�=���r�<t(G=���<��r=ۨ�<R�<�<=�&f�̑4=��=��h������3�H�{=gI<
.&=)��^M<�H�<�>��é:=��<�A�_�>�ǫX<N�E=�;��}f�`D�<9~8<�����<}��<����=X� ���`:���V��<su=�������b�ü��c=D*9���O�����]F�T �<�`�;�W=������)\�<��\�� 2�9g$�Nz߼X���R��eR�<~�i=�ߩ�2C����4�_ ���F<+$/;B'��,�W�0q�;�C�GB=`+F=t@лX��qb=�\�d��z=]��;!�⼧3=�"��8�<����j�=���4��a�=���<��O�G�
=p�ں^�O=���\��9�5S<b���J)��
=��Ѽ1}d<��<Yh�<�Ae=��μ9����V
=�Y�O�H<���<q/��|����-���Y����yO�<Z���>__�2�8=��=�ټ�Ԥ<f��<+��2=�@:�*�<��h)�??�;
o�Ǎ�<��<.�)=��!���<;:μ>���S�<w��ϼrO�<�-��;�,���#=}Z�dF��-��+(�����G'u�](�<�xr=�W =�Vͻ��!;.lY;c�=l�.���(��v��:C������cH�;�X�<]a_=��(�N�<a:(=@2=L	�˼��-J=�;K��<�݊�����=���tB<��5��	O�7F���ѽ�����o]<�\һ�ݼ܌M=�s0=���v��;�:�g�5=��=�S<�U�u)<;R�<�`�Ff=X�<~F�:�Z;2v�<A�	�h�X����<MT�< ����<��<���� eS=�Z�<���<0l<��s����I;��4�<��4��y��`�;� #��F��*;7=�Q�	��R��n^�ƐZ=��4��+�;�ռ�â�,�H���ҼH<.��&<Ϩ�;i�c�`�"<���<��Y=ߔ3�,?K=Ԏh�x�B=m�G=ʔ<d����i=��s���]=�
5=�O,�G����9+�;=��;g��;�/�C�<#��$�"=Ӕ�����<�<S��<�B:m0�=��F==�����-;� ����sv��R��\�=��)=`ԕ< M/�1=lQ%=��Ǽ�H�:v�G�"�:�_�9��ߔ<غ���KL=V�O�~��;�,=v "=7)�<�M$�Th�:.~����d�=�������<��^���A=�Q:����b=ΕJ<��#<gE�ʪ=�.'��t+��CY=s+=stμO�1�LI����<�q<�;�<�:=4IҼ���J_:<��=�$=��c���f<���ڌ޻��Q��-h�F��<��<N�Y<���<ej{<R�\=��!<���<��F=�-��ځ���v��3�;�zT=7��Q�%=�	@�.�;P�\=6�ּ��*<w�$<�N��4= 9�=��=��r��ɼ%诼��M���8���<�/=�����
�LbּX�<�r��'��ST�<�	=hZ�<jI��.�`9�:_I;n#�<Ť&���ٻR߻���Ƽ���������;�ݫ��~��>=���<�F�<�N��;Q^��VҼ��=�p<�$��ex�<���JC=s�-=�!V�u��<��%;d�G=K+h�{�:=j�����<��2=�Y�<kT�;�Τ<��Y<��	����;?D��k-=>*�;Z�=���u�="�@��CD��d���Vļ�R�����/v=�"':ߕ���`}���=�vO=�N����S�a=a^=oQ�<:D=]�����W�	�
z�y�)=�<s"=ʄ�=i�E��^�?+f�����̼��K�v18��Cϼ�)�����;T�<�.=A�=8���.=�O==瀀��.l=|e{��_�����<S�(�4�������<詼h]<�P���x<*���*��Rֻ�U��X��<�m�;�p=��=J� =���x���ͺ6+�<f����jq=w6;U�=��#=(�~<��;�GǼ��F�D=�NG=B:=��:Ry;<�*R=�?C��X�<wm=ʄ�<�խ<L�伢ݸ<z2�<Np=��-�pS<�=�;C�[�ȼ��~��<��>=�v�� =��;��!-=z�H=Ԁ���@=F�=�bĻ� = ?꼮h��q��!�����qv<����,=��~<�(���1�*Fռ/�=]��;}`��fs=[4O<�hG�g_��٧=���bl� �+�u��<U��;�f=�>���=�v<L�m�A=��=��I<�A�ǰK���y�O�;��_���"=���7���F=[��<��<��ȼ��)�WU=���<	����b�<��;�[��}�i<I�.=�3)����� <�^3��Y�.�I=���<��!=��F�wɼ�.,�<H=��=[�̼3&��j�ü��=�jh�����H=��?�ĸ"��s"���<���<L�J=��<��B=9>:*w <�#=�3C���>=P1S<��H�P�Y��-��1��;�<��2=���<��=��T�0$l=p10�pN��b=�{<G`�=¤=	SD���Y�^ ��Z�M=��
=���~�V�O��<6馻y}s<I�B=>{���A���8=�F<����/<=}Z�<�Ԕ=�<��z\���%�R`#=P��@��/ڳ<M�<��<]X7����<)됼�2˼ �y�͑��w<�i�5�Ҽ͕=J�<AO��"¼Z�M���c��{(=�n�<;5T<&d��
��=$*)�d�.�+:�<7��R!�.�d���*�ւb=��7=y�#=س1�����!=���<�T�<�C�<�� ��wF=���e7@�̤�<��x=�LB���>� �2�V�>�n=hL�;��j�/�޻�&ĻR���w-6��F�<�۷�7�=��=�=���OY���=�� =݊�<*���&���m=�=�;�'=�bh<�7μ�@<�8�<T6=�}ۼ�DI=���;��<] ��pݺ�h�<�J��b�
�<�%y<G�u)E=Oe�<�J�|�����'��!��Ku��"����O7�%纀�
�̍G<	�����,޼@:W�H�<��I��M�<9�@�����h�>�n<~��<���`�X��7G�3����3�Q
��y�<���=���̏[=�Z��6�<��n��� =V7=:��;��`=1@�<P���3q��_���2�+S�;z�`HܼW�D�Y�����i=4n��_l:��s���� ���8���c��/Qx<����1s�<��h=xAx�ɹ�<��!=aQ���i�"�⵷<����-�,*��.���B�H_<� �ѐ<��m��u=�>G�j,8<� H=m���7�N��	L=���<#�=�ю< �}����<�>=��^�C�]��&E=�@=��W�.u*���I=b�`�l�u=��;R5?�-�A����;=�<��1RM=�e4�3l;���w�"'�<K��<f���T�W<_���6��Ą�M+a=�LA=ėȼd�<B�&�p{E=,��}O{�#4�(���y漎w���m�PjH<5x�<^��<+�e�L�^��=��s��Dr�0�=�6Ҽ�Rc=G�l�AD
;�6P=n�ɼ��x��Y'=�����V�<�B<�x=�'��8=���h��<gf��|�.�� ռ����N�O:t��H�F�s��<L�n���'�<�M=��<:�Ǭ�W��<q�<��;�鑼M~&���;tB1�p ���=�M���w=��+���W<���<��żbtt9no��R���W=�r��P��<g�-����2ܼ���;;��[n�@ ���{�V��{^�.f���0�;W �:�G#��⋼M�7�a�<g6;��`=�!�>�:�G��y�<c�W=��Ȼ���#�Z=�<0�d/)��,,��Z�� �R����<� ��z=<d��,���S6<e4=.��9r1)���>=��Ѽa��<0��<H�7��FI�۱a=�<)Ax�{""���4=�E!<bV0�+�7�3� �&#h�7G��^�<��<=ģ���;P=�� =I��U�I��^鼤�û4=fL�;���H=2�]�B*��b7���.�Ra@=l�Z���?�?C�<vD�@�5=z���?�q�/K-�cA<$F���KO=�N<��=:3=}|��;HŻ��"���a<�4>�D|�}L�:\,��߹��7_=̨*��D= �� =ި¼�2߼?Ͽ<�!<�g=��1=f߽<�E=>���|�:S8��j@=�����;W=�M�<N�/��fk�1!�<�[=J��<�
C<�N�F!�<#/��˶s�f�0=*z3=�d�g�_��F�f�߼�;$=h��<^�<I��;�K�"Jt=s�f
�`H���`��	��;�����ͼ&�U-&=��=��A�}-;�#Z=,$�(��9B��<��!=#&C<�o*=c	"<3�y�X��<{7@�x=���;g�<+x��7�b���
p�3��=�� =u�ߺTB�<ծ4=<����<�߁<�[=[���D=R��<��=�c���*��i�*Sc<���<S6�7Z��%���^��� �V�=5D��Kkf;<�<6=H�U;m�<I�=>ۼ�@�idE����:��Y�G{A��v���k�/�ɼu��<�ϝ�"����&=�ŋ=�<�L<U�<۸���')�@0�9���t�n;��̼F}g<z��XT�<�B;��&�XǑ<M"_<PA=�9X<�:=�~�װ<��*�鼸��<��X��3=��>��O;C=*k���t="^�*��=�y6м�����J=WI�<�W���W���h�<�zv;#��� �;�B�$i@=&v�Cґ;^?t��]=�=kpB�aX��񸴼�c>���,=$�H=���<��<�P��<)�޼Bi�<��<�+><��<�k��E=�[+<�[#���\��qh�.�=~����b���+e=CW<�c�; 	=>e�� �]��zn��Id�JqW��[�-^��F��0�<�fܼІ=�ｼ�l3�b3=���<�8^��M�(�=��D=�0=�(<,7�<�l�<���<a�<=E����8���X=iI�<ܯ�<���ϯ#=ş���<�9=e�_��M;�����<J"�<d���{p=2�`��� ��c��|�=5μ<��<)e*=�ǻO 4��]=:v�<>^�;6����&���]9��<��*��<*x;�&���խ;��P���<��n�Ś���6"�`�
=!Y����Zy=�bc�<O��<#���3���RF=��q3=���xj='�<��W=��6<�a=6z�x�G<�<�Q=#�=�F=yL�:�6=��#���o�T�s�CyA���4<�*g=~	=�=���"=���<�l�n�S�MX=��<=&䃻5��<�jR=C� �J �<�G��;��>j=���R�N�1FQ=�Q%=!<�<�7���{���(=���ъ���"=��F<���<�-ۼ,�C=%���	=���=�^���M=��ܼ�ѝ<_�.�c�ܼ�\D��*�Ⱦ������{F�@[��L�W=f��<3A�� k�e
�>
=Az�&i'�>�H���׹ü]E=��P�� =�I�iټ�B<�^ ���<���<���<oBr=³���!�0n=���%=� �<�b=ڒ=v_�<1�Y=�U��(���伣3=�?&�=li���k<����!=0|��L;8��qu�����pm=��B�#�=b�ȼz9=�!�A�ʼ�J���=C�<��f=�����њ<�9Ua��^�<x*�8R�;����;穳�[�F����<��깇o��S�<J�=��ֻ,^^��=��<��m�e��M����;	�< �Y=���A�r�_�D���	�<��<�`;�/@������%漝v@=r�f=f <wq�<y�+��WI=~8���8�������=��H�I<�-�2�E;�vI<���<�V:<�I,��ϼ۴=nP=͝���y<�ༀ�L<��v=��=A�V�!9���
�%��+��Fp��x��
�;��A=�5j=��=%Sڼ�x���.~���|���z�Դ�<N���c�)=��=%�=��<��8=�}i���=<:�'=��e=��N=�/���39E�:`��=6<qȢ��밼S7i;oS��c��c`k=L�8�ğ�:�ג<�=�6<��=��<�uy<�_7��'=x�<� ?��}F�DI<[�2��[>=dXݼM���=��;<�V�lY�J	r�]T�3:��c�;aɾ<3l=���F{#=��>=C���\�O;�<;�!o?��(����{=�/D<�dC�g�=�K�������2<�+<C�9=LT<܅h=��R<BJ=Ԟ޼����<�v=ՙ�<�Np� ���=5�e= ? =�3�<pk�:����a�2;΅�<4�<F�!���=��,=�9���(4<^ƼJ���<�=�N����^3i=��=H<�<=ܯ�>�j�*�U#=���ۘP���`<��$�s��<�����<$�=�X=]�;I=��={?�Nt��>h���L=u1x;��C���#�����^E����<tG6<&J��)O�=&�(��=u�F=u��;��\�n�ڼڟ���==6����y�\<Jl�<�Mo�3�Q=}cX�!�4�k��n���H���5=T�d=���<���4�=V٪�� �<&1�Yi;��<��X��'M-���
;=?_�<�ˊ���D�ɂ=�=7�6X.=���<k�<���;M�,��<݃C�QἮ�0=�p�:`�����,�:C8=Ev�v���/<nY=�!��of��v/�|{3=���;K�!=�:{;���
l�SO=6&�<�����S=FF=%}�;&�R�$�Լ��\��ԗ<�|�<hG"���=y��<�E�<{��,=z�Ź}�[=�&F��$����<&��d�=l؁<�C���I=�dj�ʣ'��9=�/<��<	��� %���=�NN�y=6=��i�s���
��-<K,���vM=�\(=,�Q=�&=�BF�*�+=y�@=�
d=3{5=d`?=�=�}K�4ć=L]<��u2�c�<�	��C/�<�\��2�?<������;�Ss=7���0=��;��0`�<��=�u8=�j��yP�<�2=Ŷ=/N=��=Yɶ;M2O��?	=�����+��u�<t�&=O)��m�=<�a=��Լ v=k�%�>��g��d2�:�ڼ�B���=U���X������>x�<;Hy��z��3"����KL��qK=��<�<�No=��=��O��l=$%=���=�梼d�F<��=�Q�Y��<	+���+=�Q�^5G=��켥am=Fx��s
�o�� 9�<�C
=E�(=d�=|r�< SD=Sn�<�$9�uqU=dO=��/=��G��I�<U<ָ��N�3:W� v�=�vU��*o<V�U�,J���<r5�]��Y`=�
���*=*=ق�Id�ҷ�<}v�C��<(h��8�c<A�J���X��P��	��#�<Ȍ���	����4���� ��}üQ'S��<v=���dp��Fg�k�|�?��ը)�� Q:��R��<� ��u=�m���+���SǼȤu�E�B���U��N�<9�伟�U=�i�y��<`ɻ��h����s/a=�����S=��<���:��;� �<oq���=���<Ӏ�
�2��м9W���gO����H���N=?��;:e���<T퉼�ʩ��ꬻb�7�Y��5#f�0�q=ҔP��1��'=��������Q�<$\,=c7O����<EW=a]=9q(�B��<J� =�D�<(d���<�"�<��<v,=nr���$�<�c=�b�=.~���D<��"���<w�=�j����%����6�<Q^�<zj�m�P=�A_= s%=A�<.�X=[�м�ܼJ����=��<�u[�>B��&J<dY=� ,<���<���<�X����u9y=��ƻjG��)��q�=/�����5=8�=���ܼ���$,T����<�ޓ��唼kɋ<�-+����������0<>�G��0�<Md=bq<��=���;*����~���=/z�a�6=E�����x<�9<��=\\=s�7=��<�)i�O;"�2�Jc<P��<K��	��a����/�t�u��<�����]=���nG=�0���p�:�<�P�^꼂f�U�!���!��Je=���V�	|�<B\�p�,=�|м�ӄ���=��t=�%�;�{;����`=į%<�E_=� ����Ҽ R =�Z���<`/O:���� l/��L;�m�<_�;=5@=�b�r��=�W����NS�<���;6��:;C	��:��?�?o3�� =�#$�n��;H?+���J=�-�����R��>;�d=~�컨�Y:Rm=�U�f���<r4��mV��]B=��&�a���<>#�\T=��iܙ��v�<";�n���� ��d<�{;�QܼGv�<��J�Yʃ=݇j=Z%μ�^<�6a�3P(=��g=*ԼX��Ȟ=���*�ؼx�X�C5��4<(�<�P��V�<�ȼ7㎼���<��3�p�Z��<�{����1=���<h�<��<�U'm=x� ;�MU=� e;��I=0΀�mZ�<}#���'=>�c=��t��#=T��Ӓ��0=�3w��Z�<�輑��<��!�=>��<�T�<�\�<@;K���q��u%�w����Y޼�����	=�n�<�I�)����*��)�:���1��x�'<�q{=�ň�"�W�L�1=��f=%5;�#�R��F)��$]=�^>=O��<sF���P9�:�<랬<�B<�b�<�ߛ�d%F���w��|�������F�K�<dp=-�X���;��B!==#��7�b�tB=�==�Ӽw�(=N�<m�S=2�=�v3���;�ԇ;"�+=˸&�E�H�@���H�Լ���;N�����;U��<&,ϼH~$�=U�M}�<������<*��<�i�<�q�� ��[yA=��^���>=�f��뗼����Dt4��-�¡�<m��&r���z&=�գ�f���ή<�UN���0=4)=)"�<��[=)=����i/ü]��<��5�ϗ=1Kۼ��E�]�^��J���`h9͐;|fD���:�=2��<�l����<�b�ZD2=�y:�E���Au<��1����<�GA�*T�
o@�%_D�/mX���x�#׹���P�1�"=h�j��.�<���<�-�������6�<�r���b\=��;� �;�_���7=�62����;D��<wT�=B=$Q����=ױ[=	=ζ�;,�c���=�I,�6JK<b������<��&=��IMP���@=���U��|F���2=���<��<�0�rg�%��5�<+q�\�o�*C��΀;���-=��j���L�<�����K!��3="7=6C�r����I�;�#���Wȼڂ<C�,=Ȉ�;Ee�=rv�<M�S��Ed��j?�8ۇ�$Fռ3�O��<���[<�1���'��E<û/=]P&=L*<=Aն�.�<�A=a&=�BG=�f4���ǼE�8�̩�:�!O���;��"=�g��E[�h�-=�=�������qL�����B-=��9��#P�[׸�0��:IU���;�;�mW<,�a=�j;Ի*��V=���<�O>�w�;i�{���-��2����F=��;?e����=�Y�<�Q<��==�{��"}=9v>��w=�ʼt)t��憺xK5=�0�<#��<ƹ�Y<#�7��=�st=��h=Ԏ�<a���ˣ����B���<� ��X��/T�<���h<�I=l$���=��<;2b�<�l='��f�����<������/=�y
;q)h;�$��Y�B����<3�<�P���7=��<��*=���7N���`��(���
=��b���Q�F	=���<��E=V��<u�O<E2��b'��A�D=��A��ur��a <IF���ü��:��=[�'w�<	I뼎b��n.�g,=>$=1B����<S�=�c�<O�V=�#&����<1�+�|���H�;;��C"=������+.; I�;�:(=� �;D�w=����_*C;���<�̀��N�x>i=@�W��`R�X=�Ѧ��=`�X�z������K�<
���-���bmD�:`!�^�=(�=q���������)Ǽ��K=�½�3�
=�ި<�.p����<�R�;}�=��=�%=�;�K�<":=�?����~�� =ړ�;%���d?=�<�P����و���C=��.<|W�<أ�]��<�?���7�<�26=,]Ѽ��a���4�Î}<���������wB<�r=ǧϻ2:==���<��	=��<j�<��.;rq3��2x<�k'�#7���K�kc"=q��<k(�N=��#�am�<kr]�eL9����*=��<y�<g�=�<�<��ɼ�T�2�׼4i����:;���<��R�]=��ȼ�ʦ���Nۯ<��?���<�6����i0���A=0a޼���ej�<s����A�:�+;�GPK� �K����<�&üx=�2r���<��w��=q�"=y�d;gN��s�����<��	=b�&��Z=U��X�G��g�K��<#����l��k�M�hVi��#'=��.<�����I=�8����9��)�u���P�I=d��<�6+���/=��=�����l=4p��Y�& �<�Y���/=�|� �<�1=�e��b:R��V=�+�MT<�|�<�����F���b=�9�[��<��v=��\�?��<@ސ=�@=��»-)^=V��<��<50�<�`L=�X9=��q=T� =i�!�+�\��_O=@^H<�8�<���Ի�9)==�g3��]P<�o/�0�v�(�ļHj=��<v%0=�*E=�Mg<�!��]�=8&_��~�� ��� 9QX��jm�<�"x=wσ��?C=�/3��OB;w�9�2�=u�;=,w�;�dN=N����ͼ-	񼣁�;~�	��zo;�/����6<��=-C�<my�<Խ���P
=A:����=�I,=�v1=� /�{+�;�OV<]S�SY�=c9�<[d_�J�S��^�=�^�<��=V��<��&=����W;fp�~���um
=�:L=P��/�$�)�4=W���d���<;��<F��<(@H���F��o<D�Ĕ�u���<�>:<Q�<��m�Њ,=�)<=٠��5=m\=0(t�S!ռvH��[ր<Or�<p��<.e�<c���/�P=���<��]=xW��8un���=����p>��_���=�0S��ǂ���=m�@�0#=��=:\�ֺ�{�>�O�� =Y�A=�8;=M�=W��<���<�;2+N=LE =#x=��o�/F<]}ݼ�6;���<��j��4G��r=��<
�Լ�&I=Ȫ7�m���A�M{�<?=u[	=��;��:�<�R�q
�>���% =�ƻ9��$�I��<T�:=��ʼIC�< �$��{]���
=K9�K�v<\^���w:��܋=�g0���<_�;%R!=�6�<�̀�a%��U{%��7�<�3=v>8�����/(�<��<J�:� �<�=^_=!T�m��c��<�3E;�9<=�u����j�=�><������μ3P�<�p�<mI�<��<�\����(���C��;=����V�A�F�(��Ü�p�x;l�d<X@�<6✼J3=X�R�R)�g��:-P; P=Q�8��y='�f����<�ߥ��[A��Y�f���Q�5<�@��˼�3����S�3U2�`��<,UF=�pܼ�5N���'���L=H'�oQ�<�s<gCȻnq3=V�"P=��]���h='�<���<�B�U_�����:��u=ꎷ<��;j�>=7\='�-�U��פ<t��;����?@=��,�lWM�~B���A=���<�@���3��M<����kC<�ל:�0�K�<�ջ!4=^ =�&L=�ї���ͼ�v�;��#��\\�;w�=�m;��c;�	<�V=�`ȼJ��<�ˌ�E�9=0@=��<����{��[�<���V�}��i=P�(�(��<�q��4��zQ���*�<J����랼��<�Q��V<>�.����<��z�j�^<��=<@�m8�;��+=�Q`���3��6ؼD|λ2��<'��=�Y�<E]�q�,==P <6S������x=��/��A�<E�V<B0T��8�n.����<O��:��o=D]*=�i����<�����e<�+
��䑽��B=�I= �l�y�:l1*����<|U=�����=;��[=T�g=kGռ��
=G��p=�9E=��<�O<�)G��o=�A%=��p<��8=��'��:E<�)��oi�<q��<�Ӽe� �$�;�������� =�� ��w<gC_=�!�<e/Y��b�<�c�<�ה<��<��u=�wd=�U��&�ۅ<�=O�Ƽe黑�J=�\�vN�����Hi<�"K=*��.)_�z=;=eR�:.p�D!�^Q�<Ds�<��,=d��;Xf�<L�����G;n��ϩ6=/m(�|�O=w����<4�=Հ�i=���=���<[�⻶V<������X=�;v�<�sڼt�<�P���B?�%x��#H9���<.�9��ڤ�ڀ	�jL=����[]<v/;���<Z����<���5�=}�k�Ձ�<�9=�`?=�"���Z�G^���=��|w���)���S�(�%�`�<�T�îQ�!P;X�ur�V4��J�*p=�������H 2�&(�<�U=��!���0�H̒=�?��W��h%��s�<��`=����,)�gG(=.�O<{�;�S�;��;���?=�0K�'X��{�wC%�/[J=�D\�4q1=</�<*�=�$r=yKZ=��<�,����O��<���<pg'���;�L�"��<�ִ�z$�;�M<4�!;�0���A�<C�;N�; C��l�3�qp��02<��=� ߼�v�Q#"����<�;�2&�.%����1=b^�-�o<�ļ�(>��V9=�y�<�Ĝ<x���d��:Kj��;�y�:�O=�
=h�%���yn�<.l&=��d�$́��+�;�H\��*�_ ���`�c�^=�8;=H��u��<� �3�a�g��<��¼3��ԁ=X6�<d}����<��<d 0=,��;�|A;�v���H=���L�+=RM�=�w=�#5="��`D�<�4O�v�ź�Z�Tl�<��<�3����c�(�;5]=r�2d�<���<��;��f*�k���3X��YҼi����H6<��J<�)��o޼�Ơ�e�<(�=԰@<�}k;,���Fs3< �=0����u��3���ټ���S�V���^=c�(=�%9=�ߡ��a�<��-���m<@];=�l���t��ޫ;�=��|��z=%%3���=�,�;����O_=����l尻@���m�n�C��7J=( 4<�0�����b�IF�2Jv�b���6=rG����;��^�ëk=k�<�R=�>W�Tt=��T�ŷ���;��j�PV�<`���Z��<�Z=�&��&R�<�<��<�X;��3��k���=�C,=Zј<�R�O��掻&����<�e��,3����<C��7Ǽ��:=�yۼ������<��=�o�����<�U�<3$�;)����j=���Ħ<�t&=}��T�!���<�@������=vyC=�
�<T��dtؼ\|�̏;3�(=�=�<v�=!] �_?��k3=;y�<P��<�%=Q�u��.���*���u���J:���=�9;��<#p��
*�¡_<N�=!/׼[p5�e�#=��������L==�L����J��<����<�,�h�*J�sc�s�5�BK=�UY�d~W=���<�ģ�"�<o�=��Y��"��<���G�3�U��'2��K�=桽<c����׼�,�<�D.���<�A/=/W=��'<��v��i�����<R�����5=��y=Ɲl������<�W<��������<PO�]�<)��<����<�R=��O<�_���.@�|f�<���<��f�a]��{��<�����w�|q�23��V�<�v=����������ȼ�+=#F�+,=@B�����O��ς�Ѯ<��>=�Z����<*�=.�N� �$;�MC=��U="�; ���<~H��"�<`�d��;�_�IY�<u=c���v�;�ud=��b�%!����`� rI�7�*�f)< 	��a�<����>J<�)�ỔT=Woc<c�6=}y+�h��<��<oC=�n<x[�G��;�N��Ĥ��[�<��2;y�=Ȣм�v�<��9=sV��D��j�: -=}	�ˤ�<KLo���=%���92=�YC���:��Nʼ��Q�V{\��1�;��<���I�缓bu=����'�;�7=�����	=3�A��=�kI<Pt����^��g6��9@=��1<��)�]�-��v=K�O�E�N,�<+01=�)=�毼�4>��� =�!�h��<'l�[i�<BE¼�<����P=#숽2RJ��_@��B��KW�A�3��<֋�7�������� =�i��꽼��U=&��:	�̻�,�<`���I>��w�4<�d�<�eüT��<<�E=�j�=8U�<�|<1�E<u
"=դ��2t9̿u=��<�v=�������<�Q���.�����%&=�R�L[~<`�<�B�
�Y���<E��<��;a������v�<�@��M�S��<pB<��\*�6�<l�<$��<�f�)Rq��μ�y�<�=��h)�<�<��	�;�2f=�=<����<���:;����\;h�=��=@����<g<���w�D�'��K��X�<������n�M�P��Ja=���<�����b=�3<��=�-��⑻V,�����@=�g�Dg�=�*�a#D����� �P$Լ�%���P=��c��.�<�a/�{h?=��<�j<4��<�4��ˆ�9�B=J�0=`9`=�3��?Ҡ�P��;��J=� ��$k=��^�|J=ּcR��)�i��{D�a<����QJ���&=@��<�%:��3�W��?�;h�3�N/�<��d�<=��ʼ���<:c��<�9x�;�6�;�@<=�؏��U�<�=�_�b�a��=*f�l=�~�<�I�2I
=2�4=����E�<Z��<��C��0�ُ=�S=E��q��O�<{~�����͠<�^m�� �s�:4�R�l�==B]����[<|��B�<M����ܼ�̓�Z_!<,p=�<O�(=���X9�!	���}���JR��b#=�t�b��<�4m9���<ԭ�<�o
���<#%f��ϒ<�w�<���<	��	.<.���y<@�#=DXf����C�<�(=Sg���\���!�;d.=`<*J	�&�=�=����$M�i1=6ދ����j�נ4=�#(�G�;����:���U!f=�K�mF���ޯ��x<�Y�;�g���i&=��Ǽ��:%`<39=��pR���+=~��<�P���	����*=8zL=����<�ϵ<O�=X��<�_6��E�\�)�+�q��.l�p��<$��<���ܼz��;�1��4�<������Qq=X���6.�� ��'b���H�z�&<[�ʼ�9!=W��<#i0<z༻
m�[%��;���μL//����v��<h�N=
�#=|A����<d�4��K4�}����>��9Q��9<0�T:���<t�ϼ�jU<2B=	�*=�q�<?G>=���<HQ�r��U�ܼ����� �<Q��[����j9���=_��<�b�<�?�<���z1��x<��G���A�e=���<o�<=
�u9<������%���D�t=���<��	;��ؼ�� ���ּ5gW�íx;.�=�o� �G����<>��;hλKi=���_ȼ/+�;j;<��<��;3NüwvP;؉���9"��μ�ޅ<�C	<�u�<\Vż�*�c��<L��:��=ݓ�R-	��v=RW���[=�xD�5�=�8˻jh�0-K=֠=�d2�؇�<ޫC=��<��<�>h���/I6���-=��?=hq�Y�#=p�ڼw�F<�e=\�㼗�<4إ;J3$=�T��v��<kN�j�F=�Ṯ1u��#=�hY=s =��n���ܼ��@<I_��}�<S5<b�{<nh�3�K�d��<�}:<���<1A�<��ּ�\��=���<��y<��9DY�,�����Ν=]<C�<n�q=�u:=n���<+�<Df���<�:��Z==[�(��s;��5�<�叼Bc�E�0=���<]�=��g<�QJ=�K�<M����9���z$=�����:&=E]*=��y<� <$�ټ�AT=';�n�T!���b�<bA=!�<�QD<��S�T=o�=�y=4)9=��
=.S=��[=����4���G�<��*=&�5�ʐv�a�s��ڪ�0�_����v�_=/tm=;żz�R�ب�!�μc;0�:�E=�Mk��C���M���g#�(ƴ�'��9�+=h����:���9=#c=�V_=.�R��;⶚�uhp�ܹ=?3=����/��Y�
	�$!I=��輡�@�5ț�%L�<v�=���;���� `=�+պf0�<��J=g�$���==%��:MY==�u�:���<��<�xs=�%�<f�9=ÿ��?�M=��3<y·<�L,=��𼻌�Yz^<�DE��"�<RVP=�~m=3{	�!5:<o3];�M�u���aB�;K�;ш��]�(<��n<��]�7Zs����;q&����<�Z2��*�=��i=�T���!=��K=�;�H=#�n�1�;;=��A<�Q��.�<Ԯv<�軶�ڻM�=���2��~��p+ǻ	�<}SM=q�s<5�̺�������<N��<�q9<	j	=h1w=,�=�=F��<���<ns�������Y=�	#<�9�<`�<_��1Լ̟�<�"���=�a����5�h=�Z1�B�j�Y <�h5=�k=��9=v+/���;��;<�����O=l���u޼��;\0�<r�=C��<Nff<�8=�pռX��;s0��r�WJ<��޻���2>c=X�?<+��<D#n=��f�(�=�d=�Y,�w��;|\=�<�`9=�Pi��Ao<�n�)�=-�<+V��ᚼ�	=�.�;��;J>
�2h컬yU=�V�;�m���g��<v^0��,=_F=�"2=Ոh�͜�=	�/<�ϙ������.�<QM뼙g<=�<����e U�ʕ=O>e��ͅ��Ua�Q��;�<J�<�a=��=�0�����$����IX��q���)��<i.�<6����Q���c���#<�;弓��;�U���R��<�ͫ�S	[=���<�g���o��L�26;��c��uϼ����<=�<-:*�X�$�G=��=��;����ge��?<==�?=��ͺ<YVl=��L|������3���#��#�<��<=�p��<�c�kM�<�Da=��c���8���/���5�pW'=���<�Q�����;�]=�M�u���IY�:1�6=��>=;�?=�˃<c]�:�$O=��d�)�,=ɫ�<��9���L=)MK��r�<R� �6m�e*A;�{2<5T#��r�<W(�g�A=���<�Ɓ<5��;�5=ߋ�<)8=�$�<;��BH��Y����(���=��<��ż��M=Qj��0d?�����02=X`M=ȲL�1�׼2V=H�<�c���=:W��	�;��+=�cм,C+=AQ�� <�i��dN=�L-=��<�G���k<HG��� ��B3�qH=��|�����{��];\by��x=��<�Up�k�;�(��@[E=��<��<�{�$;;�8=�r<v�V����:+^�:TM-=�Lo�kԜ��u��<wp�<�V$=��M�)<s|G�]��;̓=]F�.$J������<|��<QsV=�S���B����<̔<-D�<R=��U=�t����<��6��i;�����-=���;:�<%�n;
�{�Y�H����<=,R<1����<��(=������ =?/V��+ϻ�:4=�3=N'=�u��b�=l�2<Kʣ���%<����v�Q�#�;at�<V!�l�Q��p��i�=2�b��Ep��[:=��;'�]=҄@=etӺ����0<��<?)a�|�0<Z�Ӽ|R��m(=�8�����C���U={����<e��$��<�\=i�Q;�M�9��<��ۼ��q�
�N������(���>=�����޼��G=��S-����y�T<"��<QrP�l����<h[�|�<8t2=e�<A�v<_��<��v��M���N<�Z޼M-=j9�J5=�
=vM��CA=�=9<HX����:��۹w�_�Z-Q=F}�<�i���9�� �<�D��uC��=y�xL�< ��<�o`�kN�<#�=��=���<����ހ¼؍=Ѷ;;�.��X�(�=�-v�����<`�a= k0=Ճ`=3�K<�/�a8�"7�<t�S�<�=��XZ=��;U2=��=4?:�E�<w�ɼj��|�<�/=5߼ۤE��J�<Y��~;=�0��=��;Y�Ǽ[u�;����AM�<66�<�	<�l=�Ў��t�<x�b��=��=,=&��:Ҫ�:D���}�Q�<�݇���ܻI$�<K�;�Dm<��<�ə:�ݒ�C<��:.�ɼ��N=�i=�q�^��<�j=�Q��K�<��<�t_<7�Z�����-�U!=`E��K԰;�]Z<��V=l6�<�hϻ��)�PP��ᨸSѼN	]=�j���J;{蚼�,=u��'OM�l�ϻE@ ��Y�V='$�:�<��<e`=���Z<a�=Q^�H��+�==����q=A����X<���<K�-��&H�Z�F�[�����<4	p�Μ�<7�<�j����<��G��i#@=C��<;bt<�*Q<�m�GZ�<��u��/��Ȯ�;:;��!r=� "���B=�RO���=ʵ9=�W<>ܓ<|5黪����\� �4=�w&=U����3=��9���2=��G���
=��-��`�:~��
��;5J��[G=m����=֏)��(=��;o����<qx�I̮�Zu���N�����N�O�OuD=dɃ<��\�Cq�<X!�;n�<B�y���������S�X�<bl1�����]�B^�iC\�`�<(�f��a=�9���Q����;�إ�-P4��l=�*,�+��=�+,��c�=�mR<�ʼ��V����;-�;��<�v=�Mƻ��7������v<D7d=*
�H?J=5�˻�@=<.��<��=G�-�?ql����;-{���O��\����<cxA=cy�:�n%��z����;��r<�,ځ�G��<����Zv\<��;���;��!�-/���<��;N��<yB =%'�;q���ʒ���s�Z���@TX<�=�b�<?m���x�Ku����N�A�=��Q=�͖;�+:�K� |����=�(/<�p<t�<D)A��N�;��	�m�,�-�W���W=C��<�*0�[-|=`�������DD�,�<J��;\�\=��=.I�|W=<r�G���0�(4A=�,��w�;�׼��<n�*<�V =���9. <��>;
�6=��=R*< �=��P=j��%o�1z<�
=׊&��5�XL�� QA=�ؼ�桼`�u<��I�Xm>9�ʼ�l =�k=��A=��>=�Ԓ<�?=��=;x��~���=�tf�I�1=$�w=I�M�8;*�p<m.��z�,�:=��,
�<?W<Ҋp�
���b=6��<{*ݼ���Q)V�(�=^��e�v��L�<��`G�<xtL���I=s�}<�����[�K�J�<���<��(�x�<؛=�	o�~�<�\�3�=S9�N��$�o=|�C��(=l=�n�;T=ݚ;�jLE=�o<v)m<I�{=M�	���<�A/�~��<��=�oU��Mּ��<��=�>��G�`d�[�D=ػۻ5[n;f<�Ɏ;ܙ=F$
=�A:��-ļ�t͸��\:ߕk<Ԓ.=�^L���_=�Y�<�;<j"˻P)n=�{�;]�R<����Ww��Hb=�M��'J�?��<���D��򇲼;p=�$0=Bu<J��a=c��<:���BF<e�<C�D��	=�⼞�<+9>=���^�I�B /<�#W���9���<�!=R������{A�;�a����<p9=���<��K�����=��=9Q=pX_=j������Ik<]%y��R5��?=S�>=���<����C=?�;i�4<%Zy����*Q�G;ü��<�F�;� �o7��Y�����</P�C�"�{o#���O=94B=�C=��T���=JQ����B���-��D�<�i�z�[<9�;�oQ=&O}=�U�<$v�:�u,=Г�<�L�<�4
�~S����=��#5�6N�</~�8.�}��]�v�FԊ�.�G=(�1�ߤz=3��GȻ��<����<s��=m=?g0;�;!<ҕ�<�
���v��9��N�iz�;~"4<��A=H��<FK2��ü3�żn� =��=A�A����(k<�'�;��<^�]���b=��)=֖>�H��<�⪻�c<G�?�jѐ;B�ɼgP0=�Y��޼�2u�_4I=&�ݼ��<S�;<
N_=�.L;�o�pHJ��'%���j;�-9=l#���z"=(ͼ�@p=�{�r�� 
��(rq��Ɔ����.ɪ:y����f=-�>=I�D=����߼�ć<��7<~�W�lMM����<L<�"\=N�k=V6��o�<�+�Ai�0V�<M�mQ:=���;|���L3=X�!=7/?=u�<�2J�?�g���A�����=	�V=ů&�,�E����� 	=I�<��=D�[<�� <J�k=ڸE��k����=��ռ���ܹ��
S=6�3�2�_���9�5�<1=.�G��ͼ��g<�����<���<��;2�(��:�Z��2�y���k=�H�u�-��e;=�?= s�;�T<�q\����<+�#�{��}�o�8���G�$�M������J��@� 򯼒W<��:�~��� ��=��=�X=u�I=�(N=�>C=x�|�8�:�K����;�b��M�b�V<�<����<#�.xN���-��os����;?t�!��A� �cW
=Ҍ>�@Z���O
=�~���;�,�)�<��0=��Ӽ3 �:��^<-f�<��<V�0�X�S=���;������d�]�]=��T=J"<5�Ѽ�.=lG<Uև�v}�<�M��ټ��]�+6=�����<Q6\�Y2-=�]�<&�Ƽ~�;A�H�9�g=o�><�`H��ȩ<�������<��:��`;m�=��s==�v�м�>=���=�`��R=_}���ټ�~p��ʹ����<�f��_d1=�vT�ej��1��t-=23O=��?�����7ɼ�r#=T�<�@�==�K=�g���)=�D��(b����/=���Z|r;"�-�h (=���gI���<�`=�_��wh��d�Fx�_`�<3�(��U�<,�&�!�=BkM=q��Im��B[�<��ݼ~A�^ 7=T��BS=ˌ3��H�:����P:���<Ӯ���s�R��Hs�x�=�+�<�M6�渡���H=k�U<v�M�0u=ʍL��G=������qrP�r��3'=��C���;1X:�rR<	 =����X��.=o���뒼	�<ߤ��`c�7�5����V1�<��j��2�lV�(��<�q=O�=:��<�'%<�}�C�B=���;4�<��OM���e�	a=��F="a���`��)�X��Q=Y�B<�*�<R}�;C;B����:l�㼝O̼��6��i�䚃� �?=ܾG���;@"y;�}G����<��ü�*=O���Ԉ<p��e�t<t�<ؓ��m��߱��}�ӀC�)�
=s��<�b1=��g�7=�G=0�=��ȁY<�e��OC�4�Ɠ���ǌ���<�����P=V`D<~/Q<�4�=�����R;�!�<ˋ�9��=Dh���Y�v�?�����ϭF��H�^x�<X�	��ݼ%��#g=M�f=ƌ'�i�<t.���Ȉ�+d=�w=�WE���<�Ou=,~ռ��'<7�<�+�=)H=I�6=�w=#�k;�D��l"�ՙ���=�<n�=�Tr��;=[VE=��m��p{����<�3?=�����)=�e};{�m�y���I=Q�p�K&5��>Z<Dv����@���<!�t��@[�3?:=D-�<;�)��è��d�;�� ��n =H�=����.&�ry��g%=Z�<�X.<>�9%K":+F7��z��/Q=�h���������3���Ѽ��S<�mF=�7�1�=L.=��Z��25�z�/=-z�E�2�6�����<�m��f�ȼ������<V"z�_�=�J���͙�PLۼJm�ё=��b<�<M�'�d�}<�e�;м�<��=wV�<'���J�k�T<��;;8��<�<6o=?L��Ƽ�H�f��<�GP�#�;�k���ض�b	=�Z�<�)���+���6G�ɹ=�	�O�8<�7�1�S�U�<"�G=��.�f�(��8��#�� a=��f�})��֒���<��=Y:˻ɳ�<����>`���<�{=��;�%=6)��x1=c2�o�Y=��=��HF=�
=̛��#�nO>��y��3"�<��<(f�;�o�;.��(�<�=9�/��[L�+;��<�]=�CO=�R�a�6��~=@	=�\��6�;�o�<��U=KC�;Ok<T�^�߷J���-<��0�[��<-s*=(i=�,=c���Ob=�+<�A<sJ6=��=V��<��R=��0=!��4I�j5�;��<ү0���;�v�;<P=]j�<������À�sa�<��Z<���<ʧ����B=I4�;mʕ��Q<0B���<�$��4s+=�7�<YB]�m5D;��<��U�3�B=�j	���+���y���s_��ʦ��H�<�x= Ad=��J/=(�O=�=0��iۼ��A=�!=��c<(v��i<?��</A%��-Ǽ�C�;�rI=yn�
����=a�"=d�M<_�/�-l�<�]�J�J�<w�@��q<�|>=�%'=3��<Α,=�P���';��c�[%�<3x#=4\������!��p��7���zL���s��4\��n(��k�<��<"F=�y�<�fƻ���<ա�:��A=�`��<-	H<<�߼7?�5>a<a%=Mob�C%=�h=�/c��=�+����<-a���?����</F=wT�<@�<N[<�z<��$=��k�ǲ>�ã_=���;�u���!="@�?�<6��;�Ut<�!� �h=�����p��*5=۴	���_;�p�����<�~=X�Q���[<-�3���/�_dL��葻�F@�hmH<��M��K<p?=�YU����Y��<�Q�e�=�Xy�:*����f�P���H���4=nF�<1�[���:=�.=��;�C���<U�$<ʵ=� 4=3�p����OJ^<j�5��ģ�H���BL<-�<�hc=uiO=bv�H���侼v8�<�q��-<�,���: Լ��������n��2�{�۵	=�{�R ��_��0v@���<L<��^�>������K���)��&�;���<�(�=��,�1���S}|=a��<KW=�ѷ����<5Q���c����(�=�ԻS�4=?�E<�>Q<����9���aT<��\�c&<�	��K]m=]�>���y=���Ů]�� �ku����<B�I=`û�֔<*|����q������o<}�;��<#�=���<��"=�H�+�c;�z��q��;�5��5�<�^�ڏi���5��Ј��7=�߻9�UA=a?&��=K=���<�b=�]���=��7=)�׈=Ո?�%��;�U.���)�<Ph�S�'=�U���ҼO�<�j�iĚ���'��Y=5��;���<	�4�A�V�+rX�SN��h�Z<��"�B �<��<�J)=�9y��P¼G
�Pc��|�<?=u`��#3i=5�$=l�i�x��=�(C�A��U=�e%��ji���n<��˻��߼��A;�uy�|`��-��T}����=(��=l�D�ce��f��#�K<�zN=� =�(=���x+>=[��<����M�=&3=��<``��-�<�Nn=���X����ߥ���ߺtt^=�V�<+�=��=�w0���`�q�x�;(���<=;=��ʼ��<t��5�<�1���ݼӗ=.�3<T>�<��P�6�<�����Nk<r�,�[��;9�2�X�ջ
�	=+����vI<}A�<����â�T=~+���B��<}�m�վ=�����;��H=�!�"�B=G�H��'�����ƀ��5�S�Y�`�:>a�O�ڻ�
�_�M=�`_=�(O=�d4=f�$��y;�1�:4pi=���F3�E#ɼFj�<��N���;_M�<H���R�����<�$�;2%=���\l���8����<�6P= <�\��q�<=U���[��䊽'U=R�ؼ<:=&=��<z�����<M�<+� <���<�=�N�`�4��=Ѽ��s<��_=��0=؂�`�>=&�<mI =3]o<-cV���C=+�C=��:��6�:Tq	��nܼ[�"=��˻���������e��l,���-I��W�=?C<$��<��(�MM$�bJ��}jr=,j=��ļ'F�<ǭ�<k�;��j�$ =Olb�k�ݼ�<e?F=9i.��!P���=�X<=bR=$�<j~����C<-�����<`��<O�,�T����Q����d��+�1�^�1�m�<��"=��W��<&��=��d�y*b;3��W=qʝ�.S�;}�����|����<��j���=貒<�<0�:4�S_�<�\3��E��@<$�y<mIV��1=����a`=�;�cƏ<�j'�D�m�%)��~�ۼf]�;fl���^R�Z�<Ԫ=�1
��S'<X�� �?��<v���sA���z��%=�ҽ�N���Z�޸G�=� �XW=��&=-�μ<k=�'<�L��Z/=vz��<%=E>�<]$�<�0�ylV��[Q��t�<��ż��?=<�#�Pq��r�G'=�%ټ�����.<5TQ��¼*	%<"}W<��=&H�<sK\:�iu�`�l�.�ռ���;F�𼞧������Ժ!<p�#����ѫb:>����E:<�3�&��;��=�*�;�jJ����Ž<^�8����<1j�:\��<��<� x<m�*��_3=�C/:��<��J��b#=�94�dv�a��<��=�Z�<�M%=2��;��<��=���;$h��œ�������|�>>n�,�K=�Q��J=Nd@���<+���#=C!n�F�; �<��м���	:=༼��=c��;�T�<1�[�t3V��� =_G���!=��&���Z=���;��;���:E=�<fπ�5��<	]�<6^;�g=��X;]F^���	<NP�<Q==��d�s��<�
<�P��_�<�l�5Fe���=�Qk��ym�F����!���8=1ŭ<ب��.p=�����Q�Vw���:&�\F�x����/�	6��6b�,(�K����]�T�$��ă���[��;&���<m37<*���ub�:�P��m)�Q+�̕*=��<U1'�DH��h'g<Ȟ<�=sb;=Jh�;>�<q����iX<ِ�;<ZJ��!�E�=�� =�o���X������^�);�<�T*<zt7��Z��x,l=:$�<6�k�p]C�Rܼ	�Y<l�-=`=?ʬ�o\��B��H��C��j=��e���Y=��i<�EV���<>Ũ<�˔<V�i<�xF=�	9=f��;c�&=�Լ�G�_❼#�u=.����* =[FW�B�j\<U5μ��[<C4Y��l�<I&=��<o��<t�2�{�<�C��v=:�	��Ne�ѡ,����FC�<�-E���v<Xz��Ļ��<��Q=yj0;�`�=*�)=��W���<�|D��u[�A�W=̔J=9�<#w<�CL=���<����<�<�8���J=�����#����M<��o��<]��;&����H����<�o�<�"�����w0��8O<�Ke�X=�<K�	=N����M��u�;���T���H=�O�B��8�]r<�<��=&�g<u�L�b/�?L<KbD�R��˘޼&Q���\=��=�9.<��j�3�ü����6���=e��<�C�93<��)=�z��-s<��<b���2�y��N=��Ƽ�kj=훇<ǧ�:�Jz<t�E=L�"��-G=��=�4j��b�<�E�<#�=���,�]q9=;�.�2��<F�<*�#=�8��w�R<�=/ W���<)�:��=�LT<ٰ��"B<�Z�<*'=-��/ܼ4�=B�b�J��e��5���<H/=��{��b8��rļ�����)=_��;���:?n<_\��N�����D���C=,��*�;�ꉼ$lڼ�c<>R=���+_�<$�<f�y����<B�=!}����-���g=Nua<1犽?��E����< �W=��Ѽ7�%����<�m��[�<��=��<��l=.c2=�#!���;��<Pf�_�BV�<d4*=������#=�,=ʯ<=��
��}�;Z�>��]3=�ā���輸|8����H=r�=��<����;(�X�߶h=+b�;�<�N�<b�<_���� �����<l=y�z��@Ż��X=#r+��ek<��;]v����<�x�V���¼4%V=��9��z-=9i�<F�8��e���r���(<N��<QT�:�im�c��;��O��3�<�8�c�0;�O=���<���b�!��\�<b�N���{����<�z!��c=lw���b=��]�vPZ=,V'=�.�3�7=>�"���m���`�[<Ѻ�<B���+d��Ok��c(�R�<
	#=�aA��U�;p�v���<=aN�<�}l���h=w(��H����'<�j�<���#Ed=9����AD�H��܃<�Y�<�Z=	"��^L�J��:�����_l�H�
=�����@�����;Q�;=��r<�0Ǽ`c8�՜�<�
�(�>��<q�=�R��Z>T=%!=�[q<m!V��f!�̦�����< ����1��G��݌�<�x�<�IO�L��;:2I<.E��f|�<
oP���<�W:�eF<��Z=��<N�B���;�Y:gI���������?���<=��M=`F
��V=�P(=��=��=�RP��L㚼.:<�5 ������@o"=L
��/&�6D:=?/�@����W<��+���N���+=P|=4��<3��<���$^X�fun=#��fh3�˅"=�T=��N=���� �#=Z@=��u=4}	�l�<�;��+�A�Ǽ��ݼ�3)�P���Q�C�:�W��5���=0컼�*�b���H���μ���h���~쁼f#r;�;\�WX�<��X�^=z�<�0��S̬�@�<�x�<-�;�/�<���"J]��pѼ�i�;������>�;�</m=M��<խ��u	<��v�n���UP�ˏ	<k$=�Q�<����O>���<� ����?��7�<p	�3�3��s�<H!Q�mм� �;(|=3�!={��<8���׼q�n;�{0=S�n=I'=͵;=x\��唌�)s;[��;]��:yk=Y�D=��<-R��k���B�w"�>�O��:�<��<=G]�<RD<��=��<�A6=����D6=�;���<H�=�Ö�)1��(���Y=�g�}];�<���;0����~<JR���޺l��g�6=*�3�Z�m�W���G�k����5=��{�**��w�<.��E����꼅�H�hʼ��I��<�Jp=��4= �W<�o��&o�.56=�'�<���</�Z���*��������<���<�D8����� �&=��<wD-�Flh;G�=Ϙ,�M^�=y�=�����^=�Z�e/ʻԐ==`�<��=��<^���A&=�h&���-����S�?�<�J�;���~�g���B��k=L6<Q����n����?��'Q���=%���y<ǒd<\_?�N%=�] ��'�<��<P><Go=���<@=��<&�]=�<a�����<'�G��^�Y8k=X�ͼ}'�<�!�<������ �t�<�@Y=��	=����m;=E4޼kJ<,v<:�<���<�Q$=.�W=ji�<�L�$�<{^/��o�&�<ƻ��vj�T�u���Ѽ���<���<�2r�� ��	��+�M=f�*��=�I�A�Z=��b=t爽ʲl����-�<�x=,%L��/<˨A��Y<�c<t�==�>�ٕ=�̚�<�#<�6üj��U�f���"�P�^��/���
�<`�較 $�A�ϼl���G��{>�:bc�oa�<l@���:=E�<=	&D<ܩ!��xP=�G��- �mz=����0��:L���i=DX�<_8�E�`=$�=����?��V=�=}<�S=�'{=����S㼂��?.�E�B=�_μ\eK�<�U���	=�M��2T�=6��]c�� ��T�d6<�=�����|0��=�7�;$Oƻ{N=�ހ��"��0<:��;`z?�%GF�S�N��8�<�乪� =��!�\�����	<�8��y�=��<*���.����L���h���|]�;��1���2��[�<�� <�4<ڲ�<���ޗ<��»�H ��
=f������<K;�2���9e��=�a�H<�Dp=�<��a{=r�/=���6k<��=LBM=��
���i<��'�B#����:~ѷ�R�
=��C�G=9���#5���2�=P� �O)X�+��4�=�q���ڱ;�)!���^���w:B�e�X >�7�9����<����?'=���;�=ȁּ���<=����T����Q�t�[�8���A=�#q��rD�&@)=�{G�VѼ��<�9�9S�@�����Z=���<\#5����;�r�<0��<��t��I��<@��>B?�>a=F�Sǿ����;C���k>[=�~�Q<�"��tz��L�fU�Y=!�e��⻣�^�|�ؼw�;�����h=�c�;Z;=��*=2>ܼ@8�N���@���u=MF1=��m;PRż�i=N��<��� ]�:i����"�gfC����<��F<��0=(�U����<��>=H�;�
=aC�z���BQ=3CP�͝#: =���:p~ļ著�g��s�,=q�U;ż2���=�5¼GQ��X�X={0=�^]=/�;��b������� =_4b��<��+��)X����<��(�%���/=B-�;���%]��y@�K�B�P2=C�S�]\	���K=n�<�#�<�/=S�߻̐�='Ղ�G)���j=[�i�Fa��Ƽ(b�bx�<�[�9��;��ĻA��<��S��2��h�ٓ����<�]�;���;_'��=<R=7
��PND=��<�8�T^��qA= �4=P��<���<v�=���ֹ�`=nEɼ<,���l�޻(�=�ي<6�f<�5K��.%;lb�!�-�f��<@M;�$<�ć<���<J���2=�x���2=K�4=��Y�Y�C=��=�W=��=����R�<���F��<��<HO4=gu;x�2��߀=�,�<æ��"f� K�EI&�Tu<??��
��<4�<:6X�<�2�5�`�X���+u)=�b�;�8J=�?�� <=��<kU<:�j���ļ5_j����;��<���7��u��:��N=	)=ν�<��=\<K��<~��׈=6ʇ���
;���<����U��:Mv��U�f<ۀŻ�up���X�4�N��}E=��q=W����=�?Z���<�X5<;mӼ�� =b����)�f�}<�¼h�;q�=-b|��L&�̱�<B= 9(=�=z<�M��=(Ƽ���<��
=��j��*m��U�,|�w�Լ�A��`r<	?6=ny���9=�0�n'P�}뒼�&W<_�/�M7�@;���2�~΄��B�<ꚱ��pW�]V�<�k=Ϡ�;&U-�67=�$����<-={�$=�=0�<}�<�-�;�f�=�=��<u�s<`�Q=#VR=,�=����5��5����P�N�><I"=���͖f=�)>�wU<�bw����;hjȼ��틻's�ǰ3=P��X���P<�����E=�P������,5=O�=i:i���E��,8���L=�d���3<�bA=i��<�u�<.�}�$�L<�¯;��n��S;��v<A� =[(N=�`<_�;��<�6��<��=Hg���%=��nN(=l�=�(6=� ��yY=K�ݹ�'F��{^=;r��0T�N�*=�3�<��=6v2�y��<u��</C���<���<�ZB=��dC��0�	=�#����&��=�OM=��{��Y�A��M=�=����nVv�cw	=�ڟ<�C��+�(=Ϗ�Kt����3�<�)�<��<�/=UwG=�R=B^�1^U��=��4='�@�?����<��<Hkm=�e=��<�*=Hſ���F������]���T=(| ;�#^=3Ӌ���d<e�u�4��V����<?0	��(!<o梽 �<�v���F=ڰ~� �=��O=!��<�=׻��;�,;ة»Oe�[�[�0G7�)�<��@=n4<��=�����X8=�(=�5<�K=lz;��C�<e�/��h�<��_�s'�;�%9���s<�}�;���<����;��N���=D����<z"=����M��䇼����6R<�3B;�N�;$�׼�&=���<>�=B��< 6ȼ3���G=� 9T�e=ܦ������� =X�ܼf=L�<g7��L6r=yڼ�F�<p�;Ȑd<�H���r�me=� ?=P�@;S� =O%"=���Լ����������%�=	@���<N�%=���;,���q��h�<��z�K�c���� C*=��g��8�<�ǃ��}>�%=!N��x�n=4��M*�<�i�<W�J;���'/<�y=��m;iA���4=��<Y�M�P����A�an�<�ɴ<�hռ�	���=qf;�	:��<���<7�G=�mC�oW<{�4<BL=;)=|q/��o=���ȁ���4��5=��x=��y�B�S<���ePw�<�y\�GM<m�=땶<�C�;���<�4\��` ==��He[�V%�@I�_$<���<M�=�����W�M����{A�N$��X�~�,Cr=A d�p���/����<���<�ټ�=�t"�A,�<�%?�[�$=�����o�8:�kA!<����o����<�JN=��A���m:�������<C-�HA�:���a�r�u�:��F��@���H;�B�;ݧ&=�!�;��/���<=Sk�`8����'���D�<�㼁2==�.�= �a<�a���0����;�m�=��<v���{8=�����:=�\=��B;e�Q��܌=�6=5C��6;0؆<�3=	���[l<�d�y#�<�1̼h��<����~8��[��R��y`S=��H�y�;����Be�{Ӑ;ެ$=c)n�T�P����w�I�I4=�J=U�9��Q���<=�W=E��V=����7�,b=3��<wT<��j���YG�#�*�;�;��=u��̭���=��JH�����ź�1Z�0�L=���ˎ�<H����W�$�H=�t�VL%�Ɣ/�,:�x���j����U<�nX���ٯ=`7�<�r��a�7=	o�<�m;��!�kG�=nca�:��<�27=q�==h�<m�߻c�O=f=&ؼp,Ƽջy=����I�< ;H=M�3;ׄ�>6,=5ü�ǻT*�7VY=o��$�<���<u~B=���<;<[Vq=�W=�<ޠ�<kYN<�.~��fJ=t���D�<��p=���n'�ٺ<CڼW����=a�8=~2�<(pI�Q�<N�<�
g�9i;=��#=��=��<����D�3C��%Tj�����u�=�1 ������x=�y�H:"
=�����=A݊:�F�}u< `��[�A<0�һcy�<Y�C����<Μ�N�0;�u�=��<!��=_��e�=>�8��,"�Np�4[U=�����<e4��j�4��B�<�=W����;.y�;��L��x�;�o<N�$=�U=y5}����#ͻ���z�Լ�=kd��h:\���Q=��=4lE�'0�:,d�<�C�ե�<�U@=�G�<�����n=2L��	#����=���<q��<�ݭ<g���돼A�<�Bp=D�8�����Q�;�	�N�y=� ���f��<�t���f;C�<��<E���]�=��6=7}�<�5=��=��1=J4�<�D��1=Yz=��c=�	�;����.�<��#=7-�<���< ��;�w\�φ�"46=��T�~��<�T>��j~<�Dc�?�P��
���p<�ۻN�&'|=J'�n�s<Ӹ�<��{="����~һ��0=�Ҙ��v	=
d���[������#=�
�����Q˻z����Q9��Ao�Em�oP�=�h����<h]=pvy=x�<�:��p���0��ׇ��	�=j��� 廎�[<�<x;�'=Vj��Q)=\h,���p���+=��<'2s����~�)!=�uV=4�$<ٚs���<Ab�]��&K0=�s�<��<՛����:k8:ї������ �8�B�H�I=R�n��J� =��E�Q�G���0�_ʪ<5�8�=&2�Oy�<���öD=B�<����
�L����;[=%P�<�h��_������<�sW���=�\��m<);E<��4����\x=U=˙=@��;��S=�=�=���p�J=/���O$��]%���<V��:�?��d���Q�`��<S���y�<���;��J�ò>���G�1Զ���4���~�3��<�;g:��̺��5=�qb��\<(,D��3�<S�;�(���q=�3D��p;=�&���>=*��
)��x��,�qɼ�栽�t.=���<������\;�������;{��<[�;*�<��<P����π<������=�S�����J�<
�>=z=��9���H��<Y�ۻ8N�T#I��/=;=�~�<��Zf'��`<?7лop�<��)�Fa��Q=r=��N�+��ޮ�UԘ<ra<=��A��`��_��bYG;���<]��<d�);�i�_��<���;� ༽E!�r���)I=�!伐�<��<��<��=:e�<��#=�!=(,�<�g��6o=���<�f»�=r�����e��;y`p;�]߼@�˼l|=l���5�<Ҹ�;�8�;;���cA�e��MK=�w���\=��S=ܪ�=ġ&<�#?�m=���<Q'���=9�*�x0>���Y�=�&;���<�DK=��$��>=�v��>�V���B��R<�7�ر6<B}�������g=�F�<\��W��R�����a��Ǌ�:W�;�A<b�;
ӌ9�j7=�,<���<�h=����d=�n{<2]��3M�D�^=,'ѻ3�;�Mi<�L<f1P����O
��?�<C�����6<Q�.���%G����E�����N� =eܖ=��׼Z$9��漓�d��.U��<�QP��4�<�<���<�&=�x�;/����<s�$=��^=$�x������<Xy!<��(=�� �q!:��K��a����<��q`=�UM=�W�=h����ϼZm�/��~s��=�Y<�=�o��Z ;&+��ؐ�i��<@4]<��*�N}<=w�=AT�:w_����=�}Ƽ�I�<V�J=s�=��x;7�<5��<���8?[;��n����<��h���ݼWy<�C��{��&=ga<��=��
`�N�k=la{��y���1=�t�<����a=��C=	�O=�40����">�v&�77����@���H=EX�C!�4�ʼ,�y���L��'�<����a�� =��3=� �+=)]��4���=�ݵ��U=^1@=�[8=�36��.����c��xm�����T�;=ݫ����=HS�㡼}`==��E���S��+Z:�c�ρ��!��<��9ƫ����<���K'=�.C=����30<���w�;�,B7�������<��Ǽ�/�0ӈ��vQ��o߼��<��3=Uu=]3Ӽ��=M�U=�S'���x=�=E=�r� ��t���7/<*n��w%���D={��<�.��fz�>T˼�X�ƙӼP�h�ć�j�&;�(o=�U"��'��0t��]<)���[-˼����Ou�X=�b�h��;A�O���H=W�D=;�:<�=�<�=A�A�=R�v���=��<u=�b�wњ<�>�=�r=�G�<3��}���+����^.d���f�=k��_�^&=$��h�<�!���<e��<Q����ע�hA<}�B=��<�f=� =b�������W1��1ͼ3e�Ζ�<	5�GW��XO�S(;`�3�����
��������r�c<A瀼�?K;S��J��<�	���f=��}=�h=���<u��.� �=�v	��+̼��.���%�e[=2nR=�I=�� �ehL�= /�pR�]�@=?O���<�"��f��<x�_���+��@����4=�,�b�
=[��;I��=�@���e=�.�]�<�a5�M~Q=S�컃�>=��<��r�?�h�Ym�!4=�#)��9�����<��V=�=�b�;]i-�N��<5�=]"���z<1\�<q�>;M'�<�XL<��)�	��C�=xt�<�m����#P����]冼Gӭ<�*�<G����@����;Eʬ<\��<�N<Tx=s�=�Eݼ[��gr�;�q�;8�#);���=*�=,jӼ��~����;���<��*=֝%=��=m�/��=�$�W���7=�[n<Zk��y=ږ��f=#��<S0=;�D< �L���k9=�	�����<�8���v�Js�:��q=��X=���;_Լ�����1a=b�`���=N�K=A�v���^=gB�<3d�<t̼z$�<BTӻr�<ũ��������;��=ض���"=
&�;����w�<�1\=�t�;XOn=�yG=��z=H��:��<��C=��d�Kj9M��0�R��=:���<u"�<�|d�q��D�˼�܂=��P�� �<W���"2=�
�p�0<h>=2w�ؗ��,�P���-��5-<f"��.2��*.='֜<�༇ؽ�ǣV=�NO=wNP�)h=�p�<��<�{4=E�>=XOۼsSü����GJ:,�%��9���<���<�)�<��/�SBf=-kj��C�M��<�Ya�(�r=�F��Û0���	�Q����k�<����(��~=a#=t8=
4=��L��B=��̀�������K�>�����<c�s=Չ�<�nI�9�,��<�F�u�Z�5��+�<߃N=���;K��xB=�dG=���|>��W��ؼ�I;�Ż�t�^=H���u=o�q=F*-�ѷ|�x�$���мN�V<z�U����hD�^"輣�P<���;�ą=��+=�*�~��\��<�q��C<d_�=Sya�e�<Th����/Ɲ=��=�"�S�:<�t;�̋��u@�-��=�(���Ë8��^=#�3=[ݟ�3zQ=�`���B<�bH=�5<���<w�F=����k%C���^��$u���!=.{x<�W2=�,=�	�<]Ǌ=�`���������; <HM��#�<��꼞ow���=/==YȂ�OO�;��g:f�+��6��4=&�<=o3'���/;)Ț�ݛ�4Y�<5�\<w�<��'�x�<:�ּ�c�<S���Ͼ=S3!����0>���[��ב[="B�<v�<o�)=F	=G�=&@=�>���X�����<�M̼8�=��|�M�uR=�C^=T�ɻ\B:�=�g<����.��^Lb=�~�;12?���û%x5�䎼�[��0@s�'z;���<�Y&�}DD=-z3=�N>�cӻ
��hjQ;歼;�.<���<zvD��C�<-0ѼD� ��ӻ ����=���;��97u�<��ͼ�L2=O�< <�<�=@�.�l.o<���<�H<�ق<��¼�Q�;�}�{>���=�������E=v��<-�<����<c��
ż�*o����F^=���<�c;:T���w���<v�<�l����:{�0=�(��>G��Q==��=ռ�}=XDǼ�R�"P��j%t=Z�/�v��<a��;-�><�e<Oc�<@O5���;��H;�4[=.n.=�c<��ļ�Mk���<z�o<@�5=b
O��;�<�*Ǽ:�7����9��m�atλo�P�Q�GV���4p���$<�ja;�~���+�{<��g<�X�<��E=hC�;�۫;��M<,y-��P�;��;���D=p�I<�R����y=����w��=Q�t�#���R=�f���~�X�^�ު��?�=�pջ��<�m����b<A� =��b; �z1�;z?鼙�S�[���d�Fw=9���T����=x�t��#	=��<��<��=���;b��<��.=��`�{�W=,	<�t�<������<=v��;�oL= U4���Ѽ%c�#��{���>�3)5=�Z��e�2�1��<�!�<��,�B�p<9Y�<bb�<Z)��]=4�=��wм.y����>�C|2=����r �n�L��%�<�z���a���g���<z��;L��9�q�Rh���*=Ć���-:�Ψ<�B��ѻ<��#�iEG� ��+�<�4꼿Ή�|r�=w���β��J�<��y;C��<�8���j<�Ϛ:�%=��=f�<?�:��=O`�: J:=^��<�ug<��L���<�Np�<��;��L�����f=n����a��Y�<P��*�/�:л<��J��h&��>����=�F�<L��<�}*��^,�8<=<���&�!�ռOR-=��<<��;���� ɉ�*�p=@i<c�4��Ta=�&���v�**м�n�<�;f6�P�<�q=���<شA��~?=W
��VӼ|C�����}�u=�Tm=��n;D�<f��"�<� �<�H �_�,�@�
��� B='Q�;>L$=9M=e�<�v= �<�<��<=�=��'�����kb��ku9N,=���<nn=��*���_�W�=ٝ@<o���h�:�[�<.�B=�;��S=�/��\=5�:=5S���;8��;|v����D`���T����<�S��;i�<�&�<�~�<�?����<�[J��L/=I�V�t�"�=��7<L~T�3�T=Z�O;
V�i�<0�:��Y=P�[=��a�78s���}<�'}<��<oU�<�l6��
=���N���J=��^���-=�	�<z�=&���
c#�5D#��<�ׁ�����
ϼ�r=|����mQ��IƼ�w��V�<��N@=��E=sjA=�s��ɝѺ�	\�q�t��=T�u��M�)���T:��������PA��?.=�Aa��}=�_�<�1���
�����7���M7=�-ȼ��<���]4=T���K<�=��'N�k��<j�'; Q3=A����<��
���A�5� �D�8��;=	��W6��¼�_;='�V=m���ڭ<S�4=�HQ��Rw�g0D���=��F=p?�<��;�1=O�E=}��<�-��r"<*����j�N:q���?;;|�<�jo�_{U<��=�!o�O����7W�N(c=��<�p(=���;�	=��ƻ��<��<����i���qJ���`:�����a�R���W=MiV��J��s@��v�����;�F�tK���>�]6=9>�<G�>=Q�����b�#=^ב<��=��:��s�00�[�f���:=O]H���z=�!
�t�<�J�<i�%<E\�<%��<����-��<	m=�E!�P�,��H=���������ȼ���;x�<�D��,r=,/��8� =-��;<�ё��3=A2�h*�<�= �ʺ/Fv;��&�{r��<2�<�����м��V��F=��F=.��<Ž�=�=b	���j߼��0=���;��a�'󃽿��´�=M�>�����<�C�<x��;�W����=3��A�<�Ϧ<�O�<s�/�j��<ު�;a�<P+�<�~=�?=�y�����b�L<tAD=��� �,��R=�H��K.��m��]�!�N='�����N=c���Z�<��<R �<`�,=��:��N=_м�4���H<X������B�.s_���D�|
:=nCr<�X=u!��>ļ��x<��;{Z<�N�<�����1<ڍv��}Z�j9?<
�I�h3���<��$��D�;>����<�2���u<���<�$�<�G�az=N�(�A�<���<M�T�-��<�#=w�==1=~[�e��<�\p���}���L�D�R��8(=d�@��y4=~��<�"<I�p��Y�z��B��m�<n�ռ��=�
��wq2�8oK������M�qNA= ��<�� �r�Ӽz�M=�i=ay=���<� ��t��B�޼�c���;��<,w��4;��B��F=}ܵ< �F=.̼lG���
)=	����<�h0={�J=SM��2�<s�K�7�Z��{���O�{��<)�
�Շ;=*���'x�bP�φ�-Y7��g�����<=�N���?=�}%�
`={����;���Dv=7!<ҽ�<��8=G1����{�Z�1=ň�<�X]=��b=L��MF�<������<
b	=�4Y=h9:��<��<�����-�3f=���<Sa�<��F=o����O=��<ǽD=��v�@R<� r�����Rw?=͎M�2��;�;���.1�*�@:�����b�=��<!V�<��;�͸<]�F����^q(<��<�+����9	!��k=E����=:a��ڞ�<�����;n�����=	=N�T�d��R=F����������<�\<��9�k�=m-<���gż��A=s��=J{м�Q���|���s��1�]��9}�?=�t:�]jP=��!=PJúq��Z�,;L	+=n{�Ki�<�M>�( �<K��<�`r��]=4����y�3�\;��X�U�<O�<�t�8�#=�_�<[P.��+=���;=��p���<�]=U�o=ê,:j�E���z��9=�}�<��@�|
R�*��<T�Y=��f=�^=_�<1{s=���C�<]��<��K<����e�<�'�C<��o�g��.}�rs5��=��N<��B=�4�;x�I����;�=�Ȯ�����<���P={�m�oܸ�"{Ѽ��Q�b�<j}�<�B=߯�<DG�<�'�jX�:6a-�W7��7�8��S=c�<�CѼ�l���`<�DR��;�<�n�<���<V^�<��d��.�<��6��AN=o����<[y_���8;a7!=�i��Jy�<�*=0#u�`r�<��P�L�E�9�L�YY<˶<>pT=s�=�e=4B꼍�~<�7���	<y�"��X:+��4�~�.�r����	S=a�h==��ri<��P=.�c�2�j=ط=L����5=��A��!���צ����<�(�<}�*���>=ZLr:f#����;˘��F��< g��=�����VS�e�=���|Wd���;�S}=��B��케SJ�rJ��D=t��#�����F=f#���|>=�X�<u�/=��[=K϶�����9j�ZB�<TKa���4=���e�h<�ɇ��N=���:�T0��fI;Uh=S�<�W'��{��$��<[32��V�����f�<W�=��{�5F/��K�����<��=JC����&=�X��Ӟ:I�r����˂Y�L������<
w.=5��:�:]={Mu�^$ػ�y�v�<��==P=�|�<��˻"０Z�c-=4�=H�T�?��<�!=6��<=.=DfK���<e�.=.L=��y<"T;=LW=�Ö�z�<� ���<�z.<*t�<�I=-'�Ъs;�$u=	�����a}�<��@=��<�IF=�T�<��F�U�<�w=.�ϻ����]=o�V�lr�J�s='F(=���<6#�<���<(�4=�tp����K+=xO�<�k���6=Y���D�Y����<����0�S=� ��;RL�<���ʂ�r�����%=�� �jh��s�(=�o:y(i=��=<�j�|��<Y����L�}?�;���W����::=nLx��k�
˼�1n<��p<�Z�=� =^�Ǽj<=�tQ<��Y=C=�B���;�����R�8뵼�0=Uh6�����<β;ۚ7=�J���?��8ۼ�����<гv�Ly=<j��z/+����=��4�C#�<��2�$�R=��D��~<a�<P��<��X���n�q<�<�]<��s%���C��#����,@<���]�=U9��==����p����Il=��e�_W�=}�<������$���]�	OA=&��O%y���;�QUż�K���A������_�<�l�9JZ%�hKI;^�D=�#<L4�<��=U9�< �Ӽ5���x�X��=;��7�μrm7��1��cG=�`�<:�0<ۂ�=3���\�<��$�����-r�<	̈�����vWQ=�����</+��A��<�Z=1�߼�;=�`=���􅡼�\{<{�<h4M�
�����= ��[��T����/�fh���=c�6���>��i1�E�=��z=&�	=�w����[��)�<B�=�H��A�J��������y�<�*k=nv��3>�\��<e�1��/f=�P�<�I����'��L=6�:g�A�O�T�O=,�Y��*'=�d=��<�3a���;i,���k=ω3��W����˼D�v���9�;B�R��9��<h�Y=�
=�����}�|v�<���<�z���E6=y0=F�J��/���A�`�!=�0��N�����5�%}=�+=F����� �� �z{o=��/�[Ֆ;jP7��s=]w��Y��0G=\�9��(��������g
4��NB=b3<���;��1�M=d=M����=}rL;v�>�`ь<^�=�E�jnB�q>����;�$4�o�=ƅ�<��<U8ڼD�<�O�<�Ϝ<S0/��1����O�_=rA����67�Ǐ9<�P�в6<�c&=���lg���N=��G=ܢ�_�=��=��&�=�a<@c��wV=�m��5��������"A=�1$=$�,�]p:D;���2?��/�<��#=��4=��;T��<��B����=E���`��<� =���)���!�?���<ܟ{�ǐ�=<�8����:5�Pd˻Z��<T#=xQ�Z���4��gN���!<M��;o��<����J���7=�A<�w]�1/����:,7�Eu��h%�:;9��<��==k�X2����
��$�=�C=L<�%Q<u�X=/ =��=�����G�; ���!i�<4�3�^l<���<��������><�����g<=(ͼ.� �^<=�=˼��d���*��\=bH=��<���-;�o1<�9���(=e�<����e�ӼZl<�,}=&���aQ�<d�	=|�;�7��)ټf���X:7<�e�9��9���<m�+ #��ر�*Z)�m'W=�E�=ĝ=�����2����W�����<�0}=E}�<Gk=���є�1=���9�<=�_���=ߩ�$=��'=��1�v�"=*�+;�h=��W�֯��ּVo���<�4y<�Dּ��B��=�]��2;<�q#�$h���K���ȼ�ͼE��;��༡�N=�Wy��Gl�_���IwQ���;��l=����j��"�W=��»ɂлvu���=��A=[5<~gn��S=��<vڻAp�;�u�M	�5F2=W��,W�<���9{	=�pF�8j=�_M���b<�_�<l/�<(E=���<5Y���P*;|�������,���~<��;) ���[*����<���D]�<�༼5�<ʣ��4�7��y��yz<1g��(��I�<B���g	=�H
����;���G� �)=2�<;J�ހ=���,i�<��k�L야�6�!'*���h�k<����0e�j�o��:ļ��9�b�;,�=j@���(;�L�<C�üt	r�Ԭ��f�#� <_dмbG=���H=���o�<��l�<߀�<�;J��?,j<��=�.;�a���<�M7�jV=NRw���=[ֱ<�[D�/��<�ܻ�v�;���;�k<^���tк�+�<��9�^C�<�<=n�=�S=^<�g��AL1=��<�~�<i�a��Rn=�ʆ=���������<��<�/�<�.��;|=}�=@"伾�K<bZ��~<�<dZ��;=pj�;ϩ�<��<	7���铼�O���;�r=_9�<����a�:U���q=C�ҧ=�8"=��_F׼;Ɨ<�>D���=on=��H�<@ힻT��<�:��pQ��9�.|漱:7�R�@=�Ｄ�<�"��7�;��=�q�=�C�Dc��w+:��ü*j�<>%=�C����E�5��B�P�<5�X�:9 ��c˼)�[=d
��A=�9V<Ƙ��=be�B�=n/[=T�=���zuj��W	��Kq<Y�Ƽ�|/���n<�%=��f��kb��8��=5�м*�;��q���3<
7��?3���߼��W�_�k������I=�3Y<-��<�������ť����<��a==��<��;(��o�������2=H�H��w�<�2�u��̾k<[����H���S=��<@P���<]�]��
=@��:��l����<f�<���#��.I���<=B({<��=������_�?e=��<+o3=�{]��/@=:�^=���<��r��<oK���5��p5Ṥ��<T<0� �
�t�-��;1 ����T�*<��ϼ�������[��/���c��t;�{=�̼��鼤��B��X>#=#j:������;�W�\~����S;�k�+��v��<J,�������+�_��:���?�&����<�o�<l�����a���#��-C;�T=�L@=�)�<�9B=z1 <q��;�<<��=3%H��E=q5�٨m=���暨<�s���$��d�<�'3��������n�:<��<z�G=d��;Ut��2�5g�v>�
�BfT�r�e=İm<���o�,�Mh%=e?$<�T=Ki�<oW�9�K�eR=�&=� ����b=��=�.�=g�=��%���K<[���5;L�6�,ܰ;k�7���T=r<$׷<��%�#�m;ʖ�����91�D�N3A=�+��u�޼����Q/=��g�������s:Ef뼻�μZh�;@�<x�-=����t8�L=(㫻�3[���v=���4$=xZ6��7�{����<y`=�=H=��@<�=;�Pv=�#�$�輄ś����<�su�?<$�3=H�Z����)�=�m"��C���:,���4���A���=�qw�n��t�B�;�����Ƽ!h0=$�ڼ��:�b<z��<n���=ؼ�m��C�J=B��<:g=�D<$~��g�#�G�h�>҈�a+`��=,h����e=!�{=h#�<�%U�Y&��gM�5(=��<��y� ?=㝙<�@?��c��۵^=y@��vk���=��4=���L��I/���!=�y�;c5���(��2G��dE=c��<�2�i!E�[�q�+�;~X<Gд��E�<�z=��=	JQ� a�<�P��"�G;d�=_{����o��6�<�5U<Q~ứ,�<����*�O=�G==�<�琼ni��ֳN�X �9�<�����Mۼ��*=���;`H�<��#���=�Ȁ���1��*'<�,��� ���g=��;�P:�;�<��Լ��K=�P,�ǳ��@.6���=?W<�G=�('=��ļ0��-e�=y=��4��_Z��t=Z�<9��/����<$."=mX3�}���7=�<��':o>�(=�y1��(=�<�Q=�>���0<�8�<`��<��0����<Ռ�<7�L<��!=�b=���Z-�<�,<S�8=h`�<iD=���~�H<�=�� �e٬<V�D�M!W���|���<Ԑ:���C=�X==:~<�b��n߼� �<ߕ=iL3��D�:�v�<��;��\V;Ǎ����6�[���0��<>ﱼ�H4���p=��μ�}=���:�D<�t�<]g��<<�Wv=��#��נ<b<ڣ�<iS3=��=�a�<�V���*�;�ׅ<԰�:� ��종<��t<��@�X�='��<��<�5�Ry����c�sv�<���<o��i�����$�2��<6l�����Ni�<#x<�����:=��&�B�@�c1	�{����=0Z�������<o�����=Z���y���o�]5�r{?<T�:���;ͼ�K=�Ny<9)+��p(<NL�<o�<�&��sy�;�(�����<�wy=�U��Ю<3�^<K�5="�Ѽ��B��]='Nh=��=��r�x�=�,H����;:)=C��<c<�n}^�&� �բ�P�u�V� ��>,=�ō<��2��å�����P���-�<Q{��`j=.�8H=C=gJ ��;p��_u���;CE��4["���-��w�P�<�a=�L;�#����R=��<֠�<��\�Ѫ7<�1�<����o3<���S|���W�<��=��&<M�*=��9����-.=a�<%��>�6L%=��=>���AB���<��f=e3��a`��߇��3=�~<ߓ8=�GƼi@߼Ң���t=4)<1R	��}<YE��)���[.=�a@<�ɺ��ݔ=��U;e�B=���<����X��	,���<�d��G�`���ἡ���/�<6SJؼ��;'i=N0��V==�鬼9SU=��w=d⼩6����<H�Լkϐ=4K$��T3�1�<��E=��=\8�<�N=��f�0�&o6���	�K�������9�"�<E�R=`��|6=I9=,�<-=�81=���<�>�<�6D=?=V�18Rk<�s���]��-=I=oW=/�Y��{ �@��<�}1=�3�<9��'g�<�Ƥ<����<(�"=M�<=N9���;�ͼ�<LY���je<��A=u��m�'�ԝ��m[F=N�<�e���%c<�Pq=E�J=\#�;�4p�D��<��<�a��t�����<v}?���5=oZ�9�m�2��:
�a���[=���� 4<zV�O���q�=`l�<��=N[=p{�<)N�����BR��S����;/��:0\=���r� ����<�@F=?z�9�q��~�"=��_�ٕ�;q��9�=�"��ط�<Ԛ
��r�<G��<N��I�l���Y<X�<��*;�i�v\�<y��;��F<x��=G~=�q���m�Rj�<�:�;2m4���<K�<=�����$�h5=5�,=h� �v����I����맼�5=�*=�;�;7:N<�������rZ�fv_���=�=[��-��İ��9�;�%�</������Fwؼ"R�<���<^8'��5p<��X�����[��&��`=�:=j;=�2��X2g=)�-���8=��d=�ؼ�^<�M=.ғ��7G=���!�=��'�u� =���:j8�;p�P=N���d��<ii0=:T$<�A;@�ƻAcZ���	�Z��<����/�D%X=�C��xF=T�C�GkJ��qU=}v=4 �����<�!����4�O=K���7(=Ttټ}�"����<� ;e���6�<����Չd��@�<�}�<��;��ּ����%�`Km����!�-��:<�Q��y�^j<c�!�B� =�Ȉ=I=���[==glR=*u�<�%]<X�_=�ڄ��A�:��=0c�<]��<�wA=���	�=h6�<���J;���W����S���r
=��w�+=��ӻh�0=W�=J;V�~�<f�:��=4��<XF
��\<�W=�2E�;��7={�<�e<�V<��<��<��F}K=!bǼCW<NH���b=�PW=Z��;�����.�<8���/�3���p�����<Q{����}�I���Q����|I������@<3�X=5۽�p*ؼIܩ<��q��N]=]0���^=���W�_�a�D��Dg=��<�ګ;�Lq;G5�o�μ���ڣ:�O׹��f=p��;�QмbEq��5��g	��
=a�'=�T��� L�H�4=o;�es�wȇ��H��F��-N���_=0���;a�"<���=S��F=�g��-r=��=)�?�r���Vd��Xa;�x�;��;�YF<�}�O�B�f1=�+�A[l���<�n8�b|�;��<P�ό*�n^K=E�B=0=�,����'=����:�<f,ݼ����Ա2��MN;B��h�<2|��)��<9U ��Y�w�G=d���"�!=<}���o����| =T�=.6#��=�|=g�-��{=S�]=K'=�J�l�<(鐻C�;�Z�P���gԼ&��<*���t$=Qo	=�n<=�o��M��<w��<���:��	��є;�E�j��m���s�<�t#=b����o�<Dw=���<��<�I���#2=#'��b�<ig�<j}>����G<�3��)��;���<c>�X�!=ğ�<(�<ܣX��P=�a/=�%E�YD=�6����;�;
k�����X�O=����Y=�I���-y=�@$��Rx<);=�3=�2����<j�;=u|<��Fn<�h���1=���;�A2=�/�<��h<��f��߹$ǣ<��<���~���x<�F�E�u=�=��*��[��=��=G�3���E�����N<Э<�}^�X	�Cg�<�&v=JE=,?R=� Z�_�=b�,;��<9^�;���l��[ :<B%u�������02*��\�B ��]=�!M�����
��}�=��6�1�`�-1=4 <Htx��O�<��Y=J�i��@=���;z��<Hyۼ2�#=*2&�W�<o�o=��*=��j=�y�n��<��!�`0%<��DX<f�9�c[<{��C\�k�����<@���#�;kE���Һ�r=;K¼u<���<���XCN�ۚE=��V�5:}����/vs:�cϼ1�<�g�8x\R�V>0=�w����<��=\Y�<��=z�>�������,�n@M��>�a9Q�N2�HD�����������L����B��/<Q�=<���>~<�ŭ<l�;�<�:r<N0)��L+��m����<�"=P'ܺ�9o;9���w|4=B����'�bk�:�N�;k�<)�<���L���A���6м��+;CA=,[��w�<Չ�<�hM=�Z���<?߾�dOD;�AR==V��w���1g<!q<���׫˻虜��Ao=�{u=��,�V�7��f<�����V<�6���=�<d;�<=O4���<+��<��z<�#�W6=��=�`U���<Ǡ'����<�_	���6A�<q�A<30<�%���ђ;}g˼�N�V�o�[^T<��+�S���Y��<��-=c@�qJN���.=�$M=Zk��.��<��c�Z8��X�r\�<X{5=�-�o<W�7=��=���74=䘟:�2���
�m�F)=��=�,��8}�� )��K�<�<+��<�9=���<[��<·==��3;x����!μ))�h�	=w�^=�ռV�P;t3R�J��<�\��i6�W��<��b<��h=�hX<U�h�<fd�<k��ɚa=�.��8�a���l�Ʉ���:-<��=����>�;��=�h-<�N�&����û-�*��i�<q�U=r������<�.<��E����<��	=�,=dؠ<�f^��Q3=q��<:�*���<
K��뼮	"=�?�j9Y���*�^A2;�3:�+|=���f�2=�^�]��]��;?e-=H��<�g1�),H<��b���-<B�����J���o=��=�n-�PwQ��<�ny��k��=0M<��ϼh<��ܼ�$l=��	<��O��>n<�X�a༏ݾ;�T��N=��N=`>~���7��,����&=�ߏ�I<�lH�*:�F��<oP5����9�u߹��W�Y�>�Ӹ����#���=�;c=e�ɻ-�1��᯻O�<wn=���D�dR�=zz&���-�y�<?��;�L��/��F�!���;<gd����_���K��[=I��<�(=32�;~j�%6=\��w�e��<o�K��J׼;sƼ�I�4��<�>�+�	��ӓ�o�@=�<h�6<�7^=���ECB�:�<f�@=#�I8K�8=
����\�baM�y|�0G==��D�
%�;�Y�;��<�M<�Q=�=.=q�3��YM=��c�,_<�dNH�B�=�%¼c��<nc5��[��x�\=��l��<c?<h�=�� <O[��<!�;i����U=I�<����.=��� uC=a��K;��h���;FR�ܴ,��w���ؼa������D#��/O�;��=E�=
�B�Pc�A3d=���;�6�;�:�A<��&=�9=ɇ2�jS�j�%�Ɠ�<�0Z=�e�3�2�?|����:;|�<a���>OJ�����������ڨ�HTV�R;�o�;�<J`<k���z7	�%�=���l�;Jn=���;�(=\�
7�[&=Ҩ�;�+����;]H�<pZ���N��j�<�X�<��>�(�X�^�R��������|�$=<o!�g�0��$:�0�=�cżi�<y��]LU�@c�<����54�3���#1=Jh��y=� �<���<Q�
=�Bg=�1��{=�(;���<���Eg;�+g�x�U<,:=k����iŻ�h�=��=�H\��#����<e�[�� E�\(������{��]V=�]<¨�<ʫ��@[�<�R;< v�<���]|�)�*=�8=�=��C;���;N�1�Gۇ=Qo]��a��h=��뼚���*C���&=wC8���%���P�%���G���s<j�<��L=�5#=�0�y�<b7=�Nv�b9����a=�<�=�|9�����2;G��<x]#<�&�Z��;'x<�0=����/����?<�@�ly�;��R�$��W�
=�����3�e�ͼ�᤼�M�&D��=�x��q)ջ�eG��R&���@��`�͑�;��T=�zp=ܮ<�+	�M�=:u�;5T庳jC�g�������J=�����g�<��;=/m�<��6����<��<�~�;�!g=�	m�$���A�/�O]⼊Tʼ��<��=�|�����<���ӈ����<E.��0h��d��5<=Ҷ<����9��<�;�=���<�gn=�=X�8<�)7�B�=���<q� =<ռ�#���뼼s���A����;��A��惻�(���=+�S�:��+,�O0߼�b��I=5�t=�C����y�9��<�">�w�<��5=�S-�|�Q�[;=�O�<��m��5t�缅�<�߻G�d��p��-�<�ŧ;^f!�7=/��\܀<a�:i��<@ͼ�P���v�=X_����%��.z'=C�<�D��A=�f5���'�ZN��zW���@=}w����E=bs��r�=���<@%Y���ȼ�a_=�0=���0t�<~��� �;��X8��|M=Ef=f�@=�hܼ�m��J���)=>�����=��k�Iu=9=��r��I="����u;w
!�w�<�P�<n=�<�}漯sT��E�;���;���<	��<�\�<��j=#M� *t= QI��j����!���<hw<m�t���:<�1@�5=�<������<���?��ߴ�����<��T�� X��J����:=� (=1U>=Iݼm��<P��~�����<��O=m���J	=���z@K��,���)��j��r=g� =�b�=`�ǹ�G;�J�<��E=��1=��48��!.=.W��=�<�H3���c_���	o;^l��B��;��<`�=�R��� �a������h�<TA�<��@��d=��!!=AМ�A{5��wb=����@ռ.�<$�༱��7=�z�<��<�����DX�;���l�M�Q�G�<d����T��+0���?=��<q��b�::��<�V=3�;o�P=�jw���<K�\=��	=X�-=0�&μ� =S҂<>^n��޼�''���:ޅ=�3=����į�<<-=�'�ET�;��;�m�<�ǻ�c=�?<'����;�%g�h��`�PV��+�����)_:j�O�S	�����<~���s�Ƽ����Ģ�Ķb�#�;4.w= X��M���o%=o�=�;N<��<?��2�G</�<�_�R�R-�=��8=��<<��!��V�"zL�t���(I=��w;�����l�I���t\뼋�=p�C=6U�E�!����K=pN9=�x,�$X�<ﴓ<�=]��=���<ը�c�=�lW��~=�D�<ʣg=�=
� =o�N;�%|�UĻ8j=���<�(�<(5	�$�����;�8��GP=��l�QRI=(�4f׻�n<e�S�z[�<��W��^<a��[�@������H$=5�i}}��e*;�ͼ Q=a����	߼�IQ<m�t<�*<<�쑼�͋=4� =W+/�ȩ����)���=x�<p��y���/!=����?�ϫ<��<�M=dQ.=�#$�H�<���$ɻx|���46��/"=��:��9���b�<_*��B��#=ѕX=2a}��;���<X������*y���������:p�<��_���?������<�Q��%�<j��<��==������:���<BZ�=t�`=|������;ezJ=������<�8=�nU�1��a��<�� =�VP��ȼj<�=�
��8\Y=� t<Vm@�.>��""P=��^�Y��<,L�=|W����;T^�������<4;S=�׳;�!���=<�R�a�W=H
�d=c��9j�<V��<�'��PC3���v�n6.<,T�r<�<���<Sn=�ņ��[x=$x
=͗A=��;)����<�F/�Ǭ�[����i<�\��<L�s�
�<���<������1����;㫗�XU���}��!NA��j�h��I�i�;g��:=��M��u@=8\9<��;�L�<ͯ��8�*��um���<�E����<p�	=S ����ĺQ�,=����	=納���O<�J;#�m<pf����)=O*!��=_2$=h�g<uS=U9W=U�p<=¼�+=�#=zq\��� =������O��kn�<��!=p�"=%s+=MQ��
�	vS=˛!=�6�;_�E�8j����޼���<��x��뼯A���<�C�<��=ݚ����@�
���=[m.=��K=|n<�a[<�p.=$��<e��఼��^��9C���a�|�,=#|�Db����<��j���<�#̻�8F=p�{��qm�bE3=/*��ǈ=�,��jU�<D�w�w==��������:==,�=:�[�An
=����*��p�-���<&�!=2}�;CԀ;v/=ͧo��t�θJ<����
=I�a��J<�3Қ��x�<}��<Jym����<4i<^@=��=A��o1=
/�Q��%�6=<�
=���<G�Ѽ1ZϼD�s�L�M���<p�!��tZ=�4�N��;*`�<�ż�hb+��&�ʴ�<>�d=�L0��&;lo�aE�^=&�M=�-`7�b�<'j=%�%=+B�<��<*�<��C����<bZ�<ux=տ���:=�N=E_u��KZ�e�;�����J=
$�=�M	�Ʌ�������ƻ�1��o7�=�Y� y<=�I!����;N�;��/t����:�~_��2��v+�<�j{��Ҳ<w��:��;�&�1��H=P �kM�<k���� �%lL�\�z;a���f;�<ي=�L�h'�mrb<����S)=v��<W������e]�p�ü�4�<3��X������6>=p7�O�e=����i�)���ͼF얽=���<��(=;?>��$���5�B�:-=���<!�Q��'�]�ѼĪ�Dk�;�j�< �(=V�	=j;@=���;���;z�o��A���$�������W���⸼$<J�x��<#ka=�7`��S<�AE��@=�����<"*��-y��j�<5�4�2q+��/<����<'0�C9+��6k=	�ʼ�=�<��i=��%=��<;�)=��0�oڇ�?X��v[�<�N-=�e�,_�;s0;�6�@=8�
�1�=���;��v��Ǽ�
����
 �j��a���!;Ke��aI�<�����2M=�� �������m�A=5#�շ���2=%e��I�z|��b޼'��x2(��?=�k�|�׼l�;�kB��:�<����t����:�t�<��<����������K��<b)��C=!
�<2�Z=��x=��,=,N�<YO�Z�X�V�F9��<��8:��,���J���:�����-3<Q¼�7X��x5�G�ż�=�-���}�����;��I��ʁ�|a�=p�8\�=� h=[����sj�T�K;`�ȼL =�`�;���Y�
�uy���<޼(=�4m���<W20;}�
<�c�CN���m8<S+��^�;!%��f�[=R5=�;C<�V�=~^=�0��3缚�G�qC�<'X!=���:��D<+ ջƣ�U�E���N=ǻ��s��<�1=��`%=O���v�����y=�j<=�/�<2���}
u�4�4�L]=Ա;� 3=v~F=��<��=��;5�=��<��9;Z�<.��<A3=q�I=40=qڼ�}�>�SO=���;֛�<r��"�F����;��b<|�9=�3����<��H��=�!,���ܼS�n�W�J=����׽=Pt���v�k���Z.�if���;<&��;�?㼙��<\�W��`�<�'��z�:θ@<���e���?Y|=��=����&*� ��<�_�<�	�º��^�<,枼��n=�B=�z�;b��<��ʺ�67<�T��f漦:=���?�O<m�p��v�<fe̼�$=�	��( ��	�����yY6;Ke�<Xϼ<r�F�=��5=���:�I��8ޕ<�� ��뼼.��rV������<��'=�um<Mߚ<��i�P,���»��=h�(=;���脼ƅ��L��Y�s��n�IQ�<��t=մ?��xi<qD�=�Œ<~=��I=~�<�!*=&�Ժ��=�_ἜX=�LQ=��<�����=d�<�緼C���768�������<=�Y=O=u���q=��r�^P�<(����g ��N�!+���Q.=�m���I=3G?=!�2�K�3=q:�<��=e�+�;t>;��v�<�&��`��L�;5�'�%�Ѽddz����Bd�v
��h��jE���<}�D��_0;��-����vU=����-+�v�F�{L<s��-N�h�O�5EX:Y.=��&=M$�+�V���a=��=���<̇�Wwʼs��<�=�<>0�<��@�o��<��%<��:<�=r�&�_���g�C:��<���<yH��&��4��<�ſ���;�%���V���5�=["�:9=�?���%=I+w<^e-����;w%}�(��<�7�<[�2�<��R�<�E���$�+j;�c�c"�<r��@TѻP)#���<6���:�=�G�<����F�#<c���	��ZؼB�Z�a=բ`=�'�<1�S=�(!�X��<��(�ə<*w:,N���v;y�VK�<�����!����<-_,=��07=K�Ӽ��8��Y�V�=*ܼ�z������]�9�d�4��3a<�O(�$N�6`���=���=�4�-�j��=�Dr92����7J1:=����&<(>M;L�����<6�O=�q��B���T;�� ��!�<Td=�A��ar�;h{:��Ә<�����I<}ɀ�ʹ(=���Oɂ��:�����P�'=qu�:�~<��8= �=gxҼ/@=�:�I��<�+��bc=`�;�<x�A��hM=�y�@0�Q�<ģ�R�m<�R�>3���Y=qB�<�.H�:�������&>=�pv=Z�D=5�3�H�<���=��=J󐽆�ӻ2��_�X���=?=��J=Hh��OW`�biH='=�t̸|T=�v�<&��q=J^s=c��</�<p��nr	��ss= �<��C�.o�==�<��t�� ϻ��.�m����=�X�78;4���Nا�}�;�4=��v�K�:;L�뼃[<�E�ˉJ�l�<�Uq;/π���<��Q=���K�D=$T<==a=F��<��U<�&<T�K=�񼂹\;�����	�V�T�:]�I��P��_B=�E0���6��s%=��~<��7��QҼ��_�-�;2=���́���"���?��[�;���M���	�\��/���='��,h<��=S��;�h�;+	�;ۥv����HG�q�m�h�Q=�M;=��4�������/=����f<��!=7������DԼ`���ë��Z�<�D��P�=�,Ғ<�N�;���"��<��Ǻ��<�UD<�^<_@��s*��B�<�$=
A�\o�<�,�����<a<�f�<;�,���d<�fC<���<(]Y��������1a=��=�[������V(�nu����:��;$<�4���e=��$�v��`嘼V�+�28<lP�=��=W�W���������T=ӝ�&b������[�<NU=�9;g	O=�~2�\ <£�<0�g�h[<ߏ����!�7��ѹ;��T<�-z���ۼ���<��=ԍ���;�@6<�W��#�=at��5:ü����v�<��o<��'=4�1����<18��#��͂�#���B=�O0=I�<U3�
G�<�z�9j����[P��Y�;�����؛��=�EF<���<A-8Iؿ<gQ�<*�E\;�%u;H1v�+�D�L�J�6��<m,�<]=_�?D=!�7=���Dkd=�o`�n]2����<���<�O�����F�C���<�\= �q=��K<����D= ����<�K8=W�=~�=`,J�/��S=�����.�Iw:=|O�p=��O��#�<�(�j
=�^f�P}=�U�4KG�b҈���h��n�{�A<qn�~Nϻ?����)�|�T���<��4<�fc<W����=����"��]Q=.�&=�i�<dx5=��Q=r��<��Y�׈�y6;�2=��=uq�;:Ǝ�,&����?;ʛ��X��<'�M=�#4=�A���B�<!|�<��r��f�<�R=kU��#b����L	�< ������Ih��)�;
?���^�I�<MB����?��J�@<�ޒ�|<��;=xZk�	}#���z=�';/u=���;�I��F,�N~=�qQ<��9<�1:�Vkt=���]�P=�:�;��;��=&<y����o�O�����E<3�"��/B;��|�"�U<�Z}<b��||`�"���-C=�m���oz�<1<��:jg<=%�P=]�����<=��y���<>ZӼm��\@�Ԑ˼'7=L��;��X�/�P�3M��='�<���<�	(=+M;�<��{�^.�:��A="����&�ˢ;=������.��F=��<f�ټ�j<(%<	���&	��6l<tYQ��i�<Rq=�I =��̼a!M=P0��#d;��B�O<�i�<:�6�"�0=�߈=q�<�$w��~�<0���1�z�+<xPk<6�4<m(<��鼑
=�_&;*�i����<��3<d��<,������$ʼ��<d���T�<���9��ش<Od�<��B��z[�S�<{&�"�.�@0��A.�;!�_=�ύ��l1����UM��Kv=��Z=7d�<R���ow=܀���@=����2=]�=���<5Eq��G¼�=��=
=v3�5O==�ɢ<h��jG=<뎶�/�x��u%�
=��;M�7`Ȼ��f��q��CH=��0����:��q<�u���(O�y��7�[=����Jn�;�l�"�F������A���Q������ټ��g=��=��#=i(=���p�/�@�X}<4�=-?<k]���*����<<�Q�D�(=^@���}='����R���_=���;��S��=e������<�|M<�2=g�P;}�)=�}p<�z��Ii�W�-���=����;<�\=��#�ʐ��z=���<���{ɼ�D��N�;�p�:��<'o�:��]<D5��* y�
1<!x����&��k$=v3l���e<�4�<Hh_����ٺ<v���u����J�0=�aR��xG��༺� ����k�`V�<�~G�"p==���;}�7=Y��<Q�`�S=H�V��a=�<�i�<�x�<N�\;��4=(��)�6<S�.����<&��#&5���	=��<��<��-��[��v3��v�<%�<�/<�[9=[u�4�<�a'���<�"�<=K��_�r�<��=Ga �Q�j=��/�Ǡ��UV8��u[�R��<�y�<3�ºe��<F�~<�Ke��S�;�)4��6d;BD$=7�J��؉��v=�~=���4< ��o3����<��*=y9ɼ����]���5<B%:��>4=�ҁ�79=:���9�<E ���{1=�4��R��34� 2&=Uud����P�'�����_�D=�(�����\t�C����<x��=:x[�
�x���߸�E��(*P=��L���ü�z��n�;��4�z-�<�TI����<�'�&��<Ax����w=�u�JsA��W�7w�<+�<o�=�k7<W��X�1���:3]��p���<[�=ς�<5��e𭺸�K����=1�%<�[=�=s�4�)��_��<M�(=j�C<��ڼ�m�<��x��堼�_ =���<��(�!�̼��=��#�{!(�	�'=�:'=!��G�<�"�<�^=�3v<��<�r`=8�9�5m�;
�<?G��S0=��%=�i�<��4��*���gX=��8�og�9M��9-��J�wB	=|p=�=z�d<��C=�r!=�)��O���)��0=�9�ϳ;�{N=��	�J<=Ѻ=��6�7�]��<�k�<VD�ų�<}��;O�v�6��<x�@:<$.=~I�<���E$=��I={�;Z/4��k=��Ӽ�==,0C�R��-G=��ϼ��<�mV=���$��<���ak=ţ��;�^�!U��`;���8�Ȧ =�츼�؊���6=�k�}�m��'0�)�]=D{�<������A=a<|@b��ɛ��0�<Z��<Ӆx�X�j<�aw<�
P=�.s=K��L$+�}��Q=L�<����.�=�<=#�R���n=��Q�=*�a<�Ut=;��q���&=�x7�ϕ
<d��;�)��W�=��;�R�_��W�:8�=Ѓ����߻u;�7i;��J���V�%��<u�=�=�v[=%q*=���<�� ��6�<^��Tj8=�M��!M=_����j�1/(=88Y=����;��H��<��=
��<j�/����&&<�F������ӻr6=wy~<3`�}	�l�=�0r�J�==P�c=C(^<NCһ�C��m��n��;��W=����n���h��� �}~r=��'=�tڼϵ���0�|ӺP'��N"f��=w�����b�=���<�|L���(=YH��ę=q�	�z�/<��^��4м�`ؼ>1b��L5=��_=�1�<�?�9�޼�|M�Eؽ���5���
���g�Y;��=r�E���<�<��l<��=iQ
��ʹ���<Q��a�6��:*<u[T�Aw�<
���C�<R������<�����W=CI:��OQ<��>��c�m$�ό���	=��<�1=�P<��꽼�H�;Ґ��·<|l=6-=Ś�<z�7=���[x/�=�=�yټ��/��:=>Ұ;=CC=}�<6�y<��=���<�hE�X�<�=�@:t&|:��;��N9T�伉��<�29���<�Jc=��29�=8=��x��\�<�-���"߼/i��������� ];��;-��/ =Wg��=+Y�6�ͼ��;6�Ǽ�%��+^�(�<-RO=�������f��}<�pS0<.V=��L=x=ڃ��+h-=�g2=�I[� I6�P�(�&�=��;�Z=�QU=�X�Twм��Һ`�C�/�?`༔}�;��R<p�@<{6X<K�����<.U;�m/<�Z�<�E�o�<]T=���;[yD=�d�(��:�& ��S�	ŧ< p=1�;;cw�����<)»<��3=aN?�C��;�7�˞Y��Z��=e���x�I=�h��e�L��8��/=��M=�׶;n��7^I=��S<ФM=�1�')=d�Y4�j��#\�=E�2��лֳ���<ϼq"'���<������<�O;��R=B�;�Li=kn=��q��7�<+�<�r=<u�;�����^8=`}�<��=FG�<�����U���C;�Z=y�=km=�w�<��a���漶L;�2s��3ͼg�Ļ�C	<G���5���*5����'-=2�=zA��'6����<��C����<Ŕ�<��A��P=�J�.uo�Y&���e=���<�N[=f����޳=�����V�P���-%v=��n<���m ���S��wg=_��<���:}m̼���<Bt<�	� 2	<�,F=�>Z�$&�;a=�dp�ռ��X�L�w=�5,�R�ռ������<���<8��uMO��St=��=���<�;�V&=�-=�]'���޼�~I��Q��l�;���*<��N����<��K<�?*<q��< 
2�N���ړ<�~>���2���#=�=T_}<~�=�u����<�D=��X�UF�;�Q�<��]<�3���5�|��8~�r���-�Ն��#҂����<�K[=�_�΋H=��^<�D1�k5���8_�9�9=�8=�!��A�:����<7=���;IO�=���F=�%b��]��x��=�J��=�i꼴D8�t��9@;o��� =�\�=|��<y�;ҕ<0�v�w=�=b�o<�T<�i��@=��Ѻ$��<��I�npJ�ܝG=_�߼0�D�����V2R�~XҺ�&A=Yj�<��<�v�;�Z.=}�Y�6�t���W
=��M=]�|�ǻ��л�W;��x�d�s�;~.=6�/�UH=�>����=��(��QԼtT>�^�Y���!=���ܩ���G��ܼ��=ͼq���Kua=C"r�I�,=FV��p�h:>s������e�"��<McԼ�4=!��<�ş���5�޵�j�����FZ$���x��,��������o��O�԰��u��@�8��U�,�+���y=�uM���Q�$�����8E��R�=*?=��ļIW=����Y���u=o�c�y� �K'�<2	c����V��<Xt'<�,A�|� =x��<%���}�<����0=�EF�=����KJ=�ƻ��ؿ�Ս���==`J�*�����d�2=�[*<�	G;d�<8=3o=���)��<�\=1���]I<��;S	A=X�ּݼ �5=�]��>�<�֛��Jt����c=�,;�����(g��+��I52=>����A���\�(\���;=��=2�¼)�;��</m2���eS�<@>��n�<�}����<��I=b,ػ�=��D��`���'��Ȍ<[�s<� �ZI=_i=���X)R=��'�34�:��h����x�=���;=����O���9�� �9=�����d�<�����Ⱥ�"߼�d���9=�Q�[=�6#�s��;8h�<��<=�����*�]��<\���<6�6=��l<���<�Ւ<�\?=3)=�!��� ���;�t��l/<�)�<L&>��<�mw;��T�����>�o	���мG���$���A;�4=�'����<G��;k�<�{C=��>=sI�<���< p�S�U=i3�n2����#��8�<i�5=`�=��ی��"*=d�8=@�=g�<�М�� �'{=8��<�*O��G=Q�?�W�R��Ǽȃ<�y�^�&<�߼_�&�n�:�t}K;����7�<_G=�Ԡ���[^=R���<�G=*��<��e��a=Iy�<c��<KT"=���<�{�;;���D�=�(=�J�<�e =����9k=�V]=�u���|�<�V�<��C;
�[��n=��<�0���
��c��u=0�x=�*�<��:�HV=F���.�<6�,;%�L��	�<XZ�<��� �Kx$�P�j��Rm��:�.�:���<���eON=��<5 �<na=��S��ߎ:�@���x+=^�l<�L=P�;ۣ��[[=�g��i=C��;� =��H=�����="���Ff��^'=s�c�k�׼�	ۼG��X��܎ؼ�H��#=���;:-=ͩ8����g����6=4�|�U�;�٬��o3=�*	=���M��������ܼN�w=e<=K�C��E9<���;E�S=7D}=��:��=��n��=��3=�z�${=�"7��E�?h����E</��<;@><�g>���<0h"����S�)=?��Qh�Uu%��#a�~v);ڑu��S�<E�=[{n��B����L�*�Ӻ��λC֌;ki9=Y�<�| E<�@��e�B��/ƻ��-=��<â��/�</�Ӽ�iK=z�*���=C|�<P�D�B��7�<H��;�G=�=%��e_��et�]
�<gZ= ��<�;�7$��&'����!wQ=#�
=�B�}����NR=g�J���=��,=Yg��ӷ�3\��/��#�˻)����hB��f�=��=��޻_W�9�+=e�9�g =l�|=i�<Q#=�#;��L�b��;�P���=�;=1dq<�\=���p�+= ��
�<��%=l��<S 
��Z��q%<�� =�Ҽ~�E;��M=�Ea���;=�A�x�=$����)���Aջ�u޼h�F�G��;{8�<8/i���(<�Q=� O���@=\��<���<��/=�t�.#=DfB�,�=��<�7n�}����<��I=Ғ�<���1���t@=d��=�����f�����3IT���=���<��8�6��Lڼ��<D� =��&=b=��:��d�<��<MO=�~���=��=l{,�r��<;f<H<�<��
=8�<�==t7��,��D�X=��<v�:����6N��`=7��nB�;:o��t=��w=(B���R�G;o<Ɩ�8����d=�UN=�7��L"<���<��a��7�<Cv��;��,=�<Y�W=���͕���Jt���O�+xb�	q=ʽT=˾�;\����)<�kfW�!O��!	��i��<�c4�/�<P&�:m<2�d�o��<	:�<-��g4�!�;�;��ji��%=�^=F�9�xǠ;s�=avȼM���=�^=%���D��j��k$=m� �=ѦB�5T=Z��!����Ti��/�˧=�K���=15�<Aw=��=(�D��y����==([<�.=!2�<$��ZQ)=������<��R��<�n����:�����2��A�(k]��N�d��;��<��<�Q=����<y��s+�<N��9�^4=�I�< {�<m��<Ϣ�<�5t=k ���<y�=)uz�Ö=@�%=�0�;�F��.���j��#��<z8=4tk��)	�p�2��Y�I~=<�Y<�@U�����ub�<m ]��Ro�J��<���+�M���6=��~��P1=�ױ�#,=XA�<�IҼ2��<.F�<3�^=�Z��[=Z��:���-�k����x1���$�<�`�KC9�m��p��;K͍<נl��	��s�*V���N�t.;�1�m���_���l���z;1*s=����޳Ӻ��=s�G=d�x�sI��DhL=�<:��<�==�'@=Ͳs=~�=��4=��f���$=$�=^)7<�&=���<q�?=?{�<(;<� �ڟ%=�:~���=� :=��Ѽ�e[����<RF{�G-U��R�<�4�<�<�<�W�<�,=�=�6$�7"���.<%e��O=�r�=V�ؼ[;g�T�S<��<�>�ަ�<�9����<�K=��a�<��=�F=Œ��K�8�N=�����#=����n��մ�<�t�<1�<=����T9��2)���[<&Kk=(VӼP����g��Y�:�����E����=г3�f�\=L9=��'=@��7'���U�+�H��k�^�;�c=	Ċ��5P�׆<*���%nW���(<�
����<Q�=�jN���+���@=~���!�<���<��;��$��;�����m��M=(�=���<�a���K=�Ny;i;G� ���Ƽ�5�; ���t:=3�S���!��м�Wp��	9��%v��Mi=X�L����0�U=�R�<y	<G;=�韻P��: ?�<R��<i�6�m8�<�_{<�0=qp��� ��)��z<c�ȼr���s��<rS.���e6���c=@9K���'�k]4;GK=W�B��^��0�=��<PռC���^�`�;���<}Db���n���E=n�=F%9�7��ܛڼsT�@�캕�=���G�q����f}��^�F�,����<L	/=ݎ/<������=�Z�;�q{<Ч<S�ļ�:�<�N�1`�rw���)=��;e���$�T:�<��k={���G��:K<�<`";ρ���W=��H��8=~����<�5缈 `=��:�o=l�<�_�<~J%�j2��|����~�к����8<��?�5r =ɤ�<Ce��͙�<�W����>: ; ��;�0=c"&<��\=VS+=/�/@=���<�#�[��<��4=j�ּ��5<�.�;��D=�L�����s�3�F���x!=G�,��R�旬��}����`��8��
�<�8ü..)��}}=t��<����~w���1=����x켽�=�9=i=}�����!=Ņ?<�()�p�=,�$7��H=��S��I\=��0�B�5;T&��U���`<��żYW<�v=�WǼ��n<��߼���<.�� =��n�B�X<�=�Ϡ�㯃�u��;��k=�����h<���<���0ٲ��\u���=5$ʻB���
<��ȼ�u2��G����z��|<��@��=��189��`¼*으��<~�T=�͜�u}�<S?��:=�ѼQ�ф�i{¼|�F��I;�b����\=�vL=�%��5�e=]QZ��yG�:��t��؉�L����6=�����B����;�7{=�n��j���%=�.2�'j(=���<1:ʼ��;��m=p�=��<��	=&vܻ#����Q<�������<b(9�Ch; E��/��\;�G�G���V�׵�q�[=��;竞�{�<^U���m�b/8=�u �jD��U�-��׼�r��L|�A���V+<���9��=�����<�. 9}�=&�׼��⻛}=�T=�&�YXL=�6I<����z=�6><�3\=D�3<�B"=B'<^,�<Mq<
~0=��;���Ǹ�<��K�����m=��Z<�+=k#��e��l1X=��M=	b����<�U=6cؼA=����~c=�a�;�a!<dl�=���	F=;�=���;�t=�-B��h �k�G=("=˝���2�,�}=]S��{k����;�����,�浞�a����ݼq�G�frB�z �<��8�h�=ϯ漳b�=��C�;/��<���<��<�e��N�׽*��1�z4#=8�ݼ_1��4�V_l;�vi����=~JǻE��:2_��h��;��8=�/���=�����r�ۿM=\4�<L"==�D�6p�#=�� =0�<�
��-o�<��� 5�5%�;�l+���h����<�ň��F"�ОN�r�����k=�30�:��<r\J�P�9���W=G��:��~=�IU�CA��͆���k<��)�t �K�5���<��̋v�I�
=�R�)-�����~'f<{����ƹ<0�<�/�7��<q^Z����;Y��UCW=�P�gV�������<�S9==�2=�޼��;�ُ��l��[8��̱<$�e=�2�K� <�N=����<�ۿ���<i{S��Y�<�B`�i$3��.�<��B���6<�vX���'��W(���;3A#=�U���#<�*(<��;h��a�Ի��9=.x�=zIL=�Q�����Q=L��<��=�e<�o�<�S���r
��һ"}?=h:�<R���^#���1��%�	�;D���Vꢻ�	�<���,ɼƷ<�Mμ�U`=�I_�g�=�'o;�&&=�C<���:�Q�<�:���u���[��p]<��E:)��T����8����a"z��S=O��Q�[=>���T�����<�kܼhv=G�z<����=x�3���<��t=�+=(l�<W)=�M)�n�=wd�gC�v���k�Z=�\`=�`ټJ�ϼ���x�a/���}� �8��H�=N�ڼ�q0��^û& ;�b����e�6�<�)G;E�K�!��Dc9��b=3��z�O�R8(��%=QA��<�
<B=���k���0=$�=��'<$���],��Ђ��,b��=8�}=�	ɻ���;%;d�ɓo<�LT=vt�<0K=���:JJU=���� 
����Mn�<WW)=�D!=p�!=� �;�ߗ<=`+;��3=����m�ͼخ���*��}<W3�<R�=͢B��ꧼ_��9o=
�Ѽ��u�⎚�[��J�μC��<+�;�&��(F��!vN=��b��;�9O��!�<�S"�.j0���7�mG3��`ܼ�V���'!=�FE�kl=͔=6�˻�V;|  =#hT�����{p��皌<%�>=��<�J�<���<u_=�E���<�@=ڵӼs%��)C;����</~(=��.�G=@��<$:��O
�Jj+=,�!<�XT�4ļ:�]=�=����O'���}<�=��k-�m���,u�η�<�|X;���d�;8��
�s�w��m��Ƽ6[��U�f&�ߕ������n��w=H�<��׻9^�;�Z�+v@=�킻k6=�I�<�����`=V��Z�W=}B�������Gͺ3�z�9�<
U� �S�A�i:I�p<���<���I!=��{���<��&���1���ϼD;=�is=�A(=�r�=��f=HE=�$^<�E�:�X3<�`���O<"X�=��=�!`��:��6�<%DR=^������S=�����G� ����?���#<�;|�{��޼�(�Y�s{@�pK��8���G!=h+�<#�<<��<��3=I�W<��|=2�<H�Q=��@=]�x;,�/��C�<��⼔]B��Q��+��FD< ��v,O=77X=O�ﻚ����==2�L����<��<oë�
��{�T����REJ���.�[��<j��;S�:�N��<�>ɻ������r�?�Ѽ<,���F=�⾼Gs���q3<�Π<�4��E#=�O`�WƯ�2�=�姼� ��^A��9����#=j�<!jb=�b���i��e�<ߧ��C=A�V=٬���a==v��	a��.�<d�2�T�;��3$����=�c <?;<-R =Y�1��<o�k<�1=���s=td=̼�;=7��<C=�<1�� _=-�Q;����=L�R=&ĥ����DN�@ O�2�(��#��4��W�X=`�<��*���Y���	�c��;����j��i���=�<l�,�O�T=#�h���<9� = ��:�r =��"=*5���0=��ؼ��I;{�;=n==[�5=��M=|h�<��<�@�%SQ=��!�	%(<�O����;M�9=��o��:5��v�h*@=��<T����q/=wU?���3�X�<�_;�$B��e�������\�;w��<,�<�eG��6=�I�梔�.�<��o�Z�<.�<6��<Ê=��<̈��g".��<�<%}<��<A�����LӦ;ᆡ<�H<f�B��倽8d�U�X�t�
��i��w����<49=5)׻�̗=|�g=�.m<x�'�@B��	=����5���-1=��=���;N�$��H=���;cm�\kS<mx���c�b<ݳں�N[=T`Y���l=���ϻU���/=��
<fx���&�k����j��F˻)�<�/�h���	�gu=�W����H�݈	���`��q�;�>��� ���}��g=��8�ۼz��<����B^��},=EW-<!:=�$d����;o�ԼF���p��E=;
=��g�p^R�k��u�7�;E��=:<A�c<�=j=���<I=��g�dN�;��\�N�=ӞP� $#=dr�=��-��n������i;=���݋<��b���(�<S>={��;[��9{��<��P�N�׼r� =�n�����J�d>V=}u�<��v��J�<�ă��iżzI.��5G=�4=�0���)�;$��<�B ��L=/��<��<�V��~<0�I�[�L=#�<<�>!=����)U=�~(=��=��n�l�8={9�;Ҝc<��K=������8=+Ҽ�+�<Be=ΐ��?����Q��{�)��2g=��!�#^M��q���^R;5X0=�s�%��<�=��<�ϼ��3=�t��$��<6�<�P=��^=[�<�
��7�&;ѹ<�8�rt�<2x���J�=|�;�O����j;��x���<���;��/��̼F�ټZ�-J"�^�	���!�H�Q<��G�����N��Ƶ<t��<�c*;AO&�	܍��Ҋ�=���]�C�[ *�r㧼���<�e�vY+���!=�? <$=[��<��="mG�[[M=-�<6i�<��1��P�,�<�����=���<�PB��w]�<F�=�3'��9b����_�.� ��<�y��7�ԐS���3<~T=.=�/!<��=D3���=���<d*>=���<����?1�s�S��39=l/�OM~<�$.=����r�<�5=1�>=��<����Ԋ<��==A�=5؜<.�<~�i=P�P�я=����r�Z=|<Qb=#m�<O*���ż�w	�slG��'=��e�K,���̡;�ɼ��<{�T<	jϼ��N������v����)=�y�<��wX=��U<�X=�2N=j�:=���:�G����@<#o��kE�=�cM��j�;YJQ����<�P����;r����I=@�1�+Ļ:�Z�����=��M����;�I}�*\���A���v�1d=�o�<�)�����<,����=,}�<�'u�kQN���+=l�F��e�=���RH_=���<m���D*==�%p��FG@��B���<K�-<�%���L:��<��W<���<ǖQ=։�<�j4=�:�0�(=%I��
	=o�$<���<���!%����k����@ؼ(��;����׎'�kٓ<�OF��k����5����9��n��t�F=��=�?'��'���o����<~��<��>=�1�Bm�e�=̥�'9u�yxq��[��B:�S����=d�G<c��t=׾�:Ss3=t�=A�#�I�1�"^7�py�<H��<��=�z|=3F<��7�p�~<-ۼ$�`�aP�`ü�i;=��A�[=��E�1��ļ��F�䒍��'
���4=6��<�<N/�< s<c���`=���;2�<y��;����@=0�=���<v`�<��m=�\��-���^:\���	�a{O��=bd���e�$���iy��
/������,�s�{=�0��g��<�Kv�h�;=�<��#������c=-�1<�O<��;��m���K���<L�^=,ډ�8�ؼyj<=Zؼ1S-��ၼ�Oǻ�CG=�O�x��;ϖ���幼����ĺd���89=Z?�vr��B�9���v�	==7S�]�"��C=<�o��^�;��<�0=M���N����<��:������\0���ж��=�5c<6��<�Y=�s�<����Q�11�m���F߄��#I= ��<�ET<CT�������F�<���; T�a"e�_�2=�'=\���7��pg=��W=Gj�2]�=��q<�T���<s�R<��<x�!="�0=��U��`��Ԋ�<n&&��>����<=+�<�3�<i�2�j��M����h<�,�<#�~��� �� ��L!��j�(�/	T���G�ۚ�%�_=����}=�S<�;�.C����c�f<ޱ2�5�gR=F-^=$}<K�	�E�=#Z�<C�8=U�h=!�m���X�:X4�m0�&3¼��缗f�c�C�B����;/��<2�`=��a=��L����<c��=9yc=��=��_�� 4��ϼ:=}�F_4��?һG�=�x���軻�<F~�JSB<���<*��;t���c0=���Ɋi<�*���ݼ�j=\�<&.=�j̻�J<�ą��Xe<�4`<"g޼ ���� ='ε;WE�������\;
Dx=v�~���<��W<��<9�-=���=�`<�P��
:=��-����=^t=�h=&�S�t ��Y�`=���s���=4������M��<&=CΏ<�PO�N�f=��</	���+�D�;��:=w�e�����'���n��&WM�γ{�9< =K��<T�M�
0[<qł�f"�<mT�ǀX�z�;˖ü�Op�f��<y�鼧RҼ=�;=��{@^�Y� =�(f=���H0=���;H\=l�0=�9��Gd�T����%;��[=v�;�3=b�
����<�cT=a/�<�.�<Ft��� �< ]�<��伞)���E����|�<|�X��<�d���t�e#v<��+=�u�<�&�����g-w�Ys`��4=) %����XW==h<�D��cB�H:y<�|U:ay�<�r�<�%�T鼅j���(�ݔW���H�Uu�:-(L�:ʳ<<�(=�4);��<����bJ�=�+��v��<F]=p�$=��=���<�j����ϻ����4M�v=?0�<��=��D�u!=D�m=SGY�Ԅ =)�J���B=@��;��M<��*=#���l= �;m6=�W �JI��+k9��=����<:�V�x<�._�<�߼;K[=�=�j�:3]5����;Ifm;J)k<e�^=��y�����W�{=Q��93��-=��<��`=�฻s}�<�bQ��W�ㄨ�����3���-<�>�^�S<I���31=�K�҇�;��̼�c̼!DP=<n=o(C�T�p��,=[�<���<;j��<*^;��=�������O��S<3<i�`=�7=���<4�e="
(< ='28���;�b=O�A=��s=Q��<O�T<�m�N-=�1�<q�=�u�;�2=e����ռ��<��ټ5$<N�<ܶ0=�-/9v�s��=k�^���;=2�a<�-���l=V��~�<=S>=l\��PS�H��C9<_{ؼ����M��h��
=��ZH=�w�<?z<;o�g�=��<F�6;E):=P�2=4A3<7� ��"�<���}M�<ٷ�<�E�<�t-<-N��9C��펼�q�XN<W=����;�C=�l=7֜�ƈ����4�"3^�	hW=m�[�6E>;+
p=�V�:�"=�����aE���J��������:�D�0��?�Y} �@�ټ��ݼ�u�;�z�����<���<��&=�=��P�\�����<���<�B:=�C�О*��SO<p=�t˼�<Z=#J;�k��<�G<��K��UغEs�<�D���!��	j��	Q=9 =�*��Ӟ��i͞�,J=n�<�Z�<�F7; =D=�a0=H�<�ʶ�^����}<�=�J����;&_�:Q,=e&��u`�<2S}=�=ث=�50��/��?�Sq<�7&��� <6PT��D�<��3�����F��<h�=&�
��S=J�+<�3�}�c=<X1=#{�n��<�{9�~�<]^�F������<F�7���:��5����������:[��GM;N�<��[=�{�<�
����I<АǼ���Xwy��M�;�K�QXb��7�<M��:|�)��p��Z�Է�5��!Q;z��f��z���}���R{<�.<(�k�j�5�:� �<C85=�ɞ�<rȖ<�0�<6)^�=��+Ԏ���S<�#=]n;�%	����J=��߼!����� *��c�=��<{�	=��<P��2 y��%�B�=�+�<��<]� �x���"�qJ;=��<��߻~�]<�dR=zu�<rO�>�L=;��I��̓�4UƼ �'<�)��R���Vy��*k�}Oۼ 찼��컣|#�\���7m�u)$�ͳ=[��<�(�;��(�O'i�5�%�A��<*=פܼ�z	=ӾF;�L`�R?t�I���f�_=��Y=�pb��I=*v�4K3=�H���^���=��%�����c=-Y=��:=e�;c�f�"=#<�;8�l=ݱ<�<�<���;Ȧq���n=Z���X-��f�����w�<�<#��Sm��mJ=o���w����!��:$=j���Ц=�a3�6��<NV��Z
=ƽ��S�<<P��XV#<]~%=��c����<pRf�}�}�~�]^Y�l�j��	�R���y�����D=^)+���������;�a=��p<��ʼ��=һCK��a��%\<�QQ=�q�<3'��YE�V��<�u<V]���Q= 21=�I=
�6����}�8=��)�HT�w�"=���=sJ;�'���X����<�;Ҧ�o���c�*=E񿻻��<�31��Ф���A����<5�F=)�;��@<�^ɻ�A�<��a���'=G�C��0��Dq ;�	��	��Ap=8�<��'��)A�<@=3��<�����@�6GǼ5�3�2�Cx�H�Q�w�!�)Ȃ=e'�=��<� ��|<�z�ٔ�<������=�%�XA��!=��=+vq=T�@����<�C=��<Mb=��g��?��p]���ݼ�I�l7޼�s�<�W;5B!<2e����=�)�@�p���<��<9�<dW;��%\=�}�<�
��w5K��R=�me����<��9���y<�+ɼ!5�:�ξ��F�<��N,!=ܠ:R�+����U��bT=�+�<������F/9��<��Q=� y<���I�<���{�b=$Z��5�*<�U���޼)�X<Ba@='v2��:=��]���;[R�<��ͼ�H=�M	�r  =T�<��%���<�����W��੼s�P�&�=]�?=�=�;�둻�}H=�v�n�Ƽ/Ӛ;L�<��g<˳	<.�3= uM=��<5-�<Y��<�f=)܍��� �qA=��9��1O���<�2�<9�Y�Kk��<�ď:�W=_
�<���+�w���<� '��;=��>����<6)=L�F=�K=�7ɻNi=0�F��� <$��<J�Z�$/=s�㺝�
=*���C(���,�����'<�6�=��;��o=��d����<�."=t�8+���B�7��5�����h)U=Y\��*�$.�<6�Ѽ92J�{=<�@ռd�<ݱ8=�j���r�:��<��8=J�j��}�;�f=}�W���H=�'�� �5��]9�R�(��	<��a��\�μ��Q=y�)�� y<�Yh��@�=��I���C<ai���:������қ�|���3Ɏ�!�=�Ҙ<�f"=v$Q�W� ��B�������:6%�=Hz��#׸��7=Q*�<HC���7D=7g=9U8=�Cf��)�:�]=ƧY�� ƼR/=e`D=�P �3�@���+=�[���ݻ��=YZ�:�!�eX��/I��$�<%�3Z	='k��0/��o�<(\"�ܡh=�"��X��5{=4)̼��4��L[=���<�x�"gq=���:9ռ�Q9=}T���8�=,N�S1��5�<N#�����ߕ�w�G;d�@=c��G� ���P��!�\���6���%<]�g�6=&��<Z�5=�x�<~����;����:R�<=F�,=�>���5�;�=�| =r,=��Z=��=v�4<L;<�<=�:�;���=��,�,���e�����<O���lϩ;���=8|T=ɍg�2�(��v�<����/��?,�5$&=bp4�82o��a8=l���mK�����0R>�6J=�ߓ����xI=�Q�<��=X����G}�#�p<��'=lH��-@=�q�<������E��RZ=_�=�_���V=i6=�1=k���^�;2���	#s���y����{+������Z��@ =�d=+�S����<��^�J물��;f�3��<O��<�9�ӵ3=����26=e�<��.=t���A}=��<�~�<��;�=��M��=g��<��<;\���L�o|.=��<bj��ƻ+/=eC<�p�;0�4�CL=$(�<7�;�H��]��M!��G�;�Pk��8V�0�a=#�;j�ż�)�<�C�1�<�\P��<�W�<�+(�)X���ݼ��ɒ:�mD��G=ɮb=R@G�k7=�	�<m=�|I��sa���O�e �<���<ͿM�EvT���&��[�<��N=��(���ػ���<�3Ѽ�e�+&��̽v=�l>=�	���-=z�G<�#J<>���_=��!���<Vk����<�&=�!6��2-�YŪ;_!j=��=�F^���J��m<�	��;��*=�����Q��ӏ�<]�Z=S�C=ZR��a+e��(c�{z�;fNV=�/r=� ���-���A׼���<3�T=��@�n+9�+�<���<�qv���u=���<�.=�Q�<Sʖ;+�=:6�;KL�:w�߼O
�<ܗ�3V���"��B8=��a�������fw=|�=����ʩ��f'=���<{\S=��a��2�<�m=D��<�(]=9#c�Bx���㞻���;Fm�V�\jH��6�N�漜�H=����˴���(h�Dv�;�k;�G�<��V��[=�y
���K�	��<C쁽�L=_�C��м�K��x��rӤ�فS��5=<>�� �:�B<J�!=��0<9.�.{�z����Z�S�==�9�A�A=�w��/�<@�X�깏<A�9<%�?=T�a����;������/���F=2�Q��̦<�ϸ<4�p=�~<=�Cg�~e<u���o����g����<S��1=8n=�B;��������P=�N�<v�Y<�s��w6����;6�+�-�<<	�>=$9＜�$�"5<g=�+=9���v"�@m|=��O<�?�<�:Z����:�Cc:��<�f��<8��H�q��ڼ�rP=R��[b9�Ǻ�*��U<5�?=�{��Yr<�9��)PC=���ͼ���.!=�aJ�O�N��C��T=�1�<��6=$�+����<�%�<�� =9}_�uI{��I�;k4*=P��=yA<Ο�e��<��
����<'�=��A��"I�;�Sv<	S2���8=�j�*�F=��+�J�=A������=jq>��1���=�_�=S�!�6��;|�<{�=��<��T���p��H�<�r�i�p���[�W/��韙������j=�K=r4;�׼���a��;cż�7���y���!<=D��;�鼾�����<���7�=b�v=�<�U�����2ɑ�#-5�}�a=
��<����v�=	�p<���<��w��eG=�e=��A=�n���:�4X�<p�}<�Ì<����L����<�p���)�9=���<���<�c�;T�9�&ƛ;̓:�/<+�9<]�I��#���X��<���9=�2���R<�ۼ��!�"t�<x!ļ�%�7�
=�4���%(�PN:}��<jV<�"�� ���"=����	j=��=1�i=Q:�<9vC�²S=C�K<�?c=�`Ȼ4�?�����<�̄==�<U"=�� �����	=�,=�q����;ߦ)=��;�N	�JQc=�Z��`f=K<M�ͼ>vO<璘��wG��F=/'Ǽ�U=HJ��{8�@nR<\�8��)F;33���[�<��)��� =�����B�<g#;w(�<_���:�U"=�쁽�Ǔ<�
�<�w�i�+��BF=6O/;��*��2=�i�<,�Ϻ	�ձ4���#�Z�e��u�<�d�1�|,ּ�����.=p4M<�F%�Ŭ�<J�7<for��J�+@=F!�P{k��؁���1<-"�#=$�`<��n=sp=jü�l����}<(+�4b�!=�br�aL��D=��#<`��;==�L=cPӼ��ѡǼS�"<�$���D=�0=��=Z):=Ӵ�<�={�����jм���C��=�6"<�ʋ�ک=��;���T��,��-�6��wp<�W��3;33=+�߼���=&�`���<T�$��1L=�q�gp�<ʻ�����Қ�8�I(=!Z=��<N#�<�Z�!���BnE��Us�b�=ιü�a��V\�H��;�������f�W���ɼ9D=\<��8�$=A�<s�<�W�8F�<�]����`T=QO=;z>���!=q7�<h�0�������X,�<��"�U$z=m!��,���>��u<���<m��Q�=)�i�1=�q�:]ډ�-<Ԡ	��4μ^Fw<Fw��`=��@�ȑ-�(��u2;��������[��S��<?Se��SJ�'p��]�P= :��͖�\��<��,=M]D=2hK��2Y=�tмfh\<�?�h��<�kB�k8�C���y= �o<���R�=Oኼ2[�T�ͼ(���I�<E�&�K4}:��#���<A=��f���'<�+ü�{�<{ =)�s;]o=B�R�:��<	}U�Q,i��w��X4<��c=�{A<���7�8���Q�!��}�776�ao(��C��.���=����<�m�<��2=�u1=��L�ǃ�2.#���&���;��Z=;�[�
�	�dr\��ID=�=*�<�g�;�	{<hr���=@=B$�;Zݔ�B&��~�:w=Lv���'n��Y3=*.O=���<��[=����>���'=����5�!�I��&�����<�f+�~NV<U	�^�k�W,�D4<u���C�=�{�<{�<L!���=Z�8�e�$����=)�n�=3;��L;��:�c�J��"=�&���<&!�	W���n\=V��<�D<�>�n�<{��=�=움;x���=�U��v�<�)�;m#<d��F�ܼ+5ż9>i��--<�y=U"=��$��1=��ܻ�=2=N��<��
�<�T��ȟټ�/=�G<���;�<���)E��.B�x?�X��<=V_<�
	=w��m$��x��Y^<���</H
9�lJ��!�<k���e=e&=���=�P=5�.;~L"=*�"�A=a�m<C��;��3=4^���-�s<({޼�<9C�<L��;�-��/f��A=��'�z<s�
<��|<(԰<�C7���H<�|�3{;��'���<�㦼{�:�(�'<����2���g��eq��q��<��%�S������0�<
_�<�<��=�»^Ђ��H={�^�9,o�92n=k�;1C���<=�O�<V.l=+s�<��5�
�=�������p'��g���;�8<J�M='Cy=52<y��<��,�E�B�2@=*��)�<��E�6/	��Q
�l�h=����q�<���� ��;�<�0:=�ჽL*<8л�-�<��?=��W�&�=S.�;h 
��{=�{;0Q_�ji��3&=�&��#Я;!o��=9b =��!������^�<*��;ytb=Kc޻04��<�O�f�~�Q�)�u<��?�W݂=5��<�T 8��ìD=�1y��5��|.=���;�/���=��<\��;x�<D�H<��μ)bY;��#<��i��G�<%�A��ª�A��<��<9�<=g#d���k=��Q����' =�� ��f?�}��<��;��=iW�<�z|������< 8 =���;[C��å�<G�>���2=�h���I�Y�:�9��<Ԛ��� Q��:I����<�������Z�k=�a<1����+���{������<$�Z�\�;�ǚ��)���Rc=��&��i����<l�@���%=��Ƽ1@<(���cT��E���;r�3=Iv���<�P����%=ڲ;<��&�KH%��=Y=��7������y���=���V{6�]�=
�6=��H=<³��<D�۽t�K,[��<B<�==a�*�4���]��M���m�6����<e�D<XH=��<M��;|l����=p%�%����<�ߑ;H�|��,ϼ~y=����P[�)��<b"<M�T���'�O�n��;�gP�A災��'��R�<�3C=�{�/��:��3���z���;~�O=�}̻�y�<%/=�����S���U���l��T=X$�A�����ټ'��<�J��_$=��%<A��u|��P�<�N���>���&@=��;�CW=N�7��A����<B��Z1�<r�P��E,�([=;G[�z�D=���<�;���_����X:�256�Ɔ����v4=�Z>��!;=mT�_�:��=P���?�/y���<��2���˼9=�V��_��/+=��E�u�+���<F��,��I�<1}x���!=U�<E�j���<~P����r���R�$=C�?=��=�Ӽ���>���\��LJ����~4=�bG��bg��Q�<>\};x��;[����=̄�<(�V��H�<�$�;TPD��M���J<0�f�~z[��qO=ki�<�1�X���.�;��;B�)�7�<��K��,�?��<���<⹗��s�<���<�<ʡ��xA;0^��T�<�8<{��:�Ӽ	k����5=���=I�	=�ϼj�!=��k=�7�5B1�MT^=p�=
TJ�N�t=�Zm:y����0�;���<�{��ܺ�]�<=�8�����vS�=C��;A�	=��L=J!=#��<�ɼ�6��D� M=29=kt2�����]<o=U8a=x�:�T�<-;=���;�2=�5D;ߪ=SΛ<�X1����;�F��t���a��67�{lX;�:=�/6�s��8�;�P�ֲ强����;�|�<�����j<z�v���O�{�N���Z���;�H^=���<�4<�[�*�<E+�!�;eI=�]2=y�C=mLF<�=[�g��W��;�p��ي��G3�8�����<�w�=��=�0;Y�<��<F�%�c�I<mC=��ټt��*w=�v<ʁa�_~$=�9=Y/=�X����<B���AG=ӹ<o�A�#p&=)��<�U�/��<�@�<�ۈ���ϼ,��<�#=���<����^,;$Z< ���� �1�`�ݕ�������6� ��<�Qn���=s�M�����;Gm,�A�Y=��J���7=mt=ja=i��<=E�0�S=�T�Z�<�4M=g�=���<��=�?`=t7
��ᾼ;���^���ㄼiOU�΁�3"?=�m����!�ru��܆�<9!�<��ʼ&OQ��1U=ʻ��"<$f$�6��<�ޯ�*w�#������%=��sἥ=C�;,����E�;-@��վ`=�y���=�n��)"I=<��Q�{<<i�<U:���7=ӥ<55�a*@��"���H��Z���p܍=�)�[/e��޺�dс<� �<��7�.�= ~b�f ���B�"腼S/=쯼"ޏ���P��Kr=`R<:4F=���<�P1������ � -�:q�k=8��;�;�< 5��=��;�=���f)=��5=I;�<RbX=gR�<���%��� ����1�c�q�-X�<����K<*����.3=���Bh\���~���˼8�6="�j=H�t<w�s=�t��/'Y��Q���g�<�x��m&?=�nF��P5�W�Z=�|V=�N���}���}���<h=������%��=�<��K����;������<=p�;b�/=l7�;���=�%^�X���7���-=�7�<R�>=�ɼ@�(<	�&�{�1����<�b2=B2�<������,=R��<N֎<�19=����ͥ�<_��jn�mP=�b�<� =4r����!=�n�<��r�윖�a����#��7=�zQ<!	�;��[�C[��+}�[��̖; ��|��WL=�(�<��<N�����:�Ʀ<Ͻ@��9=�M��<�ܜ�O�:=t�!�����v�[�Nݖ�w����);�F�ȫ����)Q�o�O<.�e=1�<.�����l<� =1N=Lnz<*�sn�<J���$W��p�j=;����U�^\������5�	����YR�\H��ؠ=jK;����
�J[-��U<�[{=��0=�O����6L=h��;��=�O��6�<K4I=�Kr=�aF=h=����1:W�E=��s=�V	���==ӺS<f"�;�:X<T�~���5�<3�D;H~����9�m'��;����o�<	����=�f�:����6<�s���=G4�<�1=�R%�0���Z=NԼ<�[��������Y=j���^	A�.T�1U�x�8��51�h�Ӽ/O�<:IE�����T� ;��h=�_�=�=d�ż2�
��?��0=G9�A�=�у�0r7�뀇��:?=z"I����:*lZ=@V<��
=�%�Wk�<��F=�&[;]�0=rO�QM<�7���P���n�V��;�Ǽ z"���A�t����%�򅅻�����.=b��<�a�<b8���L=I��<��$<�F;�1?�oE��;T�<'�ϼ�.=�Ў�x㟼�S�شd<�e=h\��k˼��(=��&=���'fy=q����TP=	 ;�/=y��F;b�	=��<�7%<�\W<�`r�\��<J͓<0<MQ�<�*#=��9��Z�b�<T2n�V�I=�3�ڜ=2�A=$�м��)</:�$�C=�)m=ۊe<7�伝Ў9�z`;����� =�v�<�Pu�ތ=E���d=/Z�<�W(��)���N<�49=�!5=Ŀ�����A�=�j<_^�<@V�<�91=s
�;%�����<�e�<W;=Юϼ���N�=�O4����\������Ŏ����;��=-;�~�\�|��I�X<�<�ta�<?Y=��|=�5�<�������RG�l鷻�X�o�M=����W��*��=<���e� <M��;���F.��	;���S�A�������<��<�Z�<ރL=o����3=n���;��
=��X=/v�k�=�����:-=b=�;)=��޻'oF�^>�<u��K��;<{��>ӕ�^A<v~��F@�<��K�:TM���<�9�=�캼
�<E8��C�<la<޴7<-����n��.�:m��<p�=�Y���f=�}<��<K=Q$}<Jż�`�;�3=�P���^<6�<���v=h\;ѥ�< �0n =HL����N�'�¼&$>=�mY��q�=���=�<:�5=(�<ʰ��*={#M�Q��h�<��?�i�'=(O"�D8���W"�$�����3�<�Q�<����5���%<�X�����<yR=f!�{\+���{=��Ƽ�Q��ID����	< �\�Լ<�=��<��y���%� �$��N;F��;)쀽�s�<%l=�R�<�J�;^�2<4r.<����,��EX����<@U��@��<=}�<���H�;k9�<�J;<X����]�<�2B=�2�<��.=������;P�8�S<�1���/:W�8���6�;������1\��`�'�q-F9��;=�v�=y��h\8=EH�_Rh����<��H�t���'=^��:�ۄ�캫�KI=�з��w=}���7��;���<���<@�}=�d<��1;'����<�AN<�o]:O"=�3�:����=dO$�l"I��̼�PL�f�g��j�����;<H��r�I�=.=J�=h�0�3<4�T=�,P���亦�<���X��9"�m;��~<�[D�q�<zm,��=��;ǸF;2B0=���v��˯��e�x�8�>�漎8�<�[�;�� ��f�;<�����z=���<���[v+������9�����\����+='�Լo#��������~fQ=�L�$�=E�]=�:�;�D�P�Q�Uf�=e�żi�;�=9Y<�;���;��<��Y=�:��7'<ʅ(�q���,=Y��gJ=ʇ�=��a�7�ü�7=�샼W-W<�q3���C��v4=���<�f���^3=$X��+���
�v=�z����;�O����n�x�/�2���5�R�������p��z�� G�<X=0�1�j��v��)= e=���<1�ֺ�<�%�<󒮻�6=�4<��1��;�>p=��<WT���=U���H��{�J���.���DW�@#<<�k=G�H�vP<���=��;�t?=��Y�ٽ;��	��t=o'�:�$=Q�e��:���<*=𜠼�~g��M��Y0�0��<ˠN�-�����cn5�@f���l�<}Dg=@��;�j�u�b���D<�b=j�<��,�=��<�t�` �<��;Z�7��f
<d�����1;x�&��@t�2�"<�o=O��=��{��c<�[=ܐ������h�<
��'=_*��"���,���z	=
�<�Zj���\=)��<8���<���Ψ}=	?5��!=QKl=�r��$=�=�4=�l��!�J�m:C�=�mҼ�c�*����'����<�q7�"���SM��|J��z��;<P;)݄��p.<�b��L�<!D�<d�*=-�%���j��	=�<�`�M���kS0�*�3��m8��U=�-�<��j=�*��ӄ<-�_=>O(�����@�켃s�<ќ�� ����h�;�1�<�:���a��1=�(�<	��;0�4�;[�<�
K�6k�< �q�I���oc�;�(��<]�Q=Pm/�.GK=O�u��O=�\ݼ��+����<�o �Y���cz����!��!<4�D�3�S���<Y�8�=��W��t�K=�	�<��0�@������x#=��0�a�=�%�@�[W��Լ?<�V9=�Xm��楼�<�4<)��E=Ix<�����~q<���;d:u�4c�<Z�:(�N=�������mK��jJ�{8?�H�a��^����<��	=��Q<D85=B��;2�6;g]&��d=��J=/��<b�R=M�<I��<��)yw��9���M�IX=ۅ%��<N��=�~�;�3�H2�W��<��<��=�It��Q/�7 ����x��:�=$z��{��:� ?�[�:=��;H�N��&�<��<#�x=�28=�6���k1<e������<6P��+��<%�)ͼll6=���6P��B�<��¼W/;�}�;֚<�v�K�t�g�<��M�PzR��U=�[_<�Md<B��;�y���mJ�<�gk�BYD==�B��~��`=�� =���<�M�z��:a��<u�C�R\���&�S�<O�Y=��Z��B� ��������x#���;C�C=��>�P�ͼ8�E��o?��t�nLU=���������I=�d`=�F��+"[���<��:<o9}<ת+;���<:�:<�Ǟ��c��`��P��R��2'=4 �~_��[��<%�f=��-<���=B�N=�=�� �:�
�-g���髼��<wQ�<�~Q=W`�;+Ǽ92����<2I=��<@�:;2*n=���<�dg��e'=��=�+\<5 �VXf<�틽C�j�\�<��;�Zr<C��΋L=�Fe��~o�7=�O=u일���sP=�a8���H�G#�ov���F�����𺝱N<S�ܼ~^�<s�ּ�?`��b�<;�'�#���TL�U6�;gQ=˵=�����'<-�C;L��ܢ<�1�������3=�R7=U���K�<O 2=d\1<������9ě����<|Ƥ< Q��HS��޻va��8��8/;���`O��ꢻW��:ӿ;=��v�V�V=l�q��<S�<.w&=�_ȼ�6I={�<�W��T�=��=�Ԭ�X;<]�D�鸥=�X=i~�<��=�%=C�=�$g=VC�<�D���i=��;�)�v�#�kl�<o&B=��޼\�3���Ǽ���kN=un�-|g=��&=t�Y<�w�[����'=�]4��%�;���h�[=Cqc;hW=}�����z�J=�	�<?�"�nE�<�vJ=�	F=+_<&{)��)=8Ȭ�~�<�ߵ��>�6/�<�5=ƹO�S_ƻ�p=|���Г�BP���hx=m����C=
e���X���<l�<&
�;Ξ��x���J�;Ƃܼ�!=�0�<�'�=p�μ��<���<�=�ۼf]��p� �)��<9��\j<$2�<���|��<y��<Ƴ�<��~����<X�f����jC�;��`��r����=$�/"<~���:j�r(�<��j=���:{'6=���<�P�<͜=t�;��+���;,�4�\�"=<�'��j<5X��?63��E%=g�+��\<61a���2����۲��d��=�8�^���b'y<�wk�@��;C�1=kl��p�Ѽ�����任M�}Y��vf���?��^ͼ�7�<8t�!%=݀j;�T/���N��<2�۟�;*M�<���kY�<470�s�8=�"�ǃ��<�F<������\��1W�ۙ/=���<�,��@D��)~��<=�?鼷�P=�EO��db<(|;�e�;�I�;�!:=_Et=��=�{^<�Se��U-<G�(����E����μ3 ú?�j�}	m=�c��^=�W����X��-::�E7�x�<{&�&��<��<�#��<`O�;��7=�u.��M=��h=E=:�J<�m�53)=����Q�)�����;+I�X�/=F(=3l=is�<�R=��<)�d��r�h��?3�:�M�<%��<�;=��<�+$=e�/��%=��C;<( B=w!�|$o=�E=V����3��5�m݉<`�b�cD:Z =qê�od���`�x�2=J��Dư;`��<�4��o��D�^�ul��L����HjƼ�q��X=����<��m=1`�֨��x�B=]pѼ�h=�I�c��<.��^xR��c���j6=�2d<ERݼ�xQ����<��:=?�dO��W�<F��=u7 ���2�X=��/=rva<�qy��� �-�*��� ;���<'��<j��<��"=�X&�5cE=��y<��Q�՞K�E���L=�'/;Pն���=�Z����=���9*_�<DХ�7�$=���<}e�=%�<K�X�
�<�'<�m=wc�}��=ٝY=��s<)�[=���;:��-�<�@�=P؂=I�漉Z<M�C�@U�CJK��	�<�cC���l=p==�]ּ$�ټ=�L=�\{;��+=}e�<�T<���Ƴ�<Or���:=(�8��(��PV�'0�I{=au:����,=�ļ���;CbԼ���<T\�=�D5�@��<���<Y�C=Y����\6�7uW=Q�;��v�n�b���zF2=q��;?;�`�<��=��<!� �ru�;�a��m��X �=�����<�l=c�Y=@x��DRl<��;"++�� K<f��<��W���4�7��;�����G���<�5-���:�t=�Tٺw�5�L%��i�����S�n=\+P�fA�5��	r4�*�]�ݳ�e<
�e7���6i<y�N<Fwp=��6�^Fj�P2(��x=��!=����x_�<s=��&<�A�<.�=%�=`��@�7=H���0�<���裏<��,�!{=�(h�P�X<�$�<3x��X��F3=bc��+D;�B=%���N,�<aӇ<�)9=���ƻHS=��-��o,;U��<U�+��޼��=Ժa���<= �<�r5���弬K�U7=C�9��!<d���&;���?��QH�M=fj=�.=���N���{������7=O�=���:#�[�-�I�[�3=�!�<�����Y=�'(=A�<�Z>;��==�k=�b�8�M�����=�5�3��<��_�������;�E��t=�F�<'R="5�;:�#��iA=��_=�l��N�<@�<2�+=aܝ�<P_<M�\=T���x4:��v��=i=�V=�1�D��<S�F���=�U��#g��3�x��9�.�ߜ����g��sc<l}X�V&X�tx��8�<���<[�I�:k�<o��<!g�l��<�c�<�B��E��1=���[j<��߼�T=oA=EJC�$v��Em;z�"�L=��_=э�<0'����5�^T�;�t=��/=ڟ����<$�w�B�<����b;���<7���� =�2?=��<q����U=DS==�	���E�)%�<�=����;�
^���<��6���;V�:�W=ɣ/=�qq��1=����} +=��k<C����;��G�p���CA<�43����:cn�"=���v��<[ni<)#.=��D�9�z,m=2�ܧ.=�`=-��<:Em��`<�,X���s�ix�;�0-=t������y&=M�s=�@	�[�ػqi�<�ޢ<n�Z��~�<�1=�Wr<��;��:�n�<��Z=]����(���<�G�N3m<�X�;ۊ�<W4<�`d�"ż�"=�(���=�!#��P>�@�o<�㥼w~��{_<87=𔅽�ٻ�Y)X=!.V<�	���r��»�<_̼2�=gH=���<�K�d"�<�k`=��<��؉�͊;�SL=o�<���2=�
�l�޻�ԃ�Rg���CH=M��<3�=�L�'�f�r]�:
�j=]F�<eG�:3v+<��>�] w�#�<$.!�0����l=�\<�'��Ȗ<`�m=��=ڝ�E�="�<�'=�=D\X��$~;��;�==�d;5��S�<>7D�z0P�lw=�6V;-���Mo���y)�_��K_���V�GI�<��A���3�R�j D�@a�;CJ���+���;l�g�E��;��b�<��̻�S����<A��:��ͼ6�<aw=N)=@浼:� 8�Z;G~���qV=�}P�]�{<�(=�^;��X���;tCU=p��<�Ń:J���<��!�e	�� � =2�L=��<7��;�R㼜Ŏ�OU��U�<B�����t�w��X�;:1=�;�?=�Φ�"<�<8%�>ӥ��Y������I<��z�׻�缘 :=I�(=�B=|sػ�e�<��F<g��=�Ҥ�t��<��<��J=��_���ü�+t=+{\�L_^�}z��n�� a�[v�=����7���1=<={�D���h:��<�����n�9�d����<��f��e�;��'��A=�@��\K��U�<�����5�<G"a=��\��\>=��M��-�<;�nw�KiA=��a;^���><�;��<u��<4�j=ʕO=�fh<&�6���C����<��5j;��a����@��<6����F><��<���<�
�<�F�<�̐�v�<N³���!��'=U�<�~6�w��<��M��ؽ<]>:=��>��4����9E��;�C�<9�d<�U=��3�M�#�u�d<�N2<�z�<�=�oyi�Iz=�,=I�(=���-�^�r�A�\��<<�=�gT=�a»S?��Ʒ<@c6��!<�9�<RI�<�
C�;�;��`�_�U��R�;'?I�Q���Qh�����%���<[f����I=�@?<i��b=%/�:��#=6
�<l�U�J=f5�<��;��<g���2�p��<^�����Y=�;1������PG=xU���[=T6U<�&l=���N=U�@=n�Ӽ7��Lf=�Y���=��J=�(�<��;�3�<��;��X=�<`=&Nh:��V���l�;�#=��l��p=�cc�zap��v�������7#�t"L= =�.��"=54�+5=�S�G=x�<��.=,g*��[3�π<��J;J�޼2�,=9^��2��ܫQ�/�<ǁ�l  ��_���;]��<�T�`��<�<^�g="�ȼ���<iF�<v�,���]����<���;ɱ������<��;XI����<�μ�1=|����5�-@K<����4ѻ�Ѽ�
�<�O/��t|=��<�D����<�!�;��e=�3:=�ai�[Rm�����_��3�:f�e=
�9=\?�/�V:�¼�?=P�Z�'֕��%���2�J=� <�K�=|���?�<�ʜ���=$0;�^F�c6=�t*���g�ӽ��#��h�-��d���A=yV=}4�;�
8=�_��E6�K�����~dM=�����!��$1����q<�2j��Ռ;/G<�Z4=�	�O��xK<�ʼ%��:��<I;��8�<N=�tl���4�tU���I=ԕ��#�<�j��Ƭ*<�>��C�<�
R=u���
�����5=�u<��O��E�Z:8���<=�cڼpI�<R:�;RE�Q\��	A<���1�<�9<o�s<0fm=��0=1������J�'�F���=��>��*
=���K�=��~�F:E<�̌<�4���<�H�4<0*.<L�9����<�;�R�����@V�<¡����"= �=Xg�=� 
�c��<X)=�uF��X�;�~��z�!��m�<cr4�Uo-;{輦��;�'$������<���<ݍ�<��Լ��8j����G�=,���F�~琼��c=U�<�H��NZ=�VF=������<�]G=���<�+�<#���~f=��&=����X��Y}��Pn�<�/<q�7=��4=Snh=�~=6	�<�3�<��<2B�7il�����;���_�j=�-S=�m����-<���<���<2`��f�t�M�[�o<e<����ԁ��� ���A�������];����)��.��;l�5<5b<�&�<�H��o�W<�+�<�&��$�������Z��7V��t�r�'���<5e��ļ�Q.=#;��H�1}J<t�~<�Y=��<�׃�xV*��Z�<�>r=�����-�����X�b��w�< �=9@!=H�N=vP;_���[<q��&�y=xsV�u<'��#r�ǽ�<�G;=uQ=��<���D�a�$Ff�5���1!B=Ps�;�Z=�t=���<�Q���T�Y����<���<�\�<dv=�z2���1�N���v������;CN��ݺ�g�įn=W3�;���\=;%=	d��U#<��d��ƼDl��׼�<<=����WN=#e �̋!=WQJ�
��<1>�<��k=�EB<�&F�5�(=JEI�E}��T;<KV*�-a�H]��>�<--D�Ф��լ <�bM�t=��3=^X���<��==T���T<dԾ��~��t�_=*�; �� �s�I=��)=/�����M<��@���S=�*�x�=�r��X�X��k<�FW���M�
Vͺ��n<_�.���t��>Y�l3���$=+ g�):��O�<���<
�P�<%�&=���<�͜<�Nd�G]X<���xuH���X=&t<�G��iib=V�=�x�<2��C5=� �J�Ӽ͑G=c��;Vlu<��P9�qb<iV=���g��<�i=<�,<=ȅ����<~��<�1���<��a��e�8i�O��mϼ{��<=t�<�;�M��v0�օI<k1�����n�����<;���,�~���c<'��<�|�;�iۼ��ü&]ļ�iʼ����6�0�Y��<�	<I��<��@= g�<�4#��ei��A=����F��<��Ｑ !�oN�������I<�zH=}���I�ܼ���<Dj:�����A�[�Q=��Yx=�=?�C��8�h�)�|����I��=5|=$ �N����J=�����z�<WD_�Z���<�ϴ��7[���<�-�=�'=�]!=[唼�%B�)�'=���<�1�<��
�Ҵ��v����;=�1����=,�R�&V�<zF�����8�vѼ�q\��»< �R�;ʷ=��Q�m�Լ�ll<��:�<�Cw?�9������}4=@�(=�;�6K=P�d=i��T�b=���<�ռ�h<�6 <7�<B5;�]�c�N�`����7��'=h���d��쯼3կ��{��Ӽ�qt�V� ��_�<N@�i��<\�<p��i$�4-缝�0�&)#�~K:=�����E==��<?�H�Or=���=P�^=]s[���=�kU=-H���S@���6;��!�rU����<W�T=RB�<h�+�r �<��=�5<�E=�g�� <7b=2}4=?2(=>!M<'��=�&$�k:9�E;�Q�;�"廂OA���~<d�6��=snR=N"[<�Z�<�G=|;�4���L=ċ����<o2a�!G�<'�<��8�����ˊ<�`<ac��Z+=^� �"��<u=��<�\B:�D˻�r�<Gke�G/��'�)={���
iQ�����ہ=H�;'��0r��&<�~&�[#o=M:N�QM���;�k���$=֘�<J�g=�6=�Kv�e,��)0��*g��#=oGl=!�]�nU�<�A���/=�I���� �h�;F�f'��U����<(3�<������;%�<L<`�ү =�����ۋ<��<R�T�`�ռ~�;��2���<��к�چ������;"N=�]<�n�<�Є����D�9�,<�ռ:�<,�<-����=���;:�=��<Z̥�fP=�h��$l�k=����ï�>j=R�ټ�ü�K���%�K@�;j8�h/q=/%��е��E~��X��7&"���B�����S�M�V�^�
=UM^�ķ���<'�
��B.�;�Ҽ�9�<j�<R�ܦ!=!"��?
��� ���6��H�n�<�x����<���R�w;���<��u=���;�^�<�3J=q%<:r���	��*<��doؼ��d����<�E =�]���"@�����u?���8;9 !=9�$=+v�/�<��>=քv�t=
�S=�D;<Z�u�su�<�zD=��6=��<N[�ua���<�f=L�.�$"N���:�(`�X&
<�k˼L�x=KB���]F�(N6��&�:�)���NQ=J�e=y�?=hz]=qgC=�I�����<���:tw�i8s<��b<������<[Y.=���<ٽ�=o�;^ռ6�9�,#�<�Ƽ��=%�=n	L=���<��=A"�AhI; �7-e�;�;��[<�=�PQ���+=����"��nx�<qW��T��([=a}�C��=��i<l��<�w
<=�<Lڎ��ߚ��HM<j��C+=o=�R��=�$�/�=6�)��̰���S�a�=[�R9�:�<f\U���[=w�a=ߊ���'�<���;��b/� Q�<ݴ�<����^�;;?�<}$����<�<+�G�!�<��<�L�Y`I=̌n�#A���^=���CҊ<-�'=�iK=�}����4�c뻁2�<�/���~�6v�;��;sͼ���<�@=�	@��E0�J�G����;��S�)�=shӺ�|�<
=u腼�����)Q��N���=�W[=� /=]�?����*��,=jS=���:6}o�CE�;�C=�޻�6�<�|]�#����;k-���w<Ef��}�<An��:q=zz=�c�<�]<�D=�QE=�
R=���<�6F=p�J<)#-�P�!��gh���=n�pf�����]����<
�P=r<K^=&B;0��<���;��={�=��T:)KM<�j�<Q�U��=��t�|�����Aѻ.��<O(��л-E=�-X=�8��UB<wO3=��*=��<������<�R	�0�5=$��;�v���&=&��b�y���ܼ�_=H�#�[�<�(�m�)�N;k�s=��<:�H�;��<��x����iJ�j��<�S=���<��c�=}m�<lg�?қ<�NV���;���<�@=2��<�v�<�v�<��t�/{�;�4=����K<X�*�ē=��������zb�<�2d<xl<���C��@�7�8���A��QV<e=��1=��i�z5l�� =�K=<�ƶ��@�<(P<=g�=KD[�x�Y=t�[�<���<VW==���/�9�H.��,��';�Lj=r=�0�;hoj=N��<Ar�;!�<�����B<-6]��=�2="X�<�VU��]?���;�bi�{ -�'=��/<��<�?=��=Ҫ,=��<��=��������s�D�"=#t� {��!H��1��[�	<6��<������m5��J;��/g��o<��.=��-�?:)=ѭ)��S=�=B�S;ӿ��o��3�ݼL���l�=Q�T��bJ�,�<0�e<�Dk�&P=�������0M=G�h<iD���?���]=�B��<^0�<�D��jI���1=����rb��G�<�r�!�/=�Wl�h�+�M^���X��!��;&	;S,I�)�<ld�=�=�,<�mV=�AO=�]�_G=�,����<�6T=yl�����T�?�%_�:�ܼ!_�����\�
=��7=��7�W�˼�^��N���V�S��N��<�-��;֐=�I��#?=� =��=�`�jI�<;VƼr)>=|x@�i��<����t�U�����ܼ�
%="�4��=U��<���<�N�D--=�� =��.<�YM� y3�*=��
=�sj�e"=�	�݊���<�/=/-V=�~b=HS;=��7<��Ἵ��<s�,�?<Y�.=�FI=\�=|�=F�<aQ�\�}=9!��/h<�P.=D:[=?�N=��<���<�=G绎����6� �;OL��Z��m����<��L�3�;��JF+���X��gZ�w�ޱ4;D��iϧ���=��o�<c�i�}ٚ<��N<�8ռh�{��T�<,�<};=\Ǽ�μ�U0���ż�nU��G=2.��t�<H��l�=6_�c(;�����<���:���Aл�l�;%?�w@�0�l�
��/iP;E�B�������
EX<7�^=���<Ą,����<!P�;��(<���<9uH��f���햦<?7:������:�=�#�=��Ի��4��J=mh��B��=��s<X�<b��L�<�;�9���
=�Ϻ�n=;�=}7:�M�< �=�[�����e*�խ�Z�k�C8�=�R1��Ӽ��`<q���2�<���<��M=9Z<��)=�Jټs?�<�x[�˭X�=��C�<�P�<�p=�,��%,�<�D�#����bʼ5FE=L@�=�� �uP�<�&%�rz���[�:e��i�==S?=��v<a�!�clؼk$Z�N��=3 �����<������d=�^���=�;;�
������:�<ic�$�3���<��:=��'=��ؼ�D�<���<����^׻��X=������&;�.�=Ǽ�Kl1�Z�;��y<��ۼ8��<e�)=�\�<
'�<��<�2��H��:d�;�LI�d0=�s	�#��<�� �|�-=�pӻ�W=�� �VCT=}�:Jc_��1�<�/d���L����<��
�%zI<�Me<�C=Og��fʼh��<4<;ba��?�<<��v�]K���c<��2��
#�q'K�v�0�pv�<�Z!�l��<[�e��?^���h��|&�PA���]=��<w��;5 =ZNw<PEP;�Yp�F����;�0�<{��n��<5�M���i�����HE�<":!=��#=�<�{v��~J=��ļ��1:>�'`=1���`<=��o<DC<|�<�#���*ڼ�[�;��i��ed�0���wc���k=y1�Tkp��C=eF{<���F��%=.B�c&�G8=� ��~=���;��&�N=�Z��J��<<�=���^�V�)�<ۍ���E�S�G<��<#p�;�2���;O�<l��(��<�F&�,c�<�!��LM��a��,=I����&=��:�/����j=H~3=R�<��$=�=L�l=�r���N=�:=A.�;�[:=�� =^< =��:��>C=�,�� �y��Î<S�<e<=�;=c��tqG���d�mp>=��P<'@ݼVa{=��e����<��<8Y/��Q��>G�;8���y)��E�Y��0 =�-
�ſ<�B5=�>����8=v����Q=��"��W��dԼjA�<+�6=�0e�<�t���H=u���02�+�������vdP�A�=�Kļ4\~<�E=(��<�o=�g#��,S��G,<33�
�^=FqS=ԑ$�o�<�y�<6�]=b�e=��;=�����$�<$�7���5�]ܶ���/�U�j<t�O=a� �z�A�]*=��P=���;7=)O@�~} �*�4���)�G�<�����s߻;t��);�P�<f.�9գ;Xs���H�#9��u$��m�5=�=S�<��W=�wܼ�kk< 6��.�ػ"P��k�<x�*�A[ۼ;�z�G���D��̂<--���8=�#�;�#x�Y1N�k �;?�=oļb��l!=n!;� =��� �Z���U=�#���7�<p�'=i<9�C�`[�=S�6�ǋk�F�$����h[�<ߏ�<�6��k2=I;���>< =3E�<r�<!=�;���<Ǌ9��q��ًZ=r�S�j0��g���	'���=3�|y�<c=2�Y;���<d� +=ާ`��1����c=ñS=ㆼ�)¼�*����5=�����+I��L=���<A�=�X�ǡ�<�T���OT=J j<�Fc��=�/�<����=�酼��K�����v���ɘ��0�<�iûjĞ��*�<�d5��oI<W�@�K k=_JR�6nc;�9F<�P����k�̈m=(4�<-а<a<r�x黑�)=�T�=��j<�RO�3D���<��T�|�f��=L��;:���y+��V<��u;J��<�|��t�<�,P<�H@�����H ���B=o�;]蓽�����R���1��Zn=�d`���μG�"=йD�x�<N��,	v=��<V�;f[=̝��-����<��=�)��=��1a�=��&�bȂ<8�{<�伙=H����<���;���,��%�=�st=fW	���E���8��B=F���[��z�<��<���MI��'̼��-=q�ۻ��D=�;��{d�Dќ�:����I=?%Իy�;݌�:�1:�5�.=h��:�޻V=;�I=� O�եp��
�/S��K��b��
��.���_=x���Î��[5=
��A�;���<ä���K�<A�e�ΰ/��<8�<$l����e�̼��<1ch=��_=&��<[Y�<��<#��P=�@=&G�Y�_=�]�-G;or�:HΎ=��<����3:$��91=��9=�~�<R�t=�+y<�^�*���#?Z���T���`=�5<�r'=0lk����@cǼ�5= ϴ�+Z`<���<Y�ݼHB=�=�<|,����*=�	F<v>����<VU	=�(g���ؼ�$��^q<uD=MA���?�-S�̩��Å<�
C���=<����Y#=���<�E3�=�μJ/=�ػ�@j���:�Aa;&�0�o�<tդ���=�Q<�O%=��*��X,���-�k�:;�����
_=��9;�}=
>+�-B�<@a,=ń<=?�;�2=uj\<�o��������<j��<�Y�/��p�<y8<7]�<�#x����<>�=�{9�M���$<��<6B����<����� �Q�C=ǹ!��EM=ZN(�*�>=��<Z4���P<*F!=�r#<���]=�K�;�"�:%4!<�[=���-"0=��9�$@��D�@2�%V��s�=�8�;�%�
3(���o;z�<w�<ƍ�J[=���7�V��&B=������,��8.�t4�<.ܟ�|��?q<�Ｚ胼7���}İ�����
Y��ˁ=؇�_^��A�Ϳ���9>���<We<�(����;�H]<� �̱��	D���,�o>3=�c�<<��H^=cW��FL=Zx#<�]��"L=< �3�<�����Z=�D�۪ͼ��H��%�=6@�6�=�c<��;w�V=����bb��v�<���g��;��м�V���j&�f��}�;9����ɼ)�*�+�
��إ�G�6��"���I=~�����;�W@=he�<��E%�;�U�S6*�kv.=�v'���;�c=���F�5���%�4��<9�;�n�H��9��|�
�;�a��p+=�P=tqK��߼�*=́���=j�eV=8C�<t(v�e7=
�=F�A@���M�٧L�!��Q�< Y�e�
�jq,=���"-e=d��Q��;��=v@�=����/�<B	�T�W�955�iS=+ON�ʧY�E��f�O���|m8<w;��W�6�����]=��%�Z��<
���T=&�P<�"=ҩ6=Ǻ���Z=�-=��5<XO�<ׅ���.��&�<��<�8�s��A\=�zP=��O=r��|��<[P��=�yk���;[~[���/����<^�X<���<]W2�3�m=��F�Ǟ=��H����'a�;L@�[^W=�������;=�;
H0=-�	<(�:��5ҼLD�:7��ԁ1�º?�D����4=��)=][�<!�<��ɼReW���;'��8��E<g�i��o=�¼��<�V�����;�<׿V��4�MIE�	�������ԕ��#�1��J�+��<�a��hx<�ݹ�)�<Xn���RۼV�<�+>�:��&�<ˊb����<r��<�Mb�u��;�[�>s=.�,�|RV='ʴ;�ò��M<P���(��9���?�<$�лk~��MY�<�Z<ޠ1�B���m�<q�G��o�k�:=K*,���<��Y�cZ�<ꕼ�oټpt���6X���t��л���H�<��=�� ���	�š��xr�U6'�p
�<I��!+=)d=A
=�a=%�f�kRa����W]=ޜO=጖<�o�6"a=N�s�gH�:H�)����~���=�R�����q=��	��AY�9ӗ<+�=��T�'ϼ ��q�9<VH�<��L�7�C<��"<�9J����<���=�=W6={��<́��>���+��nF=��3=~~�;��1�#ۊ�*�O�� ��r9�}�3�גB���^�2��K=�-��֭+�g�@=~��j�=x��Il,��/=�k=�E�=b[*<h�<��5�3=ɓW�G�3=;��L�J�������sQv�x�=]=0���Y)=5�<em��W�=�F�7u�A<�;n=`f<�Xz�e	�<�����d;=�޸�	����,��K|�<Ơ<�2P=P_�<k��<����I=�m�=v<�]=��{��c=�x����;b��:q�����;�ׇ;�����h;�4P���߼�4�<��=�C�^Y�#Z����<�L����Z� F=��<����F�|�N=��,�ĕ���A<�H=e��?}N=uLh��`�;Kj��A�9��A}��WA=a	仛�>=���<����@+��MؼOC4=��;����A���<'4���;���Ys��֡;���<T�T�:7&<R��9 �;�����ܣ<��A=0� ���ռ��� �<�H���cg=�9���l=�+7=wl=S��=X����=�y���_<�����/ּ�4���A=D᜺r�๜
�[A?��d��ϧ����<R �<�[!=\�c�&�I<�zS�W�Ź����\q�ɘ%;$�E=���Ap.��
�m��<��#�	/E<�K���۹��4<��ػ�v�<i��=�6��<b<+�y�&=�h$��߹����@UD;���<�$�<�
���I�<P�F=���=��=���<\�i�;Ժ�;�c<��U=ե���8μ��a=���9�gi=6!2�,�$��Ap;tw�)V�k�˻�T<x��;�ZA����<iX�s=X+�O}=)�@�0�H
��C���S<o���Q<�Gh��gq��*�<�;���w<��ܻ�����*�:f�=�����R�����E�ü���<F7�o%���K<�ͼ�q=8,=@2_���=D�	<-삻q�D��rZ<(=��ȼ���<�m={����<�F�<�L��lE��.���=�3=��=�;��삽
�Z=e�-=� =�=`�K�j��C"���(=ʰ���7=�#��ﻰ���,<�,=���<�һ��<=MT=(1�;f`�;k�[<oJڼ�a�o
<e�8�<�2 =��M=�9�<6٨;�T^��h��?�w�{}��ŀ=� ,�L�=%�*=B�<��*=�"��"�<��:=������=%W�;C$8�
2�"a������+8<�Y˻0�<\�=���<��<��=:JP���,=w��<�tI�Z�v;ˊ]=��c�m;= G��b�2�pY�<�dO=���>*Y<���;eK=^�"����xD�<+;��4��3��@<����ڋ�;���!´<4��;��W=�S=6j=�
P��1(=��=�~Q=��<�I���G�*E�<�$���(��=��<Onc:�3,�����R*��+
��*r��p�'=�0[=d���V=��<ɹ��<��<ލ�<�I	������<g�q=Z���?��<��<�sd<�р<f�D�]�=���$�?=ba@=��Ҽ��dhH�q@�9�Q��[*=�%<J��<=,=KDd��~q<6�l����<��C=��<|���m=J���:=ֽ��d��<��<i8�C������;�X�PB =~�(���	�]Fq�:<�<Ƅ5=L�{s���~��O��x^�<��D<c�Q���h�<h{�c�j��p<R�L<:=��8d<��̼2�<� �h���q�<󑉼;��LO�<>�=�=�E=��4�C�˼�ݼ��<)���^�&!�:�h�<�76�9�+=�G#==(���+=gK��
;1t�f��֮[<�G��ȼC�d��˄����;�Pc�Oc�!�;=�==��ּl!�;1h �����,�<�5=�u#�|�ۻKt���Z<R�@�>=�7C=Ƽ�^�)<�_Y���<��:l|@���»�޾�`xx�^����2n=g�)=�R�a�A�z�=(<,�6�2�<�$X��nK��<DE�<r`l��P@<�"=��L�Ӹ@=�n�:Y=r�,=0Qi=�t�5#g���<9C_=�����g=���mG����<L����8�ݢ9=�%�6���e���ڼ��'=�$�g�=�<.Q��
y=�m�<gF�X*=�;M�/fM<�j*�0$��,�����{X=S_ܼmr.=�2�<x����ż�j@=l���U�;oܫ<���<�Y=���k��<��<�uY<��g��s<d�<��8�ʼ�\�6���<_Ѽ��a=��`<��_�N/%=o��;tϼ��t{�<Lc�l	<�M���"4=�<�R
�i�1��2w<�Ɋ=˺�Ps$�3�V=�^K;C*0�$��v�K�x�;*�<��,=-w =Vs<廼����Uw<�S�Y���]�]`����<ʳ�<��.+����N�"��s����P=��I�+��<�-���=��:0=��1���{<�ٻ�!�<S ��r� ;�=GE=�Q�;J�>=�_k�YM?���ʼR��V�)�_=��$��u=���;@�<�7��Z ��C_<��¼�PG='��<��v=[,��	�>�<_}p<a�6��?ͼZzR=�vq<]�<�(+= Zg�4]�;�J�<U}����@��mk<��ݼJII����<��}x��i�#o|;+�x:��Z=aQ=�B����+�=��;�֨�)����\=
���/��Z��nɼFP���q��M��v;nq.���|=�7�LV<<��؋<��u;Z�(0Y=��޼j�'='H=F���bȺ3�-=�͖��n+�8<==T	��kN$=j�2�X��SM��e�<t�a=�)z;��@�&�r��
	��ox��_���XV<����E<��<+a��]#<��n�/r=����Y=��V���׼��.�&.<�i�[���<T�6<�Լ�;�Y<�	=�p����<�*}=��<��������>7=�==�ZR��"=��=�_ؼ�N =��⻅F7���=���a��V#$��~�=sZ9�Vpr����<��&��� �'F� (k=p����,<���<�ae��y����K�C�<~��;��\=�b�<:���@�<O�E=y�r=7 E�qc4=��D=�O��L�:�
[=B��5߻����.�/.�<�p>�hHR=z����=J�<8������_�;p������c"��^_����:ncq�����W�	���"=��=/J���׼WZ�*���E?=%S��w���d=����R���d�]wn=.F���>=��Y=by�6�?=��<?�<�c1=�O��`��k6=_f��[�Y��O�<?O6;y5���?<��<�i)�
���<�y<<��<{�!� o#��N��<h�O�E�<�
����4={�_���F=�w�9�t��Ft�j].=��h���< ��<�`=�~Լ����*=i�����k)=�ۉ<�Z��=���<���y�G�;X���,�:�<zK�:ʔD��'��j<�^�<��\=�^���0=��=S�����A=�-	�8t�<r��<w��<d@/�\�����<�]�@M]<G���	$=~����<ub=<w;��Q�=l{�H�l=_3=�qD<Yi>��U=��P<�n������"�{=��^�4��<u�=��)�^4L=?�-=�hW=��g=�4�͉_��-�м��r=��<�c�v%7=�\�������ڻK =O0����6��b���T=Vd=��7�da=L4f��&�<��]��O����4�<�#R=�iw��D���Ѽ%�������D_� �=��?�C�l=�!<�zؼ5�<�?;����;Q79=�/d<�?;K�c�6�S�0��<�Gi�}�~=<��<�q�<zHW<�X ;�U���=��==R=Ink��<=���L�q�0{��4J=z��V�=���<�UT=f�M=/bt<�,�<o����r���=R��	�Y�x�=h鼖GJ=��W�x,弨"����<���<�;���qI<��<!f�|�)=��<��f=��$�$=CI<4��Kfe<��7���ռ��=?��R��<!m�=��p�b=�f伿B�=�k���Ӽ��@���O={�$=ϒ;IT�<�"�<=�3=�=�r3�rjP��������<��x���м�nv�MQ,�m2P=�\�<k��mߕ�'m�<��;�/���Ӈ��Z=(xQ��%`��E�<8f���P=���<؋<�HL=@_	�n�d<�a��=s�����:���;�`=ӳ�=�g��C<x�h��_��(s=�@���ݱ<�52�{�K;����NED=��Y=Q�<=Wb=��3�lNq����9YT�OYv=qW=eD��Ʊ�r&|<Կ�'Wy<����0�mDs���`�{=L=������:㶼��-���G�mk�D���X
<���;�:�<G�;�F����BI=�=�x:<,�>=8=%�����;bY�����0r�<�b���:��S�ۥ=��Q<t`�C��:T���q�<H�={D��\I�B Ѽ�ow�i��9=Bo=!]��UQC�]�:=[@=���KH="	�;���<�ն���lc+<~Z(;���<��T���'�a���#S��U<v�3=����<1�=,�=���K���k�94=?u��o�6��;�j=�%�n<��&��@#=��V=��=!$:�څ�}�[=v� ���Y�L[׼��	=����%�1��<��[=!�&=�G�<��=m)��N��r˼�1���
;�M-=:W��U=C����oF�F��<ӊ
=Sؼ�_=y<�VA�{�����<��3�w:�;J��<I	�;N�ܻ@s=�Q��<���-0�D2�ч;�;:���%I=��<B(;�P$����a<_��:�}�p�=~�=�ϼ,�����3}&=*#8�jVp=!^�<!��"�=�D������o=90=�_�:(n<=��ؼ�P"=4�	��R�$����l��X���}=ă�ʍ�
C<��u"�QgW=rq���b<Ja=��=CQ�/�+=tn�<-��<�Z���d;��W��Qa��R=�F�`�{�Q�)��G�<�߃;�u��E==�8Ӽ�TH��s;�*�<yt=�$���C=��i=�f����:�9�Il,�z��<�u�;�X{�۫�;�)�9�52=�U�<�ž<�	�<Y�(=+�>=㻑�O��:�C���}<�\�<����X�5��k�<�����Sq��T�<[��<:i޼�#�;��p�&<-�M����=�<kP���f=�w�<�;=��A=H/<�S>�\�#<;��<O�y=��<ϼp`5���<�ѕ�n�3=+���ǡo=GW�ϣ��M�=�-=i�<ox�<�_��9-�<,7���=��ܼ��x<~��:wv7<�z�Ϩ,;U��<���<<	�<�K)�ЯA�q뗼�-����"���t<gE�<��=ہe�9�=[貺�|𼘐D=�\�A��<b�==� �ɞ����'=vb�R<�'=]�M^�<i�2�x}<�n���a��L����(=]W�Ӂ㼺z׺�jk=R/�=�㼑31��z=t
�<��%��o=����9=���4�=ּ;����}�9��b =�3=���<�u¼=hb��3=I!�;�P��,Y
���;��H�j\=+�=_Q�=/��<���8=�M{<�Y0�)�A=ħ<��c��5=������]|�@�<�@=��`=g/�J,=��:|zk=�����亝:~<(p=�¼���=�$=1WQ=1�������u^b<�1W�6�<l�;=��S<��X=�{�<��gོ�+v;II��2���<#=�B�=�*=<b����j�*����<1����6��L%<O:�@�=9뼨�O��?��3�A�	<"�Y^ջ���9�� ^R�N�˼,>�=<"	�i <��F=WI;=��<f=��6=<��f<��<�@*ȼ��=_�]��1��fƪ���="XR=�ט<Ƽ3<��l=�co=��¼��"�=gzc=3�=�@x�FL�Vv=�=�#��ʼl����󼓉Q=BႻ
�3�Jwռ;?.=��<n��<��u�L����vX=M��;u	)�r:=�2<no��Y�\�r�*�ybK�X�;^�μ�=-�=$2�=m�<�$�<5;=��}���<��=7s���;��O<κC=�_#����;bJZ�58J�`=-�꫃:���;u�X� =�==�$H��~<���;� 5�4���H�,={}���[�#M��WN=S��<�f�E��U�eXB={�Ϻ �<=$<�� ���=��);�.r�獁:��=*�R��,�<j�=e�w�e`m=8�<u!
�!̓=�U�1	T��w;�s��<C 9��ݰ���C��?=�t=e2=,�l�Y�D=�� �;=2�$=���2�=��=`�׼h�Ի����Q5�O�B=H/�V�=�`�Wz%�5 �0jf������L�L���X<��=̙=h0���;m��6f)�������a��<����=`���:�Y�@/�=Wh�<��<Ń��c�<VǸ�]�&=���Y-;w��cP=�\=%J�<#䔼��<	��;�R�<��;8I=)L��e����h<�ּI�ٻ��f<8��w��<��$=�<�`!Q��B�=@��jl�;$��^�A�;��\=B<����I=��r������j=	m���x=6�9��:A����O#��´:��=��<+�Q�]������r�:m��>�����4�ռ�_�<�]�<�h3��ļr^�T�;{K=�=�S=Ob"=U��<ۤH��:�:��T<J��=��+�<���Jw６<=2~m�x�?�bk��t�<M��<L�{=�=��6���5=���d=�O
� Q�<�t#=���� ���f��ƨ�0�]<1��������<������>��E=�K�;��+�<�H���<WB;��~<�R�"U$��&4<���<# �&F����^;�	==l<�{o=���v�{<Q�5=�����S�+F=�*>��*;:(�<��b�^��D<�=�@t��L?���ѻ�s�:̘�;]�<#L�;��	�2�&�?<=����3�����J1+==��:%�� �\��"�
="y��J=�2�<d�=;-�����<q�e=�|��A�;�����<�O#<��:ո'�6|�<O�=��)�e��Je��u?�
|=��<%_!=K�"�(�=�V�ϫ�<g:�W��<��Z���ϼ�=?�Foj����ѻ�b��/����S��D�<�
<8B=|�ȼ��<?�=2H=n�v<K6��P���<�3:�.y9=gj"�%FJ=զ�<�&c��*Z��?�=}�߼_b)��0<=Z�<�Y]��.<g�=^ǔ<��ą4=�̼��
����;UCR�w!P=�jB��kj��I�BJ <�'F��K=ه>�.+�<ǽ�<�+.�\�U=���;�;?Ti�v�޼>}l�U��<E^�i���Ϛ<�[�<�Z<�f�<\?��/�=�xZ���[<�S�8_�<�z�s �<����vD=�^F=�a <��7�ǋ�9f�&�f�<s,y<M�d�d�'�-Q��N=�����<=B�<8�y;\�=�8��ǻ$�<���-�<����T|=M<��M�zG<���<P�[=F����w��;7=��:А�K9�;A�"=P!���$�<��'=����3 �y�M�Ƽ�kͼ�(\=2#=�5����^=`.�<��E=�J=��Q��;
=�l���< a�t̻�G��*���c�(ـ�������W𼹵=<��X�	�=(=����]3�_b=���<uRH��$=��
=
�j������ۼb�9l�D;�� ���<�6K���t�����2=��]H��=A�Z�Z��;�m-�w8�< l<z���"d��6�<�#=T~	<����������S���=/���+M��%=��=R2���<=�]�s��=�	T=���;��;g._<��<6@=)6,=�h�;K<i���Q�<�"{�'�=w���;F�;�,��ah"��q4=�[2<v�9�jՊ; R��D��=�v�;շ꺔Gg=u$ ��5$=��h=�@л=vIZ��Y=ox=���E��:G����!z&�k�y<�z�<C�;?�-<{�4���P=��c=;G�<*�e<�����F�J��-@=�0%����0௼�76%�X�K҄<B����;�j=u4�������Nk'=���<�J��w=��<�I�;P�&��b.��F�:�>�=<d�4_ӼD���H�:N;[=��<��P=4ˈ<�&�<f=�M{���5�f@:�F�P�=Krw<���<2J�����<D���+ڼ)16��&<���C�=;{�<�Ŵ8�e<m��;w�7=��<q+=Fa~=�%�<N�˹�a�<Ҋ���U��Չ*=��7<�rR<6��<�l�C2]=�	�<�VH��I�;�=)�d�q"���绵�x��m���!D=V�V�K�#�'�LNA=�� j=�~6�$��<KW�<�d�<e�#=��=�I��� �5.n�y�=m�<T]_�;j�H�=�ن�R�=��=���5���w��kۼQ��F�=��͑r�20�a =C�N�
�=���8C�<�a���mY��s�Yh=�<}�=��=h6=^u&��ǆ���M���-��z�<��)=.���}|�9�,�<�J�<�(H�� ��|��<BU��]WE=�DJ�z����;Ȋ��?��ʃH�ǖ�<�ގ=#E��T<���5?G<?֮��$=�$�<&�[=�+b�=OF=�Ǡ<�+��/��V_=����B�x�A��Y<��n=�軦�K=���<��:z/�<!�H��8���R��x�<%�m�;���6*Y=+�|�ض����=���/1�F̡<�b<��<?)x=�a;;16��=<�Z~�/q/��y)=k�<��>=m���@d���<��N�Zl�����<��<0*=�`���%=<;=�z<�%9�?���ħ���ۼ��<߰�<�<D�F=��ͼ 搼-ab<��`��$���%< �=��<��$=�w2=ϛ;l�����.�l�l��>,=�u�X�O=�\��Y=�����;�A���ܼ��=�G��;��1=I�<񐡼�<�I;�N�<b>=�����>$=��D=��<@�=%�;��j=~��7�ZS=�{o=S�0=I�<x}��n|ټ;�^�b���2qN;�Wż�;.=�����	=2������wS=�[=D��<On*=��\=�hA=/nj;Xf��]5=@Dϼ���O:�	Q=���;��J=�A�<5=����/�K���O������e�j裻L��<!ɶ<�=�]�	=��Z�?ټ�.d�:L+<�t^<�P<U;�<�ͻ'=��G=�-;�=�z;<���O���;�u<���@7ػq5=mu�<8:=w;�S-��/<s�=��=���9%�	=�Ƽqъ��O�<P�&����o���$0�0S���B�W�E=��/���C<f�t���������D�<�e=�=j9�<�V�mD�+LY9N�=�K��`�=�$
=$��
�-���<lg]=�-=�q<��<1l<�*�<�7�<{��<��B=��=nԱ��>=u�ּ��<3>0�S�=�v�<G�=�K=��j��٣;�ۆ<�r�<�Ud�� �;�?��(4��7=�DP���<��Z=U�<�v��-�,�>=s��<PG�;�E<��=��S<����88 �@�< ,=a�9�_��<�gF�E#�<+=0!�<�"5�/,�;���^�u���	���<�C��1n0=b���_�<E��:�=��u��uS<�=Q�g=y���Z���|c�wj=���^�<�hu=r����V<F�̻��1=s��]Q`=Z�Լcx��Ә;;]�@�d",��E`=;�s�iK<�^����=��g�[B=Ym)=�U=�1�yK
<1��`��=frS��e��=��t�)=����R[�mi����<n��^�Z�rg=s�;�&��|��.�y�NT2���<�����q��;�>�<�=�K;��*=)5�8�.=����P�<��g�5�b�� �<��;��V=��Z=�_����b=]^�<��O9����6=X���k���+7�=��<�X��gμ&ڼC�^=���'��B=�J�#�#=���T�ɼū<c��<q�k�Q�ѻ��7���_=��=��W=.w�ݝ<Cm�� �=��=BC�Z2�9Z=-D<�����:�L,�),�*w
=���<O|��$�˓���~g<�v��z1=��1=�^D��[�<ʏ�0��<����S*�9��<	����<��.=22�<cR�;693:�׼ks��|	�9�h<�ч=��w<ݬ��J��=�o=� �<~8%9�&3;���<��;q/<-�y;�yY�m� �D�<|7��u��!F�<ۊp�?*�=n�<~�q<��=, 6��*������R=�q����s<"���l&=<�o���*�d�*�4y��_��;N:=s�<kp��G�r��r�<��?���7���Z�Y�I=�M=��)����<�Y;f��1�<��� ��@�Z�d�R<#E=�z�-�;4R�(?3�~�ͻ�+�<�=�;�H�όZ�T�bځ��˲��}P��;+��ᠼ��< _s<9�c=\�=�D���d.=�B�<�ɻ�5O�x�=��<��Ƶ伍p=
�K��0����¼c0S=��<���<@3g�豈<��5=i]a=$$���
<���=�B�Лb�Xq�E�4�M�C���1����<P�5���~+�ʅ̼�T�<!]&�<{�<�mU;���s��;��6�:E�?���<�r�|<�?û�3�<��*�&B,�a/�<��5=�EF��cw��ƕ;F���_<zKL=�s;�J=;�Լ�=C	=�8�A�1��y��؏�[�#=��";!��<y���W޼.�H=g�&=��<��b�6�0�Yd�<@ެ;2��<,��;�t7=0=@���<-��5#p<H|�<ʢ�<q�<�N��S�<��Ӽ�g�<\"S���P=w�<�$켌�<Uj���!�F=��h��18�8R���=��:9�I=}_g={&����=FV?��m��q1=��\�:TW�+g����-� ��<���<>1K=_%˼P�⼛� �}��=ټ"r�;�Hȼ�F~:!�<'�g=\�J=ɩ���$���S=��Y=~�*�<s=�$+�ma<?<˔.�&�y�j�<��_�#�ؼE�l��.�4��gc� ��<� ~��ﻳR��ڃ<�׼o"=B4�bhN�Ϣ�:EO�<�,�i����&��64=��_=��<�|]��5���?�ç1=��=x=�K;*��i�G=�[�SK�E�C=�ze=ѶL<�mJ=�C=ue�2�8��鼝�N<%|z��X�3=(��%C=�Y�|��;�P=���<�7=�G!=�T�<敽0���C�	��Ud<��6�H]�`�<���=%���^��� �<x��f"��<�M<Q�`=۵3=�;M��2R<4+�N�����q�D�=L��?��<¾Q���+=J��ȷ�<W�=���;n�=�A���6��=��:��2��Dp=Q��<5쪼�;=ga4�lʼ�H^�V霼�4�<?7v<�����EK�BT#���鼝�2��<=h �=�0�Z	=ع�k)��F<Gռ<�#��("��!�<�旺
�ѻ�U;��=��˼ ��;UV=��;t1��N��H�<!��v�{=����V;h{���h�u5);�#"��Ϡ<�=��Q
:H 4�HLּ��`�t�;=� ٻ����2��|<�:�	�<
`N=�W�<�x���P�n�j:�C|=����wi]<�%U<qe_=EZ��#��w���}V��'k=�RO=B2���_=��<}��P�;��<=�#U��="=u(�	��=M��"x�<��[=7��<���'�D=�;5=6=nZ�w�=����J>�n\���L���.�=&�2T��T�Z=cL��s =��3���<���<c��C��Z�=f�8�9��<]bG=��!=�p�<��?=���%C/=(�a�#/���?�Co�{IN������cdf<������<��G=��&�@Rb��@��J�0���i�e/�9���?��;H��<���<�a���-=&�]�&Kļ����`�=�@�����c�����<�{�UQ�r����<��j<��%=_�,;�WR<���<�
��e樼��<��[=�=;����<W�:=����$�_	�����J�K���<>�f��W=�^�<<�=(�<�;�#üh&�,�R=^=࿟��
�;l�*=:؃�V^;K�i=8�ȼ��g=��B=��<���<]ő<��;bb�<i`<�=PH�;=W=�ss=/9�;MH���p����;�u��=����<W<�i=��ۻ҄=uQQ����<���7=��<�Z;�%��b�)�4�U=�=�0E���i=vi<Xx�<(�K��2���r<x+�<*�z���:����h$=4�n=M�V<\s%=�D-�n�c=AK=8��8Q[��R=���S�<���o�=��=>���orc:��-����������<~�;R <�r�<�{D=��X=��]��b=x�e���k�B,=�B�H�+��<\�4�k�B����<�Q�; �r=�U�1B�<�K����#�������g=�Z���OT�t�={��E��Hk�-�w=� ;���[�7�<��ü'�<==��W���<�/(�����A�a�VL���;O�ļ;��I�4�}�<J������;oC���Q<��<ȏ���=C�k�����W=w��<aIû8p <�f?=>��:�y���;B��<�Չ�U(�qj�=���<9�=R��=VK<O��8sF��v�<g8��@���4���F-��P6=�0̼�-H�f)�<���<8_?��Y"���b=�»�4D��<�^��p����$�n�x������r,='q��SIƻ �K=t����_J<���<'�:�����n��*_=CfH������Ù<��"<��M=YsF��`"���Z��o��&�O=��0=�0=g=��S=7�q�<�޼͓;=��du���=���s�-��2f�<�A�<�e�<Y�1<�BA�c=<�]<Ǧ<��<`G=Z%9<f�=G{��֛�<?�=_�(=뜹��HC<��<.�K�nc�<��ʻO8�)|���C�;��"a~<LX<�/3� �<����B����C�.=&�����<n�!<u��</��;Й#��8��=hb���d;�y<�w"�},4;
8�1+�	.k=Xe�ߚ�;�=��O�#�=��׼L����l=\L#��v�:	�i<�T~:�f<��<�D�}g���"=?L=���{=,�!���K����<�x=�M�^@<� �<�hm<+Jh�	�?<zi�<�����{$��W���= =�c=Hs<Z�<�ջ�(=�p��9%<_<���?������<u���G=��e=h<5�[.뼵�;C]�@����K�<�c]������Y=��rK=��/�P	ӼW�=�9A���0��s(�c{�<��A�zMN=xB>�� <
K9=D�����8<9?�: L=��>����=�h=�c(<��_�kT�J��6��<�y�V�<:W��M�����7;����=�T3=Oż��.���@=��<x�<�D ���ݼg��L4V��v���ȼo���4<��z\ =*���W��&T=K�u��y<=���;��<W�N��w#=�l�<���u(=����ؔ��6y=*�/�'�<�Bʀ�Q�$=�z<7�>=��_=���<�ü�(ۼ&�a<�;����Լ917��w�<���&����r�ն�č�<[k���S=�k��=��<Z�<���<(m=:jѼ)ߤ��߹�&T
<-�:[fA=�ZF=7�<g.��V[�<z�=�ӂ;5��<eV���j�<.�Z<.59���;Y	<�+�E���<mt�<�8�; W�������D<s��<��6=�����T%�2��<f2N=�����X�=W���*W��޼��Ҽ��6���h= S�������=���|�k�vd�;,��<Z4;=dĥ=X5#�^=dq
�5k�;Y׉���n<ll�<SB7��y<�[�pH=DVȼ��Z���<QK��2?��=��9���0wȼ��Z����b@=n�K=P�2��[ļŨ1��d̻I�4��C=�/2� �W=�P޼�Bv��=�����e�<2�z<�pǼ��ڼEԼu`�;0��b]=�0?=�G��]�<h���b}�P��<lu�K�I�ID���!�>S�=�I=Cx=upF<Y���K�E=���;���QX�<���<I���"�9O=�����<�d�}���<[	»�	&��!��;k�<�.,�rGo<����*�II�2>�������<<��;mh��e �i;B=�D����K;n	�<�FX�X�^<=�R=P�%�XOB���;�I���J�<3
�<"N=�컘��;�=��ټ@71�}�'��F=<�����|)��;g���f��f�<�@D=�u=w,V<���Y������]KἫw{� �T��A]=SU�<$�;�b=��(����;��@<Q�@<Fc<C�A���<�>��g��΂��r�]=��d��B8=^�=$��<L����V�<������ܻB�<N>ȼ�1��F�+=><�S;�(��;���<3�c���<?N��U�D<��%=0C��<y#�O2=Id)=�6��ZW��<��I{S���9=��<�A9=�D';���O��<h�<h�P<O�J����/�{i�>�%=0L@<�*~=��a�� ����������'�m< Yn�#��?}��6Q==#="��:x�D��Ko=ɽ����:ս=>��<|й S�a�c�����ᄙ<+��<%�7��^(��$L<+�	�I��/�<<:=��<��<I2,<�v=��J=N,.���,�O
������i�ռ��L=8�5�Fm)=�P=��<Fz_<�.���^t<
x!=1� �ڊ��&=*a�<3��<Zb4�,Y��W��<�7�:�����=�33=�Z=qQ	��ފ��f���)���T�</�:�%�<��A�K��<W	=X�N�d+=�4߼!?�<�w�S)¼��=#7ݼ�)����7�<btK�s���S�B<M/U���]<�{�<�M�=���\�<�~�<���;�ü�tA=2=Dh=�"9<�c�A�%��<�Q�<i�D�o!�fw=��=QTl<�ڼ:!^�"M�'������c]��+�<�Ǿ<����62=�-Ҽ����W=��q=�AH��G=��
�u�Q��=�<�
<���V�#�04N<�v�G�*�Q�=�a� �<cE�Ri<k�=��X�:�#������<�
B=��7G�<��a7����<<��3<;䷻��<��W;��2=]l�=�Qk�W�q<��*<��a��/>=�m�;=�/�P�>�����%��=0������1<�(t��a=���x���
=�S��k%���=k����=����)���<�`�=e�<F��F*?=���;�t=��<R�༜vk��;c=¶1���H���Z�	
H=�Mȼ"��<�#��{����K=��9�3=,W�<�܋;�E�;�<��=�>;�����M�J��:9�e9S]�9�=&D}�F���5<+�=��n�<5B9<4Ͱ<�ټ�"���=�┼��ἀ=JP�k�<~��<��B�L�<����^���\�L��?�;L�I=P�ۺxü74�<��<�\p������ż���<eg��J�vi=.�p����<=��<��;Ϧ]�a���txI���	�KK�<C��;;O=��<��{�i"2�tW���r��v�=?o�<��:�<y���<�:T=�� ��<�:��]%<���xq5=�;��B��؍�z�:�p�<)�=�VK=p�;s�a�Q~;�M�����:��I=� @=�Iz<�}��d����LH��=�=��p�8i��j�[<�P=B;_=E�8=I)����H�/=�r2<�b=�h�z]�='�<w� =N0O��.0=$�B�n�7=h̵<�ƶ<zUE=�x�����<gq=!����W��ڄ<=,=67i=�zV=͂�񴏼��<p�o<��c=H�ݻ�Ǩ�L�l�,�%�q<Z�E<]$E:Z�=��
�U^	=�d���d��f<�\y=*R=��>�xbO���=��� Ӽ�A=F�����mz�<.Q��WY<Ե]<���<#B��<&_�K��<��:3;���t��62=K�=����:⼔相n�c;:�4=.�<�f\��$@�k�<�dc=��=z��< 8=3=O9�<`�r="�k<����5M������m=Ie��JRZ=t�ܼ9�A��,�����z�<=�W��#f,�W�<b�2�ǽe=��< cK=E3=\�<�)=Hyd�^��5=kg��w=�YL= ���Ci�?}��[�V=�����1F=cg�4Ψ<�_��3h=J�<XD�<��
�cJ<6��<�9+����<@Y<�1��Kw���6��+e+��A=d'�<D{A<��u�4��0T�X�#<�Pw:{�g������p=<_.� �x�4<��8,_��.^�c��=2Yc=���*�<�Me<aPz��wi<�t=JN=�ii��Ѽi9�CT�g�ڻ��(�È=e�=>5�<k��� �=o$뼕dB=�!=���cuؼ<F��(����<HVS=��W<�<�ȼ��Z=�9�<\b�Giǻ^�����ЃS=%�ͼYgZ�gp�<�⺼)=م)<"�����=�hD=ޡ;{@<A>���bA��E޺<�e=�i��޴����<Gh��	<�?=�j����
=g=�fC=K�"���=#��;_��<��<{�/������>A�IE<��ü�=%"�;��D<�O�^J��K�=��
�->`=�ri=WI=��j�:۞��b��p������i=̍<�i�;��=ݒ�;
�<�sD<�<
=�H�-�Լ41=�6=k(:�z�o2�#����lX=}�=�F��Y%=&�=n/A=|��~�<�;=�:/�^8<����<��H������?��<�-='T������_Ƽ�]�_d=�n�<`:�ܼ���혎���<���:;%�=���7=�U�}=�0�U#u={i=�k=B墹�_F���:�z+�$_=P���򟼊M�;�z��g�<���;Þ��)Sx�Vi�#t�W�'������:��|�����n�C=LCM=��n�t �t�m=�M��JZ=ƞ���P=sTW=.�Z=�J<2D=%;=��!����;�wq�%���=Ȕa���;=���:�7��kp8<��1���<e��<
�)<�l(<�����K���I��,A=�͗<�c����Q�2�?_j��n8*Qc=�X�����2u��d�|iZ<K�]=�6=	%�<??���=n"6��8��ּ�>=�+$���	�Z���#f=�$=ߐ�<'�B=�mz��S��1�FO�����0�Y;�.[��Iɼ3.6�S��I=7[�<�J3=�4�L�����<E�=�*7�zF��˼V@=�y;��<6˼�Ek��,8�h�v����<�A"=I¼�N��j	 <�8=B�=�`�<K�<����<�N�<�=׌�����<򔌽��㼲�=�o�<i�v�5a=��A����:K�n&<H�4;H���<��&�=�m�M�#��p���!�<�f��!0��P��;�X=�N��\$����\==��s]�<�h7��J&��<�
���푺�f�<�<l�D��<���;��6���<�|=�sQ=_�;Ar�|����;��_��x<�>=,B=�j:1��<�́<D�_��:���ļ[U��q��,��<d��o��[���Q�}��<R�C�.�~��E&=}q%��0ѼD����<�K�<��m<��ݼsa=Ro�<�'���`:�N`=����<�`ؼ�7e���	=�v�<f����,=	���N<5^�?�(*\;��=ݽ���9��|.<}/=���<xx"=�����%�=7=��W2��"8������	=t�_<ix=�`�C���W���3=_*U=�%���<�<��+���B�'?P<�L8=����Z	=h�3=\�-=��9=2�;�&Nf:Ɂ�-?<�Zܹ��;�@l��&z<F�<K�:<#6=�[�;ߊ��A�B��U�̒ʻP����9=\=3л�m�<�O:�>�E�9=b��<�w(�O�th2��}W==�<S����<�CE= ��z�R<��3�)����L =y ���m;NS��6Fo�6�<��?=��<���<L�<��ɼ�V4�tT=
|��U�&��̯)=G,#=JY��H	�7̬��wS��f��&z�?)��<F���&O�v���2\=�y$���Y��L=��⫼eQü~a�<z?=�s�;��A;��4�TUg��P=�Y��m��<��"���_���D=N�h=٭<�Xj=���<ղ�^fb� �"�����U�,�>��W��<6sO=�\A=��D=��X�Y0<�8�.=�0=؂];���
p�<��x<o��;�&�,0=�X�:��D�y��F�`�Z�����9=��t�*ü�G�:����<tƝ�_bɼ���̯�<��Y=çL=�e=�s�:��D=�-����</a���L�93o�<�)=��-:�^�_���@&�<v0=E�n�G�=��_��Z=h�1��"�<�8��m��<�ۜ��y�<|�x<!z=�=�=��n=��V���7�� �<�+
���;BDa=�=�Xq=�X�<��V=P���=۫���A�ڍ��=�9�<�=0=��c�џ<������<��a�?<BEY��!q��u<��;����<�#J=S������X1=Bx	��X���G=�����l��u��=�u��Ԣf={.I=&��Ѱ����D�$�d��~9�/7%���(���
=��Q��iw=C�q�<�r=͑�<w< ����;b/o<3��<."���@=Q�����= #�u�;F�,<���;�!=��)=Wl=�W�6�=m<F3=}���/��� ��c_��(���j��N� �<��=��	=�qh=Z	�0iͼ�� 1=u�d=/S��"1�E��<w���c=�a%����<���,	�3'-=_D=N8<A�<�ʚ�� q׼���D�;�û	�⼋m<@�C�����[�)=�2<��8�#�v�ӛV=���?`��7�;h��<���<M��<��¼-�̻"�F���M���Y�e�=(N�;�Ul=N8�<+�<�������<�E�����"�Q;"�G=��D=��<��}=@�:���<i
��������y׈<��;�R�<[��<��X�2��L�i��2��#D�<q紺Q��<|�;�[�
Q+�=�=M�7��<x�軅4�1�4;�䑼�PL�+Zw��G��<(����<�[G��B����<v�W<�B�=P�ѹ9=�O��al��{�<W׼�<=\�
��Ol=�Ƈ<�o1=>(��A�E<�:o=%#L����<9�ռGܣ<خ=�=^�y�m8���*�;K��R�;�=�_�;D���<M�
����.w8<dj�<A�=S��<W�C<31Ǽ�S6�NN<��9���<���1���!���U�:�p9<��"=�\{�ͼmf�<B�=G�;=N�B��D��"&������1�	��<yC0�-�>;,��e�F�=�*,=�伮+�;Q��<�9(=>M1<̨���=��fO<�A=@�N=©O���8=� #<��x=�����e=�f^=Ḡ9��:՘�<I���C�;S�'=Ƥ漱zz<�{�<���<�@�[�9=J���yȞ�-<mD��]��!�<п�<�7��ѽ�����<3L=;`üN�]<y7�:��N<|��=�1?= )����z��<����#<-��<��=��d=��뼖~`������p�<�&*==n;<8΂<c�"=���aC�ϥ�<�D�;��l;�_�o�;�+=�W�<:�`=}E��٦��o��h�ܼ��9����<e71=�Qx���;`�c�v�n=�6�<3�¼�' =!�/=��=N�M���ͼu4'=P�<@x;�T=�զ<���U�6�^üp��7;=2,B<�i=��D.�{�i���);د�i�ݻz���=o�c�Af=ݜ"=��㼼�<�|)�l�ѻ��J�&W�< �=��0���Ng�mv2=�B.��N�;��	��]���-+=o�ڼ�+�;�X1=�ẐŽ��,ټ���=ve�<��<�$=�w=SC�e�=~�;�� � ��"2��<�>=��I=���<�)&�7;�<Ybϼ�;�{ܻ��f����<4PK�E;*���'�0���"�H=��,�k��c��;��Y=v)�z,E=�<rd�\�A����<9=�l�<S��;��\<ᤃ��p����<qn�J5P=Uc���L�i<�|��X%s<<�+YB�R�a�/rO�VL<<q�u=������=�*�<1-�<:2�<�Y�<BS��==N;$;z�=�������yr�A�='�-���D������\�;�����<�\�Q�ż��=�b)<��=�_ =w3ʻ߭Q�W���y�=�� �v�<^N�s�0<k�a��ڻ���<@=|�G=�A��.%<�2�vLI���N��]Q�2��;p=@CD�q�T=.�
=�eA<���<���<�p��wI�22���s��� �L��<.OU�}k�<����􃽉��<ՌY=�K%��l�<�6/�ڑ��xO=f�g�ar�< 0�<�8<�
=>1���e=8��<��;<�]';��9=]�<Z#����<��/�g��G<|P~�*��%��<ʗ"�Gg�7Ӧ<�sL��_����p=F�-=��A<�6�<�����S= �N��~v<����f�;I�(�;���:��?��S1=z�;Z:¼��h=4��<)3p=�2r<���<U}d�$�.���X�֟�=-8w��}�=#5�^�@=QVb���m��'�ZD&��{�;�W��h?��`Ҽ�����<�]{�W��=�Yμ䢰��q�<�<�R�LZY=�Jh=�U"=w�<4?μ�Kc=��<���x=��A<��P�������X=[�<ѓt=a���=���!= �=){m��@=|iI=��8=;S@�W,�;9A&<.�6=-N�<Ǧ;A��n��b�<��=��$=HE�<��V:O=⼅���Q��;��B=�#S�<�6==6=8hC=�=^�1=�׫�!T��벼���q󍼇y�޽�<CU��M=Xܗ�{S= �;=���<N3�;+�6p�OV#=�ʸ<���<c9=١B�s.�;��;��p<:�*=4Bt��n�<��=��_=���<��;����zC�}sh<�Kh=3յ�< :<��f_��Ox<�Wv��21�n"μ'�_<��Q����<��_�Q��<�؞�����q9=�F=A�3��~�<�8�4^��ds�bKp�rl��1=������<iy]=�=G> =q>��-���K=��<��=Mo<b�F��8=Y�=!*$����<��y=�RK=� ���=��<0t��
��	L�����LU�<$3Ȼx��f��E�=d�'=���<�V黏�; �?=I49<�ƛ���2�[q�<_�d<��-�|?�<�t =##H=U߼n����
��/\=T]�<{W���I�c�F�y���B��<k�=�6=(��<�~=[�M=��<s�
;�MI���<�u�=Py<�����uX<��=O@��Cg��=��;�=��<(���wH��E��<5)�;�֍<�=$J=�ZF��Q���=_*���7�=r���@*�:ټ�,R���1�=<�R���S:�l\�x&W==�;c>����y��	D�	.!�����~�߼�F��
�[r6��vO��5[<aT)=W�~��#��_!����S=��F=є�L�\=5=/�B�T����<�ܼ۽A=؃f=��;~़"�8�m����;=��G=|.��r=����ů</��=;�:ǼY�0�p;n�Ȼ�m�<T-<=I�H:���:{�2=����&=�:c=�_Z<�c;W_�>��<#�;VN�Fʺ�w�<�B�C�<E�<c���W�<y���E�<N��CG�|�=M5;=�|��ǉ/��pt;��<DS=ށ�<SG�f�<l���#=b��<����w�&��Z=������=��^�ݩ�;��V=PŸ;E|�]r�<b7޼~]{<��=~�:�����Լ~Pļa�w=J���c�j;�@�ܰi�ܑ�<�#��܂�2��̰�<�-���=*��1�<�4����I=O5R=�ԼC�<�kC�˿���J���!=9'=��<56=]� =��=nfg=^��<���c05�0�	;^�;Dll��IO=����E�;�;E�ϼ�F�=X�<���<��<=��(=�q}�f))= �X=��=�M�<�i0��ֿ<�/�7QһO� =�7&�շZ=o7J=�#=� �<���8��p��`/=x�)=KV=���Y���+d=�}���[=�'�:�z&�*��i<=��a;N�ݻ��<=�Ƣ�~�f=�p���1�IC��O=��;=͈�<�����<��<V	���?��(��A���u9�6�@�����[�7�x7�V ><�-�H;���<q
N�|n���`�;|�W�";n�0���;�No���U%�<;�;��3=��&=�i��2��i�1��A�<	t?�F�p:k �k{7���<�|�<-X<X��<U[=�Ѽ��!<��м�M�Q�>=�}�<֌q�F���N:�����pg=�JO�>��<�ؼ�<�>��:��� ���ܼ�X���$�x.x�1�w<�:��5��Eݘ��i=��3�p4	�5	�;5�%�i�]=�5���'=̖<*�~=���;;�<P�O����<-�4���8=�D<���<n��<c޼"Qh=��99�l��.8=G׎<�(�;~|#��c=`.����t��]���j[<l5��f��9��H=�7�p���Q=�R�Pp=���9�y�Vּ�h8=+M�/r�<��U��(.<r��<W}�;p���ғ<�x<=��<g-B���r<t�E�kb����Q�B=��<��ļSC�*]�<�H�<��\Ƽ�>�<
�9=wJ>�1��<��:=+�L�=r��;�8aQ<(X7�w���	$=٪;cֺ;*���X62:�K=(���n���ܼF�u;E�|�8K���!N�!����;=fM;PR׼��S��8�<|�L<x�꼓��<���<����B�O���q2;�]��6�QMp��/=������a�E�<�=����rN=,�<	��<�f�wqI���� �V=q=��u�>,�<2�=Ǽz�/<�L=CmJ=F�G=���<c�T���M���	=�}M=��<T~=��K�㽢;7%���H=k��<�:��7�x=�O�<�Z$<u�H<�=.*=�C"=g�:���"������=���~e��l9=�S=c����4Y=(���X��<�F=��G��nb�zs��l�=�\(;�Iл��"=�T�;IL�<sm�<��K<r����s���1�9�J���a=T�$����<Q�%<�o=���<�//���s)=	�N= `�<��ļ�_������	<{:=W��/3?�`P���`O�X%{��w=���<�C}��x=��=�^��Ğ���|�����:�L���
���O�3#�W��;�A�:H?�<`�O���(�]]�:�2�����<��	���<��v��J��Y>=$߅<�A��*ͼ�K���Z��z=v?���<d���W��,��5=�\<���<�X4=% =�Z�\�`�!z��<��.<���^_���<��c�Wi�;�&W<ؚ:���i=�����l)!��jN��<
_.�flv�Y�B��pz=4 _=��R=b� ��!�<��d=��L</zo=6���3y=*�<C=H�p=f��<U=����-"�c�k<��=�4"���Qn8�EG(<�z|;s��<%��l��"7o=���k��$߼�-�;�1��5żE=j�==_�=)�<�CZ=6��B�a�q���]5��j�)=^!>=A�E<i��<k�?��(*�z�2=�"i=�ѣ<%G�P�"������9Ҽ�iż�<Ϊ~;��<�4=�.��!���M=��%�k.ɼ ���f<�kf=���<�PV=ڼ=�I�[D��Q��<%�-=�H��rd=�w��ؼu�ּC�5<� �<���<�f��<��=
�;�^C=\z�<9pg=�:��/�GY=R�K����Î�=�ы<�cz<	Hټ�м6qѼ<Ɋ<ܷ= �P�}9¼g:¼9��<K�<E�<���<Ԅ�<�i2�Ok����%�;?��A)�@)�:RW8�Xg<ܫ��ϟ=e��h�);�P�<�z꺙���U�S<��<=D��=���!#���ܽ<�D�*m�<�4�����}�=s�e�?��<��p<j�"���3<�<�<E�C;�1����<�_<5غ2 �;DF�d<=���<��@x���B�<)"����t=Ω-=��<PC�;}�ƹ�q�</�;����:Q�`�R<{o'=)N^���'�C=�4�M����l�;P(8< �	=	�1�C}ܺ��;3�t<�X��c���/r�1�ֻ:[��ұ��0<83�<7y�<GqG��r=VTJ=��<�/{<�<ul������n�<j2=E�O�莰;}B2���f�n"�!;s=p�r=�6��ob��x���>��<C<��<1�=%�;�*��<=�I�;Axe=m��m��V=�9=Q,-="[9��
`<�Np�� @=��K=n����䨼xR&=�폺��]=1=�ĉ�v�<04=ų��P>W�0��<%�J;�>D=7�h��o:S�9=P��W�<�p��
+=·i�Va.��cH=	�P�s<	E��(R����;�N<g����&s�-���Y=��B=��=c(S���9<���<B?���w�]@S�u�&��>3��ψ<d$��#�
��9<�=��=�L�;{�Ǽ$-l��$�{ui�2*l�ߍo<u��}ͼM��Չ<n'�*	���4��K"=z@<'��<��I=�Ӽ���L�d�?�X=Ǣ<�v<8+�� �$|_=���!oD=mqἳ7�<8ٰ�x&�="2�I} �0hf= #�;ƨ��,=n�~=�:N������OM�CkZ����4=�!��΅����;�?�<��6=�SK=z!=�C�<EW"�I�C��]l���5�1ic��k_<�$��eD�a���ڼ�7J�����p�	=ʙ�;w1Q���<3�F=O�J=����8�<ɠ��@<�*.��'�<�re=��@�Q��<맻Ѯ�<˼-�\<,=��tE�]��< ��;)��� Q�<�P=�\�< �<�T?�A��<*����=2��yZ����,�e���<=�];n%�;������r�<N�D�\�>�<"`='��;)5+��o���~9=�8=�G>=כ�7G����;� �<�<���di=I�<����jL=���Y𘼺	����20N���=��Q�d���=Xs�ZH=@&�@�<�����O*����I�=kg�<6l)<;xF�����ƻ�/�<OU=^�R��?A=(�.=�&+�n��<����y#=;r���K="�4�u�=�f+�7��<��R�G��tg=VW�<u��.�e����<�e�=s��;�;S���=��<�l�<4hd<�@�<a�4=��<q܅��޼u���
���lQ;w����%<� =��Լ/�'�5��;4�̼HQ�<�?-�Y㿼���<b�&�eּ@5	=�Y����ݼ��N=�(�;�P����<��=��:�+���;�A/�H���r��<Su
!==�P=���;Ó;͛���&!=3=����X=��:z���;m�m@\<"Z�<��*��h&� �1=��h=m�d<��)��<}���72<�u�q�Ʃʼ*���|=��=m:��='���m<�*�O�H:u��vD=�(B�L��_ż�*�<��=<¼Ơ���+Q<�j���',<m��<v�w=�n=�2ʼP��=��=
H'�r5F=��?����<��P=_Wn�F�r=�t=\��<��<�����j}�Eu�<g�<O0U���&�/�m={�P=t=~�Z�*�=f���n�o?�<���<�Q��7h={�;
�R=�S���=��<�X
��%�h���%��bqP��"7;��=�~�<S���V>=W��������ڇ<�=��F;�{�� %�?tZ<O�Z�IA`=:�¼}n(=W�t�i�;����Ʌ@�6�X��ҁ;ļjb�J"����<]�T=Z�<��J��bk�-C�,r_�|}�<6�<��=���+=9�0<Y	=��� �:��.�u��;�P=�:j�g;�[]�Vt�;{缼L������2�<+�J���Q�4�$���8�=ku=ݏ=��3;�d
�����4=��_�9�L4�<�P����<¨k<���<Uu�7�;>E=�ex�I�<0�<i�ɼ��u�`r1=��(=J4d<�<w���=�R=b]2=ˁ�<�G=].�;��'<��<�:�<k
���6���9f�<���u+�<&�{�
Ǽ��!���|Ƽ��ټ5��������/��=	ck=w���}����1=���<G������<�r=0�P=�W=�W�<�̼2^h=�%����z<_<=w�s�;�
�K�==mzG;R��w!�9���<�C���<���7=ȵɼPר��{Ӽ@�)=!�s��Z����5=��9=�Jͻ���<O�����Q��y��< }��.���P=�c�G>%�+g��F+=���<�ù�ϝ�\�2�l��:��<U�=�K=t�<=��?!G<)?�<��F�����+4<��=�=�G�<���;:T�;�ё��2�<]4<��+=�`Z=��<��Y�ù!���
=��Y=�7=�͞<=ܺ�U�2��|�v�I�O=�U�?=$䂽�3N=:H���-=�z<��
����<�=���<<�X=3-:������M=�:=t�=���q�R��cX=be+=�����=�5<���"�4>�<ؾ�<\Ϸ< �C=ڋX=�H��?��vf���<�����u<�[�0�p<,��< �ջk=�I��ny���I��E=J�g��;π�<���;�N<���<*=Rȼb}�<�/=1�<|L�:�=�t;=�f=/Z����8=�	ܼ�숼��=;����R�%+=v�<�;.F=7�u=���<�S�}57�����:o��|O�/�o�c�<�S@=|�=����NR=(�\=�=9�,;~ I<bAg��:]=�s�<�I��E���D
$=א¼��b=�/�N���'�;>l;r�s�<�=b_=�'��3I��3=T���w�g��=$���";�<��G<�E=KaQ���g�K�G=4"�/���M��<�EƼ@�<KW =Ⱥ;��h�^�|~]��6���;2uj=�.{<�<�^�62=֣��Ο�����ϻZ~�<V<�<(k(�����0�:u?�<��`=�K=��%���<��=�)G��8�m���h)���ꣻE�4��<����h=�� �9u�C��q���L�<�_�i]=H���g޼�3�5�A=e\(�YD�<k�H��P=$����S�.]=����|f=�tT=X���1�+Ǽ������<��<�<��=[i<�F�S�x�5t�<�����뼝�ʻs�<S���X��w= ��;7��|b�;xQ��M�1��<�nF=Y��_o��H:�R����@s�`Z�<c��<�6���(�<k��o�ܼr)p;�xD=��;<�����q<8�&�ó��_�4��o����<��N��5=�3=�FM�I$�<�g!=�d��C�Q<jyJ���X�Ed=u��<�9{�U�	=�`�<�H�����������G:�Al�<�=��W�9�T<��d���5<��z��&'<R�i����=gU��ü�<�'=|�<���q=W��zV=	u�<z��<]X<
�D=/�;=�[���N��<�<~R;�>ļe���@+<Y�+<zNT=��`a=�����=Jp=��0<Z�;@�����<Z�
<�;�L#��`=�	�;m���B��IB�;���W�6�P�.�K�6dP<�aI����<�퟼��6����;B�s= !p���R=��"<k[=��<�/<=p�_�a�	=᤼��*��7
=��<s���{p�<۟���<E��<��:���S=�fU�썼Y�O=>6���$�N�ϼ6�<�+��i�2=�Y�k��,\�~������<!�F=��8��u=�,m=�,F�
8<=M|������3=��<w�M��{�;C�V�#�=�g����S�C��<��-�� �5+#=h���s<=�ە<ϳG=���<�v޼��b���&=��[����G���{Ȼ�8� ����c%=l�:�t=Qª�cj����f�H~8\R�	.������2�l��<�Ų��v����<wG��:=��ؼ����?�<j�D�B�C<R���~������$���c͂;u&)�nZ=ֈͻ19���2;��g=lN���8�7�8=�a�ur��q�<(�*=��4�3X�<��T���k�Mpd��f8=﵈<x
=���<T�輲����:��o�P�U1�<�=3z<h8o��e��KfU����<I�;%:ż��J�x��S-�{^�� =eem=���<���x��<Ƭ�<�`9=�.A=L��� ����T��=v=v�%vϼ��=H"A=�Z���伴�<�˦<�a?�� =�3U=��^�O�=�rf���#i=}f�<��~�{j�;��G=�TL=ԇ==�W9���f��Ǽ�g1�õu�V�=_> ��ʬ<f��<#�E��{ü+:=/�<H��<���'�:�޾X=�5��Y�==E�<Q��?���Y��.����11���Y��=�
=���;a��;,��<��Z+�rA�;�	%=y�`=�' �J/u=�̀<�P���S\���w��4��+�=�/=�໬J:;�<�M�<]1b=��%=P+=��<Ǧ�<�mM��}�p���������<N�q<����4�<&�G=�[����^��(=_�'=�!�#.��� �����+aR���ڼ/ "����͵d�8���(dy<'��<T�b�bΫ��RJ=��ܼ{G�<Uih���B�n�7<�r��1�»Z��<��![=��7�!6�:����`�W���aT=�؜<�&�a}S�h5� &=j�<��5�;�+�<J�T�d0=������<=d�[<[��<�v�<���3L;�m��*�j�Y�3=��<=�rH�$����_<f�2=x�/�����������:�*=O�P=�����D9��ϼ�3��P<1_��}<�\�<���<1�A����<]V=��w(��͏=�3��u��;dP��0=�3�;k�&�z=�W�<K�<�,E��H�;o#"��nl��Tr��H\=hqٺS弽O7�)�b<`��6�:=��^��l����<�&Y<w�@=q$�<��@��3M��6<����0a=lz� W��d��8=���>�<]�J<_C<��"!����v�Ԝ�8b�%ϼ�0=��<���<�N�W,��0��*�<4�-�²üt���8�2���=�:�<Z�=eB�<u�<���!0:�[|=�<�<A�g<�V6���<��<��n���=se@=�2�;�zb=l�~2���5=#K+��ּ]����>��$\���<�.;=ܰV;�8;��$�4��<�$�NqB�$6�o/8��j5��P.�t>A=,U�;
�D<)W<�%�k�_�(�@�Y>����]����<�:V�� ���DT���=�(	�����&�8��c<9q@=�]��Y�d<�><%���s<��o=��<��<o�4�g��<�'P=.4S��}��\)�TT��<�D=�\<X��Ϲ�<����z�P\#=K�U��c��xs��a=�sK=�: <5��=Ǥ(�����/<��{��<׽B���� 7��i	=��U��J=�{�<t?<ZY��N���y����8�dZ�!�S�n�9=�%��>���?�;�>v���<��>=Ok:�O�K=k���N�<��޺6��ϫ1=��<�9=��i�5=8�1����:
؜<z����(Q=?p�<	=��a1=y|�+�-=���=_3=���;ػ<	=�HQ����,��[� U�?*A����}:=R 9A�:�G꿼��a�?��߫2�@?�ɨS=�-*=�`&�?��<��M�I'�<9
c�h�
�\�=w"��9=É���K�Ρ��F�#;.4��},��`=�qԼ�F =V�<��5�8Y��Ui�%�D��V4�=zH�X�:�x�º3U���<7���[�O�<����c<W�=q��1��;k���>y��D弲�T=l�;��/=x�x<���<r�"���;3=PE=����7�	�b��	O�K�@=ٮ<=�{�1�s�e�0<=���W�<���<LS�(~�<�*7��$^=���<we5����>�4�r=5�2<g:2=-��;�\�<�9���W���`<B��������oK<(�c�$X,=���<�M=�R�<��<Q�������>�,�����i==��g��]p��*�O�I�
�*.ټh=��5=��<���Ӡ�A�Ӽ0��"<cN��͇�����=�( �h �<&a��]S�2N�<�R��CS�KcG�T�ݼ/[:=>�B��=��l�N�S=��7�-I��E��_�<�a��L��w;�|{=��<�T��<�3p�<㟇=�P=3�y��0̼���<]n=w�R=W�������)@����r='v6=~�P=b[=�ZR�#NC���^�u��<n�<> +�����ޮ��6=a¶<��A���Q���L��D�;@T<�d����!��<�n;��?��R�y��#6M=�4������\=�����<�}2���/�aE=�+N��=bv�<�u ��'�<D,=�"���U=��p=���<�d=�l=#�W� �<��<��|;�<�{��(�A�m;�_�<�/v����� `j;����)���<�<4��79G<A�»]q=�8=�(��� ���;KDc=��N=F���.uT=���<�=�w�<�M�<0ێ���:ed��-�<	 =�M�<\&�<���<=J@��J���jp�4����wd���"�*=(����X<�P������)=��;;�=)yؼ�j;���:Ld`��-%;�����`�1A�:�����r=��c�=�S=54�&ỵ�L=ZD����:���T���6���,=`!F=���<��W=�|l=(J���?���z=ťH���T���ݼ<�ܼ���;�U��]o=��<�M�iXS=�q<� �=�57=�b$�jU#=Jv����,��<޾�;Kx�<q���
;+ E=��<�b=	��;Fc��}�<���<�i�<$0=���<2W���
;�.�<�?y;v�
�� T=��$���J=î<��F=7��<Ai��\�;�1����(�<G�+=ϧ���D=��+
���<�<%�,=�F.��q7���<"!=���<
�\�P�I=D�<�U_��F��e�V=�=C�<v2=� d=���<?���F�E@8�#$l=�;\=��#���:��U�� �<W3��D>=��=-�����ü�H<$f1��U�<c>=ߥ2=����w= ɿ�� k=.(=�KA=w_�/�9=Q�Q���~<��m��μ'}Ҽ�e���������o�<�"<D =���-H��f ;=+�ށ�<��"<��<_�!=��B���f�{�';�h<�}���p;
�����<�WV������_$=/P6<fF=c���k<�Ih��+o�+H��7"<U[ؼ��J��ç��_N=R�;�Uؼ�ջ���$��<�+m�b����n���<#&�q�⼹|Q��y=e%M�{A*�Gn��o����'=@x;��<��;�܀�ek=~ü9�U�ǌ<��,=r%�;� j�|<@<�4<$~=�=�n�<���;E�m�Q����"v=��\�~��<�򶹶��`�<{uV�4�=��*�P��;0�6���<�fg=�ѻ}�+=�<��/�;�S�<J�<a�G==��<����n�)D}=�ܺ��O�� �{�k=�82=u�U�2Z=H�!�9�<R��<��2�ƈ�[�=�4=�}3=F��<n� �����O=���;�t=`TR�Dk��B�<0Ya=�������C�;<��=>�#= M<7��<-�Y�K����[��)�s=�?=DN=��1=��==J�0=�A=��*=�Jù��=t-'=-[�<U�i=Ŵ9=��<��e�<zF�;Fh�<v=nn<* ܻ���<@w=�W�:�ػl$_��>=Ps��>�I��_=�Oμ��=���Z�/�$`H���B=��,��'j:�
�I%!��S�<'�$=e�<���;X*�ZM.�O�=���&�f��������"���ƼNI�<||H=�
�<3�1=��W�E����3=C���I��<{qC=�,o=��<NLl�*S:��R�	�e��%&=l伱N\�o���9�=s#I=����"fY=Fb���]�;���v�X<ʻf��i�<�;h�� �;.���<&\������a��x:���a����N�x?=�/����Z1�<��b�?F=�(ż�m�

<U�m=tP.� �,=����}G�xz5��R���x=u�<�����G9����e��5�<�,C��*;=&�Z;�F��v�׼m�,���<sx�������Y�<lT�P� <�����=b��<��^=��黅@z��=[#���Ӽ�H�;/�J=��-=���9e�'=(�;�(����Y4�HFJ=	 <<�<�Mī;ʳ�<��K<���<�;���&=a3�=��<3�ռ��S=��ʼqAz��T=qm����]��1�SE=��<�O�<9���)�T<"p�<.c��l�N�<$�g=��k<i�<+�<1�˼�:��!�R�� =�Jf�jE=��Z��u� =�ڼy����v�V�<��o��ZX�?zC;���<ғݼ�H�<(��:YO��ca=��=�77��ڳ<r ��g��<�r4<�� ��<}5k<`Zk=��N���=�͋�	�U=vjh;�����U3<s����-����"�\/����2<���;x��)a=��*��=�m��8�<�q$�4=*��o<�]�8.����<��]=<"�<�@����H������Ջ����7=�_D�L�C�1�׼�&=��<z'�j\<��9���=�<�A�=���	=��=]:=��C��eC�1�漴�7�a��X�l;=�u��6�;./M=�Y=��<���kZ�-�<�w��`~=�6��n��� �=$���y<A0�*��<�Kb=�)5=�o�<�1��۾�9/ؼ`�j<[���FE=�|��,3���.w���<��F;D����d��*�����<��?=Lm��+���`;C�V�����ie��#4Q�EuJ�G��<E����� �)�o<͞9=&�$�]M`��=P$3�Ϗ��y�����f�˼�=�@��v�
�[���s<A@+=�<�vü�/�;P�E�C]�<m]��;��13i�]�j=q&=82~=7�6=9�o���	R<�3���<@�P�1�<�J�E7=|'=1l�<�;P<�H��u@�����6<K`=�Ѓ�l�ͼֱ2=��ɼ#�=hy���P���]O=�=��6�B=�ɻ�p�H{*=�7e=`��%h��s�L5;'�=֤V�GU�<t��=�֙<h��&�=�=�@"�*���}-�DeE�ǒ�
�k���'��Y<���&c��?s����<�S.��x@�?m=N2^<ά��ޕ�v��6o�J���s[� -鼦16=eE?<��C���v���?���<]�����<�c��m�=�o���+=�_1���(� ��@�;=n�@��"<b7��z�<W/༷"b=����kY����k���/��J;��eX=YD/���=�2 �bF;c�=�G�;%S̼6�!=N�o=]b�<f}輪�@�*�żΨ=Xy0�6cX=>�B=�:�K��<�����%� �Ѽ���<QzӼ�
��DK�<�'�<U.���=���c�K��=p7P�9�ذ%<C�s���"=Z����~����h>���R�K��<�$	=+��<>U�;��<��N��
¼����B<��3=�%,�{U�P5��0�%��������������9��x&���U�E�9=��6��=�/$=�D;1S_�u�$��,�9Y1=��!=�"=�_Z�=a���Do��~u��L<=~o<� �<��!=z�'<B�.=Nc�"��;�ձ�y�ٺqe�~�=c��<�]p<��!��ˎ��֤<O
��h�.�o*� "�<@E<EEG=1��^Q)�h�Y=�t�:XH���B=jv�����<+Ί�05=NMh��ak=�0ϼ|�D=<��g���u��<�Q�x�ͼK�m=��=�W���[G�;n��ct<^H���S��6<�C���;�D=^<6H6=9�d��<;���<Ih�s܊��s&��;�q��O�5=�9��P�b�aE&�N[�2��(=w�<-c�xG�;Z����}f<��<j �:�=fˉ�v�V��'���`e�wҠ���Y�A�<�jL=��B�1�a�?�*����R���� =���<�=���;�в�Q�%8>�-���P<Ǽ���;uD���f�<m����=��=]=/�W<q�J�31%;t�T��V�<{�i�J��e��;���?�Q���5=�q�<���<����M�=»���B���<.�<�p�I<y��[5���9;=�G8= Z*=�3=��㺽�C=`5&���=�y�˫L<�8�;4��N콼\5��a߻���9�B�<�G�<-z=�j���V4��#ȼ*�»��7=	�Y�����r�ۜ�<�Ἃ�:�B�����<�>#=����0l���.=��ͻF���4=�P ��Y0=P�@=`�=��%�EL=6$;����<�M�Q+�<�j;�;;4��<��*<���<݀��C�/<�W��=���q@���C��=�<��=�9<�<?��*=e�%�"h�3��<��vr�<!���<h|ü>�7��:6<�/5�mn=�W��s�<G�򻤸-=S�<�z;�H=��=��=i��G<�pԼ �<��C�;�=�=�bM<��^�]<�.d<�_��C	��[�>X*=�K�<��=&�>�Ѣ7��d��%4=�!�=@=�x��l�<�����n���l�$1��P+�RA��;�=d��<�A�:Ά�UB`��jA=����̭<�+�V�}�tƕ;�Y��3\=x#��)D�<��K���\=�jj��
7�6=p���F��Ih�N�͌=���Lܒ��O���m���;=�H����)�b��<9���@=L�v�N��;R��<$��͐��R&�����8U�-� �2�v=�r��zCG<�"�<BJ��Y	�t\`<d�E=GO��8s�<n*��|=�����L��U��|x=U���N��;��;���5�<����뺊��w�� ��;͑h�� ��+�l=��<=�D���b=V�h�3���9��P{= 6�Y՟;�	�<�Ġ;Dgo���=Hb=1�=��K�y�<Uv�8�;9L6�/>�9�C���<=<}l=��x�@�B<!�);�긼��Z=##���n���O�%�7;x+�;�`b=�J��!�����<Zu=�8��j1>���B=r�m=Wb�~YQ�G��*�X4���	�A��=t9>=-�A=���M�<(XP��3���;C۷<W'=n��<b5`=*��<��;p�Y�©�;@T�2�����;d��=lD(;����Wn/=/Y:�2���<��,= �\=b5�<�ا<2Y.=l����<�����0�[@B=�z�;���<_���V<.�ܾ=��K=�t<�"�<�#;���<p�_N�.k�<���<k�=23�<H��{��U
�<�(�<��ͼ����n=�j;]�<#XH����<��<O=S���f/�*�����<3�@���c/��� =��R�$�U��<0e=�A�#���Ae<<���<���&�=3�Y�s�o��Fg�v�¼���<�t꼈q;=����2���2�� �<���9�<�\��@��P��=\��#W=���3�!����<ſG=�i�'��&��pe<�QM�G"輦D��9���(=m�Y<��U�2c.= "=hqt���C���`=��<�
�TgM;S7<�º�=m�-�X<�⬻�EI=��<�7a�cx`����V-�<$��;7#�<�^��E�B�1<ֹ�dS�eR"�֐"�u�'���<��<�+=ֱw�[�=׽Ӽy����<}�%��h�ÜM<7�t�ɗ���{A��Ì=�D�L?`����M��<gW.��ԋ<��-=�޼]T� =]!��u��s
=��B��dʼy�'<l醼M=-�5=B�<�>C=n��8�L�����<��A�ݰ=�V"=��=��@=Ω�;�r�<�=����<�M�;d�#���C��I�$����uJ��S=wb�=���<��3��=�N�<>�+=�X�<���3r�s�a=��;=R<,��<�R1=�aC���=���<9�==�\=�.�����l�ܼ��?�����V1=��K�b!��`�="�=Ï�=�8`<��A=�'=��O����`]m�$=��@?�tP�OCK=4G��ZG��ڼ�'ؼ�gr��J=�C���j	��D=-/ �6�ٻ~!=8I=��<m���H��vǼ�R ��V���!�;.)==v�����g<
6m��
=��A��I�W���Y�,=g�=�p<upV�C�r={���#�&=	����A��V;(��x�<��Aۻ<�E!=L�%=]T���E��f�<�/����<���<��S=�a=�J�<��-;�:�;V(�<��, �%�8�W;	$q�� J��r�:.�<�q�<��?=�U��9*=)�=Q���%=��	���l=x�<߹�=�a=�.J�̓K���'=��<�I��%=S(u��eg�e�=4H^=��=�T���B���P���p���b=k}�=�{�=�E=p[伈^;�-Oܻ-��5%����:��W=&��;,�-=�����P<=k���ļ���<���<ܼ�So<¤����L=�_�0��;�^J��m��g��>�<=���Q;=��==
���s=]/-���v�1|�D�4h�ځE=������<�ʼ:�6�\t\=7s�g�H=���<Qt�<��]���x�)=���<u��ڱr=�mj=L�l=�J���^=�^=�V<2{��H�s=~���ۘ�{�K<��W<hI%=E���=�o:=���<���<:���s�;�Ȕ<�p=;�=��J�ӑ3���軭�/<}L<��Q��0μnA��ql="��;Gݵ<���<�4��Uf<��j=bSU:��=6̼�Oü�mL�4�=��"���Ӽ�P�<��u��r:<��<�1���T=+�=�cJ=&��<�`P�k���?v�<����O�N��MY�<Sd���=���<_���"7㼸 =?:�<�۬<>�v<�&<��=��~:�=�Zc=�]=�QܼgNT��-R����]Z�6i0�s<��<LM!=��f=��<�kY=zj�<xs`�>N =WB�<(�Ƽ��;2�;J�,�Y<����V�<z�<�}��� ;p��=��Ǻ;�����<Wqd��\<d/s��y;KG��0����&<����������S=>t�<�����<qU���	������i��_H<]�:�4��i�E=�d���< a;$m�<��=6�!=Dv[=�I˼k�E��=ސ(<hʼ���<�<��^=���<(��Z��<#��<Z =U�g<E�8=��-:2�;�%�݄A�|��e�����=�d�<�i];��o�e�9�nH=�TF�X��d�;:�4<�{�&�����-'�~�,=h���r#��=�=�ڐ�����4|��a�;��W=�p�M
=��=��J��a�E���ށ�|�T��d��b4��j,<��bT�<�C�;N�3���]<��7=�-X=K�<A�C����B!�;��E;�`�t]i=�2<�B�����^=t�D��-�r��_�=������U�,s������;�(�<d;}��{���$��貼�¼�������<L{�d�<Ar<i���h�h�;Κ�<U���Nۼk�I=t��=��<!d��
$<��y�Q�ʚ.�ܰp�nߓ<�L&��4�<�����:�pD��[Ҽ�6�
�<9��R=I�<�9�:��T	V=�H=�=z�0=�����Y=�%�^M�<������:�=���y��;�"<�J�G�<��`���%�`�L<�� ��Г�)+��6;=/��<�9><~t��?s�;iW���=@�ӻ��<w�g�L2����<�a=�F�9�?=@!<nI#=a��z6w<�p=�Ӽ�%��J;*k˼2�:3��7r�ۺ��1='�煑<Ѷy<΁�<>�j���O��#��y�'��<0 ѻ�
Q=Y�~<� (���%�L=!���2��[=�2@;(�M������L��6=/ݏ<��K�;3T;r�:�q�:,O<�x�<�"��<j|<=�$S<-Q�na=������.=�OA�+Ҧ��Q'��W�|�򼕔*=cNT=F�Ǽ�3����+<��5��=��,=l��<�?G<U,�;��<����K<��=O�
�c;=�<��}��в�o��<��N=�c��Lx=�,�f����p��Hz<�n�bZ𼯿4=�%i�g�9=��.=օ:�Цj=���:�]���JE���]=~û�w]=|5�<����<��<�p�͢�z��<��Q��QK�S���zT<΀H�t�U=�]��s��<"T�PFɼ�;<�i5=�����c<��{=<w5��l�<�m,�k<b|y���u:�L=�U=Fl���8=&=xo3��'༘Q*={��<i��$�)�Ƽ�2]=��<��<�̻� R�m��\W_=��q;���28�<��i�g�<x�9.�	<}`=�2=)E�<��<]{�<a�Os��O=	=��<��<s��<I*���=�4����<��F=إQ�,�4�/Z��������<��=�G2=֧H=h~=�m1��)t<G�<�=�����Lb��G�=p�4��T����
=<4<�i=[E:�C������C�;���<R�\����/���<���g+�<�+<ęC=�`?���`����<��t<$���*3=b�_=�At=Q�U�830=G+�;�k���Q=��<�ۼ|A�;7ە����eRB�Y�%�sF~�lA�<�6=s�={d�dF=����6�Q[U��~z�F�z<��V=�`ļp���v����՛}=�
�\�=0=�ԼG�7\=̦<��%=�m�=��;���3(�<�m���<CS\��K=��P�	aB�[7=@!�R��=R㻟���5<WI=�	�;�*7��O�#fn<c��<�x�\Ǥ;R^��{1<9�;���<@�6=Z}=+�<�ټ���=o|�<(�M���<��׼r=�d��<g����U<�j�<��='(c����I�G=(=G�`:�\p�kN�<�:=���<�!=�έ�%<��&����;Q����A����m<���;�]=Xw7����<��=�ȕ�����n���T�뻕Y=�?L=��=�ѻ/UU�$�I=LW�%�7<��A�����Bs�Q×�YP=H���"p�< u��ys=<v� �W���'漫̽<��b�ʦ+=�5�;nW�<aY������n�\�M��.�<�X,=U��=��D��?=m�^��S��H,���n��=�5=��L=���<�=���:->��ϧ�<W���?=	�����>��O<Ӏ,=�7Q=���;�H�<�=�=�a'����<5�z=��U���[<(5�<n)Ӽε���<\(Y�%YԼ�	���6�<f<¼p5#=oب�������<.h%=�[O=wK�;�J�6sE�D�I�9[��/?������9X=�{�<���<x�*=D��;Gc=^[h=[�[��1.=V��</xv=B��85=�����\=��N���
�<5
<'�n�"�K�3'=ޮh;�[f�;"q�CK��M�>�|�=*���z�|�.9�X3��j;ʺN�B;k?��#=U<��t�H=�}:��|"<����9'=�ZE=5Sv=��9��& ����w0=��4<���6�N<y���)z=�a<ى:E�����ޔ����+�<�����<C�O���<'DE=�D��$Ke<:B��e�U��<��"li<v�=T�j�� >=5f�<�2��f�=�#1�ݹ"��!�\�*�X`�<FTL�.���/p����﻿>Q=C�}�y^^=dQҼ�7��	H=;�p�,Ϥ;�5�D�r���*�-�����һ%~8=��<J�]�L���_62�p.�<�zX��0�<�%H=�?=j7S�y�y=��N=���<�j�<�@���<�v*<.a=QUh�L�J=�u�r��<[":�&�H�ö�����<��;�v1���4�8�]<�o���<�:m����<5]j:��"��)�J�B=�6=�Լ�J:╀<�m4=�]J=�*
=Y$<$���]*=`wF=�#A=�r���B�M0X���;}}<@���D�7�#�I<Y5=�%�ñC=ӍJ=&�?�U~-<J���C�+������ b��v]�cS�=:|r=:�=�F=`+�<]�7=ĕ��z\=��?=.)H=�����<V�����<"[<��I�f�3�?�żq�����<�ٗ<�R=sE<�jR���g=;�=��m��b�$=�L< }�3���<�I���<@�R=.7���Ѕ;�`��X�,�(^m��q��&�Q�Z��~�0=m�8=�#�<�0���R=�A�}�7<�]'<��;\��<������<��(�|�ּ'�9�t� =��!=SQ ;�C��p��<��=��	�}ͼ��G=ޜ�ә^<�=��l=�~b���;h�O�>�_u�<�;t�Fc?<��=�/1���=B��;�����n���~Ǽ���<^ߤ;�xG�q[$;|�<(N��'=��8=�P��x���՛`=����+�@<<�˼IA�98�=�:��7=h�{<�*�=:�#��
�</�0��Z��tP���
=%#H=�R�t�=^ ;=q�>u<Y��*�������?���_�i��xw:a	9=��<7}����;z�=*�2�@��< /Q=�[ʻ\�v=�F;���Yq<���;�r��^#ռ�&=p��;�9�9[�5���Y<�1=�]���=+�=��%�
(�;�3�<'�G=��i=R=�<8�=*�l��<C�K=x+�����������!�Y��y�a��,^==�t[�A�
<��/��'=^�^<:=�.�{��<	�<o������(`=uW�<c�ȼ*ȼSך<���e �Ob=YG�;�l<��=Pf8��~B�`���Y���{=�p�;�y�<�����'�Z�3���Ay=,6�<+�?��z�;Zy</�x<w��#b�;���;o
;x���D�!��<�[�v�%�94G�2��<��j=HB����=>=��X=F=����V<z����r�<��?<�	6���0=X�;��o�{��<���˅=;'�=)��<y'}��Q	��Ne�,fS<�������*�#�����+�v�K�&���<��;�|,=�A$��.Y�k_�:�>�<����^~c<��<�Az=>{O:gY�<���;�)d��̉<�S�<�^����@���=د��jo�n�Y=h �<k�<�p� �^���s<���<)�<JټD�=�,ϼ�����G廥>��'��#��GE<6�����;�Ѽ��ݼ}��<'�2�#/=���<T�J�����,=`nD=z����e=`H�r	M��+=
<m=�Ժ�w=XIt��z�<�]$���ӼZL'��5ټu��� k*����;KY;<�S�}�R==�G�<מD=�e_=��)=��<</ؼ�7�|{�<�jE����<��K�JGP;JI�<Z�<��<���<&]���}�;�>�;�����P)=�/"��䍽�<� �<hd?=��vb�U_P=T�d=�(ؼ�=ǟ<��J�C�&<�9j<?a�-NL�S�������C=�+4=6U"�փ�B)�n1����t����d�<���7= �޼�W=��W;n[����˼�t/��N��I}&<Ʈ��}�=��=�R3<M�H�cA�wq�=�B<��<mix������h� ���ա���<8�<��+w	����<VI=�G=�F�^�m��ӻ�θ<�Th;Kg���n���"=bG=�r!��Ĝ����<^�;��<�����9����%�w�}<���1�$@=q(=\/<z����ߑ�<����z;u�
����;�<vl��
���<{�����=� -=����.=�؁��U<<<;K;nϼtgZ��U���e(��ɺw�P��;=�,<)U%<�)�op=>FG=�:=N$�<$W?��̃��������e=/6=rn�����b�����=-=@a�<o<\U<ƣN�~��
ü$���Z'<e��;��=X+�b6�:3��8,��F�<H�<R�D=��x���;Y��<���;�	�:�g���HE=60=G'��~=9=�=*�o<�p<�ky��=�<_H�;{�<=�H�v���׺�z�:qx��`�M��<�;�D���y���<ֹж�������<$za�	�	=�LW=1Cܻ����3ü��];x���G3�[���É=�`��),�xxc=��u�ce8�H 	��^�<N�����po;G�9?�w�(A7<�F�ɋ`��F�<�-=HM��3�"��xx=�����K�<N=�a�<
���;;=||V=��6��׼��>��N�<�{=N��<h�u���r=��C�=�;�]�E���O�<mL�<���]�=hd<)|����%��2��Nd=��<��s<� ���:�{r����=��$�Y?��XF=��<�#0����ł<�<��=Y�߼��I=C+c����:�н<�*���D=;��<�$3��F#<K��<��;u�3�� �����߂�q$u�w�=�;�<��������d2=�C��9��l?=9�<�Q='��m";=U=�e�<э�<˰<	��0�=<�G�5*�<>��;�Ǥ;ظ�JC���)@��I<�Մ�I�b���8=��;�~���P;�&\��&�,�H���x<l��<(E�<Crd��W=3$���'����;��?i��&��O�=3��u0=.3=ex�4�<L���*<�u<υ��ĕW=��;tV!<4�ż�Od����<a5=���9> =�M4=aWN�'mk�Ks�<_��1��Â�<
5����أ=�(^�<��+=ȅm� ��<�}Լ�4X<9.g:"HS; �^<�$=P�ӻ������h�V�;�jn�
�<�.=��<H����c�(�/�
;�� =[���Ҳ<��K=��<(����;=9�����=�+�� ���֯+=P���΀�<B�Q=�K�<O��:�w�0l~:m���y!C=AL�<���<��G=�>N����ǩ���ƻ�J}������:k�ּ�L�۠?�/�4��\����<z�漚=���A=�~�����8\;��"��G�Zwj<���<���<�E%;�o��.=� E=�֑�!A��i�<�kD=f�<J?�<��ݼ�(=��������P~<�Wh<�==�c�L���k&'���J����<��2=J���쩼i�R'��qf=>�=A�J����i�<Q����H����;�|��Y=�3<ʋ)�yH��d4<�g��_|#<��n��:Bg��S��;D�޼�Z>�mG=�E=p���o_�j3���:��Қ:ϘI��0����O=gm�ۿ����
�UԀ�63¼��<q`��"�S�����l�A�B�<��=��<�1��;=��B=Á��l�<"�;�==%(=ؘt=�<�%�{<��)=$�
=?_��y�=�d��/=/D��Ñ�<�=���������K�#����=�<�;�^����o7��/��˺=ۿ�;��/�L�#=7IB=�O+��,T�h2=7�=��Q=������<#ق=P�D�Ɣ�<ىU���N<ǆr���Z�6Q�<��;�$k�<�MW��f����������@���w��Z��Mk��A=h��<�ZQ�lK�!P�< �<�_B=*W�;���<�7�<n��3A<��)<z���Y@F= �l�� ��oR=X/V�|;"<<#8=��<sN�quY�C/���a���;��c=����n�L=�$��������	=���;,=���e=^v*<��� G6=u�>��S�Q���ZX=:�
=b9�9.�?�'-���3=�r����<�����K��hU ����;�`%<B�==\m3=*���������E�aO=&��<�g#�ϝ��n8=[��<��-�f�=S�v�==�����<�'=���<�{�;�n���D��S�<��<k��<�`�|u$=�^�<V�=D���ٺ`&��Ґ���żV_d�e��<Q��<�/��-a<������d<�9 ���<Tqe=E�<�z[=��A=J�f=����	��<̀��2���\�Ҽ#V#�_p=���<�(?����|��`R=]�R=a�4�2qU=C\�<���Ap[<.������z}��w��<��<��d��%~��X`���6�U�v��q�<�=Լ��`��T=�FA=3�)=�-�<�Օ;c̄�C*\=\��<�ꁼ�9=諠�z��@�_��5=��`��O���U<�� �N~6<��¼�c��_�=�=�<B/���U��Z
��0��+<�ւ��3�;��Z�D��;��:=�ԑ:tA�<�r�<��(�iG=�UN=G��=G�f={m�<-;����.=h#��5���a��Nih=F{���4a��hȻ��=���a.'�;$�A=�8i=|;�<��(=��<I$<bc���w=�J�;��N;��z=��i<�l�=3l�e\�<�e��;�U=�Z���1Ƽt6=�o��vC=\/���;c��8Q=�F\4=R��;�g�:�U&��~D<�hS=���<b�(=dX7�K$�H�=qG������҄���5:�T�<{�0=$�~;C>j=��$=P���M�=�3��_Y��<=�X=xC�结;�V���U���<sG��ӧ<w�a����;�P���'�F�<9���O�;B%���_��W=�=�e=?v伆p=#��;�E=PQ�S���2��Y��es3=F�E=�zV=yü��������Ƽ
��<��;Ȝ�=.��<�=!��<aZ�:����L�<��'�@X�A�ǻm��t'���a�K��<6a'�x99=>x
=˅�!�;�ibH��=�����P��
���k\~=f�4�0���v��<r6[=ٱ��*O��xI<�|=��Ӽ�==�=�{�<P<���� �%��s<rM=A����D�K�ļ��d�p���|�<�l�K�����p=`��F�����G~3=)��N��;�m�<�=h��<\�)X]=k75=Y�	=S�<s�W���F���<wU��?�8=�m�<cO���=w%˼�G�x�{�(�����<������r�b=?�>��dQ=<��p3 =˺y=m;7H=S��<�M�;(�=��"���= 2����X���6�3�;S3,�Æ<�}��9��;��<,��:gX=b1#=�+;��1S�:Ht	��ם�������<�[=�^�#w���t�[�r�ԴJ=��<Ln=|���ur��I�#iQ�xF<'d=
?=�μ)O�<KZx��7�<�*2=ѥ�<�/,=�{�N(H=�8:q�H<bX��h\�;,� ����<��ϼC��=�ü�ջU�<;5=~(��\����7-�V��=0==>��<X�<L�ּ�ɣ�܇���>$=+=��N��D���]�<�-g���ݼą0;��1=]�E=�-꼋���Ϗ��[r���p��C����<g�g��仦��>��;�.$�f{�<;/'��q=q.V<k�V=�`$=/c��*�żs�W����9fGO=�T=��������s�����.:�P><�U����Hm�d�0���><�U�<��;ڋ���'�<CD0����ü��W������<�?��fZ�<�!�<l����<�-�<��<�=�}�!���9���/�,t�Cj=�]r<��+��A=-�"�6�5= �!�T(�����s���B=V�ќm=�H�{<�� ���c�,=i�_�h��<��,=��=A?�<A_3��OF��4=;G�����7=5-�;��V�f��V�
=���;̗��Ma��H��<�?�;[����;����P�<9�;��A�%=�?� ��;���<�l<��l��<��6��*��@���"ż��E�&���j�=��D���
;g;s�3tf=͵�:�H:=��<o�[�6�V��݀�bF�s�7=�^����:;���;���<�����"=��=1�=�[@�h�<TY<������=j?,=�c�D�;�jzp��΂<�jJ=��2=��G�X�o=F�����;��K���;�u-�<��S=2gN=j� ��1���T�x�<m�<���<��*���� ��=���ջ'g.���{<�B3=��R�Tӧ;O�E<���"��<��/��J��-P���Z=�a�<96m=0#�<^�T�%�������<p�7=Y*
=��K�=�2���<���=�^�,&�<)Xr<fRT�w�Ƽ�2a==$�<���<�싻�;<���<x�=ٗ��)8���I=Ft�<h���BѼjR=�q�w� ��o6�J="�f����ݺ�,O=��b��c�<�8��|�n�$=���9M;n���͖�<�k=GlG�B�N��q=Ɠ��	��;��s�U��=5��<�P�9�t��L=�V�=![Y<z��;��T=�9�M�Q< ���p]�-�;=�YI���-������$�{�an0����<��H�J��<ڬV=�j��[�`=��>=՘�:ȒZ=�!=Et�<�<���\�^�=Y�"�&�=zE)�Jp=��\=�f,�F�=G���%f<W�o=��`<�<�' ��%�=��O=�?5��aм.�U<(�,=��&=�/���x��4H<���<�
);c����A�ltk�]��ޏ�;ge�<{˝<�V+=	�;���v�=H���+�;l���o�==�����=J=.Ý�ݐ�<_�'<�4K�!�D�>锸�7;�圻20��d����*�_C/���J'�А���HO=ex��w�?��O=J��Uw6�Pku��M�.��g�<.��߉��X�=��:��=�	��۬1��x!=��ؼ���<���<�ϕ;��j=����=7e]<&n�<���<�9���<DX=�!3�����
�<��O�X��0@��9�<�;0=��-=*J�<�F#=�{�=t �<g9R�b1|�G��<�;R=;%ȼ����e�-=^Վ��K��zA=|�<��P ;�c<=?�;�n�3m=/h�;�'�2#=m;����w/�<TU�;����K%9��"<C�3=�C>;�E�<��z=�F��n�:��<�Z���>�<Q�5=� �
gT=�����/���y=����s�8>v=� ںMA�;��N=93!�4e;��L���6��d��z�=5�I��b�<8;N����?�<��8���b<h�t���?!���M��S=ag=�z�<�gм��=�i=#	'=���J �;�i��5ἧ�=P��<�<S����	�( ��/�<���D>����t�^<��<!_K=��ż�q�zS�����y�{%k<�zn��+c�����G��4+=Y٠;W_ټQp='H�;`��;d�ɼI=��=t�/��^���=�o��<W�=�q<|�;�<�<�GF=�	@��24��+=�%�yP=>I%=bg�=x�<������K�RS�����<��<���;��Ƽ%�R=�)i��F�P�= ´<�=hV�<��л�=���$s=�4=ם�;��T=W���]�O=�3=f�;Vb��F���<�0=J��"�6���f<��=��<R�C�%F��qM��=y=�H���
=j��S�8��"�T�Ӽ��&��]q�ǳ�;KJZ=���<��==�WZ=T96=�)8=A����<���Ӯ�;�eԼ�����V���<=������s!�<��6=׆=BҼ�U�<ū�<NB=J��[@���(�<Oh]=fO=o����f��1;=	<X�=�Z�B<k=��Z��I���_=�$�< ��<d$=��ي��n�5q�i��;�m5�n<xU=*/=c�I=7-�B	��ӵ<�r�=.7J�$*=g3��װ<Am������@�<��;w�3��/��L�<ah�OJ;4�6����4��<�L���ZB<L��<D= ="=� �<pմ<�G�;� #��0�<��ٻ�;<���<�\Z�_��V张�d�E�q����<:p��M.��s�<�����)=���<T`?�j�6�g~�e�y��Z�	(�y�*��䳻.i=�_=�]C<3���@���=X	�<BӐ��Z�<��0�5�e�k���w��R=�U�5��!�&�w]8�H�s�����v�r�=r��<�vE<#!`<�����a��7���=±=�3�/�X=P�8=�>G��I�<XBc=i�;7r9=۳=G�<sc�<��<&NF=��=���(=�>=��Q��B=�g<r|�<��-��T�<i�M�#�p=ڕy�"ED���7=��8��Y=�5���C=�ͺ��A��Q��{6��������IO�s���!#{��|��c��6�<�P�<���^R��Ô;�z ��_=�ʸ<�~<=~^�<���<([?��)�|�B�z��<��:=�T���m��zT��
<9�.<e9˻k�伉˼<Ab=��9��O��S=��D=S�f��;pO�<܏q:zM ;���:O��=ɅM=7�»���<�柼����%�l=$8=g)=%=�-�;.k=�䙻.g �_L��|nZ�qj��U�������y��*�E;6�<~$�<��'��w�=^A<�;=dF����<�T�z4=�d�F��Z��8D=:H'<â���@g��л'�:�b�?o�;�щ<�({=�=�CI�~��).�;KD��7�KT���2���D�l#���:z�$=��4���z��N�ټio�<S$=`Z$;ΤD=?�g�'B<�TF���T=��3�lU�<��L����UO���X=�f=K=�lG�L-K<�ἅ8Q=p(=M?o�.Md=��<�6���� ���Y���K�=�$x��Eɼ�99�k��<?'/�@�|��'���U6�	�(=���	`Ҽ��=e���?b�gB=�'=	
<+����mV� �;Ι6=3=6��<�	u�׹b=�W6����<�=���Y=��<BL3������<&6<��c�3�<�ּ�ы<��<��7<I	&=�1x;���<�gk���	=��;��fD�MƠ<ې)<�=A��F�=t�9=숝� ����Lp:�Zټ��<k{4=�� ==l��'=����=B�;�<�����<�?F��\�;�w��&�	<Y��!��σ�gp�\fQ�9�M�7=0�;��(=�2q=.(�;V��<^��;�<���I�����F�T���L} �\=w�;_5=H�;J=�!�:B�#��Nh=Ehy�z�=��Z=>M-�9Ӕ�������9ꊻKw{���=��7�4>]�q�=J�O��q�;�6<j4>�rݼ�O���X����<�(^=2�m<��;�#���޼o ˼�iٻF���!#=d�s=��<=��������N��=�J�H�$<���<�`�;q�=�IF=0�F��c;<4$�� �N]̼y=�?=�<c3O<��!�G�z�=ϯ/=jw���=̼5S=*=�4��[
=A��Y�����J='�r��f)�ҼE= >�<��=�8E�����?)<�L$=�9n=�f=�U=�w;�32��ο����<�?�;��
��과��@=�����(c=�Ƿ�*�<(.�<���<�E\=��w��;�a���M�)=���<����5FG=k<��e����;�@��<;RT<���<�ˈ�o=�6�=������<�9�<_�;�0���{<�)=�\<� Q<b���\<\l��;��;AE�<C�(����<��5���ϼ������ ��h��[���<�:�Đ�ɽ?=(��4I�؉==�����d��Ӏ:P��;�<��2�_|�3��i�]=��r<<g�<V�&��q�ߑ=��5=h����?���<�̰<��T;�k�<���<�T]��N{<]���q�9�}^�~�¼	&=m�^��¼m^$=������.�1a=��t�/������<v��<���[r����=��=�r��3�D�q<Sd<Z����7wI=H�P�C�η=�ދ<(�(=�#�g�7<*�-<�o=��ļ�r�<�s=-s;��x<d��X��#���\d���#;�=�t1��=��5<kˍ<�V<�=?Rp��A=��>���T�����S�!����<gU��F=8�I�k�]=m�<։�!�.=��=Ȏ»�=�[	�Α$�S=�=������<�A`������!=%�6=���<�S����a��M��c]��yZ=��ӻ��8�H>\<��=<�ȼ?�O�>�j<pv�HK�;��==�Vh��W=�C=�q0=��K�ގb=�aҼ�e���U����<^O��n<=�jԼ�.�Ѵ���Q=��X=�Ms����<(=p��<�W����<������=��L���b���\��<?U=%�H�=&�/��E�<
�|�V���=�,=�R=�����9=) #=I5=TY���=��=t=�<= ���ݘ��,
��_׼d
�<{5��"@�;��h��=si]=L"`<'\�������;�ŕ�ɚ�����R��'+p�;`L��`��vx�n�F��s��Ã<�)6��o�<�*�jb�΃;�?�<�ZJ<iF=�܎<`�Q�P�K=ǥm��8��K.��"��D��<�(�<�z���W=�%F���=���Q(��2>; �߼�O�;�UI=��N�"�;=��%=�x��Y��^g��X�=A�q=Z��<R�b��B6���ڻ��D=�,�={ �=��d���$;���;=�]=��F�j<�*c���qb=�0R=��~;�f(��2=0[<�= x�=�v=z��<{b��C�;��%9�<G�=B��<��<�m�<��;��!=T��<ϡ2=8�C=��u=�Ǘ;�+��s)μ3��<Sr��f�<�?<Ȉ\=ʤ���n=�
h��V����豺�(_����/fT���<BzQ�⻅<���;Θg=�e��Q!=����ƞ�����S6:[1���r=Jx�����<.�;t�D�|-E=��;�/Ҽ��;�}<��=o�<{<o佻�K��=R���<�����A<�0b="-?�vE�f��<+�ʨ;��Qh������A�Ħ=�*X��ᴼ��=��
=[1��5=a��;rߠ��
�_�*��'ļ�����λ?�8��ۻ'�d��V�:�4��߼��$���<W�=[���ؿ�<֞h<s��<oA���;�� ����B���_�;+�d��L�<���:O�:T1z=&���u3��}=D�{��7=�"=u�˼�]w��n=��X�E��ƽ�F�;������ ��\��輋�U<��H=ƳZ<�x<�����M���ћ�<o�3=l������+�m�:=�I��X���C���>�h�o:����h;S=�s=�8(=�Ay��A�;��7=wS=(3<Q�k��<
6����3=va������g
k���&<~Qf;�K�<�`�<�i.�l{��K��T=<\+=C�=�*=%<=�o⻈����.��_�;|��;�7�;5-`��Դ<A�;=)h=���9�q;=�=�y�r@�<%cs=��<���=[
���ℽ^� =�yS==B!=��b����^�y.J=�\��
3��6�<y��,;=6P�=���<��3=����W
z�����S!<�a	<�d <�ee=��;)ԛ���f<�V��}�<o5<J�T��ps=�(4=Վ=�j4=��T�<�<�|	=O��<��\<�:������ou<=��<�T��D����<��s=��I��G����C����<�2ڼ�ϼ�b=~���4��<u�2=������1GC��I�<Hj_=��O=��!�5��9�E=q<��=��<��<�bl�EP�;չ,�npr��3=�R9=d�=L �SGĹ�X�I^��"jz��!�<~|=�1˼�k���?�(!�<��<�Di=�/t�g�<�6%=�3��Һ<�t<��H�_b�g�^=%�r�ˇ���iμJ}=�'�<q�C=Ty�2�=�@p�]?F=��= ���zy�;��l�A>=�S6=�����g4=��=��m�D�`会]P�B��
<��渔�1����p�m=�#=�׺<��b;k�=�d�<���;�{�<�A�2��<@m�<���<?Ph����-�<�L�;^�<ȤR=��M�ƨ�vb�;�ֽ<��7���)=�؀�@8߼�%< �*�3=#$<�<=�d�;ށ�!�<A�ﻻ�e=c
=��<7��LRY;H ���=�<q��T��<&_-����=��ݼh�<���;���<Ӎ�<N:��<�#~��9�<�;j<�|J<����{��jx�Gy��q'���F�<���;�@�̳Ի���^pg=�
1�8X���<��(<��<c�,�³�<���<Z=>�w<������``!��R>;��<6P��ּ��I�Y�<����}��#���=i��}54=v��:��<��/=8)�<���<"��M��n<7�%=DUD=v���(1���I=��4���<�S�(Ǽ����*=�xl��9d���2=��L=�M6=B9��l����|��*=�0k==5἗6���}����� ���Kc�.2<G%�<��Ƽ�p><��%�?�#����^&�<j�<����:uT�nW�����=5��i��<Mv4�^��i��<�z#=�6�`!��C��åD�(�eb�<q��
=�<��%=�"��aj~�g�>=]#,��p;w��;8Y����0w=w��;~5���n�<Ȁ���;wu<�U����<pI#=dm�<�=��	KX���@=@'���V�=�6���h�F�9<��f=����a@���=�-g=��	=����p�*��e�:���i~�=�/R�U���]�֚<GB;X1b�a����)&���S�ZB���>q�.� =7|�<b����+��o��<�<_�?�<Mz��`������F���6�8�;��)�<�<�O)��f�<�M�
o�;Ѭ�9��i�=�pX�� =D�:;�Y̻�+��eKM<��:{E4�{θ�0�%=T�5<�%=��[<�^.;L�c��~=/V��8�W=s=�#;V����;�u=?��ʣ4��g����FF�;�8��Vn���<��<�9��Rػ!�s=-f���M��Qq��S�S�1��="��:�1���Q?=B7�<��F=��<%��<)C9=C�\���c��t:<F�2��mw;'˻6邼��w=(q2=&Q=�,=�(�w�+��/�j�ż7�<��Dc�E��S9�<7?=�b4�W�����=7x�;�-��PV=&yG��7.=4�<�I��#b<u���l�`=[���ۊ��@����<%�=�]�<Ø���=���<��<�+��/���C=$o�mj/���Z=3u�����0�y=TJ=��5�B��;�M��vq{=��M�G��X!��z=��v�gE��ߊ��hռ~�v�^��<r��<��=c0<)�</�>=\��)i����̻�Z=�`=zә��o"��_<�S�����=eB����A=�WI=[��95'=
�<5��<��@<TE]�Yǿ;]b����9=�W#=�ɼ�x��ŧ�k,�E�<ȥ-<��=���;N�м�!���O�@H`�NJ��_��<R�<��<��P��[���Z=��<VF,���B=7 '=��q<���E�m\1=1�Q����;�F=fn�<b3��@�9Q�|����~M�~X8�?ӿ�b/���j=�򙺗��<%�d���S;[�$=���Q<5��;���<[,<���l�<�^�;��������<��L�bs��߮�;�z��*���n�2<��!�?�S=��)��Ǟ��c��=�����ѻ�Y�Z*�;�PZ<A�G�����~�E='�� ?1=^R�:��,<���J赻o�7���2=˓輑�^=z�a��T7�Π�;ں=q.鼜�������?�ao����:=Ժ���x=�Y=o��ܽ=��H=�m^��d�����8df<}"=��L=8��<�4�<O�(�[�rZ���l=.�1�Эk�*���꼓.���4����<�'<��<iȞ<g�[����6)���<׬(��==�F={4��Q�=�#�<��B�J=P^�<5>	�u���\�<� �<񇃼��G�hм��6=;8q=�˓<u$=�<�<����z&�ȼ#��;��b��8��:<�@�-z=�{+=���;b�%<K	<�׻WP<�W�*C�;�R8��n�<R��:�;4�{�}�@=3�<=)�����<�*=gT���=MI�:��\���Ƽ់7r�<�;fޤ9��<����m�h[T�a �<r}��B�;�F=h��s�V=�/=�Č�[*g<O�<�'��)�=Z�C=�k� �z="s�O{;H�<:�L=�gA=��:��=o=]�#��<�C�<a8�[�A=c�E�X2�d����Ȃ��e˼��<Po<�Z�<��<;=�7<���<�	���+9=2��<'��������;�v�=���<�H`=+�,���'�0�*=��/=e��;���ޡ\��{�0�+������^�����<�C�<��=�L�Jq�T�R=9aJ��l*�Odz=��㼇~���=��'<�V�<�=3B%= o������8=+�#���J=�!�1ª<��ټ{��_0�qF�<͹�<:�#=�5=ն����6=�g�;	�=��L=；��@�)��7=w�X�Qip��.���w���u=�VK�pI�OR=[tf�?g����=�v=�i<��"=}��Mm<6�R<�X��{����Ƽ�<�\�X=Z����E<r_�����=^��HU;=��0=P|����<C�H��$=+��<kF+��(��=��<���ʊ=����<����n������==�!�<t7r=���:��;M�1=��
���Z;���F�=�#c2�X=�u��h�태�~��[���e�X=P}n=�J��;�=@�?�M�<�f�<~��<�M�<�g\��)׼�[��gvƼ^y'=8�.�ǋ������ -�Z��$�?��=m% =�=T���<� �<b{=!�7����;ˋb<)}��a༿�漣�O=Qļ��;감<��ȼ-,/��������<�!=S�J����P�=���<(�E�%:7�b��x�<�2=�C�ʹN=RKw�:u�<���<yK=��ܼ o;�MG=ع~�]�n<}�����G��y=f�V=��߼֡�+�]���<=�Tt�ɓ��u�8;_�=&^�J��<��#�H=;�"=U�%�1���;8C���#�x)�g��<� *��~$�胼�>4�Qm���:3�:q�<̠+<�<f=m��<�Ѽ��+��������2��P����<I�������92=������3(��S���&�<������=wN뼲W�č)=>�<�ʼ�C]�c�k:�3= �
����LT=?� =6猼��b�G=7Q�ʷ߼��h�0K�"�G=�=z����;����\���=�7����I<�XF=��<]z<�<^ͼ���a�:[K��( �<n��<S�z;��@��≽���<��~=�K=��Y=ؼ�ɻ��gG=p�ʼ'K�;�q=�C#=F�(���<��<�<�bҼ��n<��<5�:���3=��<L��<s$:<;r
��)���r�<�q�;8�<��X�d�=2������=��R=��(���H=��μ��[�@�=.��n��P�Ѽ&h==�<H̀����<�T=2t�;��F�b��G�=��y��;�Q�:�%��9�k=�XI=�i<,�;�bҼ�U���%��/V��9\< �<�V�;4t�d��<�s����=|c�<���;��;�p�g�j=Q�=n�1��O���G��}^���<(�<��#=l�t��<�tŻy��<F:�NU���Y溃��<������;�����<_�<uYT=��B=�C�֗�N�������B<���L�B�S<	��됼�a���K�<75����S/U��=y�)�	Lb����;v� =�	J=�S��F4����GX<�ރ�xX�<�`�"+R��6r�i�Na��?�B�6�-����W¼��(=�dʼ9�=C=��\=U��<�Ϻ�i�Z�yE5���=�G�<�����~.<��ǖ�<�'$=�>�<JU��'�����<��K=�M=Ү6�A���
�V<ɔO=�c���<#--��r�v���I7�<��_�<~��!�<! �6/��9e����<LQ�_�&�j�<�v"=��~�<���9jZ��Ά��z6��Y �������B��V�<�U=xd�/*p=s�=�uD< �3jɼ�o����\=iǟ��1D����;�=�o:��=O�঍�dF��
.�-S�;�[-�k'�<(z�U���~��ż��ɼ�<=�iʹ;�8�9=�`�;m�I��Ų<h�
=8���L���Z�&�ռ4c��U�;�=⋠��e�ԍ	<�C�{�A�S<=.�J<��G�\�X<t��d��k �<krr=� =f�ɼ��m�L�F=Ѱ��,�:�>=�l�<�%�P<��{� :����V=�M�<_�/=���<��^=���X��|�X=F	=��"=e �<P5=ʓ2=LQ�Ic��e+���<<�o!=P(=��:C?=��Q=Usg�U�<_9�Cf =�:�q�﹆<J"\��3�<�1=�%<F`
=��:��B�؟�τK��*�<M�]��.=P�3V�<<[c�Y"�<������;�(�����BM�� #=m�O�|�O=.3A�M*<�?`�;t�<|;W=kb���<X�.���K=�Xg���A��1ݺ3�b�N=�jX=a�6�$w-=t]�W�\;Uܼ3Km�h�hɑ���=2�t����L�<�Ys��D�<h�;ڦݼnH��&��Xm`<	�'��{�<v��<�YD=�*=kG =Wp@< /7=��<wgB�M�|<��<�.�:;(�=�"f�f��<EY=��g���<�c=9)���!�:򾡼n�{=a�<�EP<y��gb=�`����n�&�	=�tn��(���8=����<����A��:��<��,��hܼFx3��un����<��(��M��ʭ�X&��������c�-=5�	��[3�T�'�|V�.$_���ϼbc�o� ��]h�qe&�;��;v&=�y�<�}<Ƣ�<���L⺋5 ��|�Z�(�lɅ=A�N;�i��&=&ϼ>Q�b\������8\���:.6<�+�<Vw����<B\P=&��<����y;�="��������<<7M�ł�:�]�:@!�z.<�e8<��;�6G�w�j=�&��"5=�*`<�4'���Ի�Jm=���:�&�<�}=��m�rq����=h�����;��J�#s��A�=D���Oܼ�6��	=� �<s�]�U�=*A�>RM��5W=�j߼���<�z/;G;
=a6��ꧼvv:=Ä�;l�?=���<*Fͼ�:M=��]<������׼#ҩ;�uQ9�A�<�,	<���;ͬǻ.����;V*=<��-�7=��[<�<-=kxD�q<jH���J�)vB==�������1=��Js�<��5=�\1=�T=v��=�<����;jϼY����u���AY��X=_�<��G=���d�:�|t���t�<oU���^���C��= �|:�˃<���<en9�gsn����<f����X&�pj-���==�Zk=7����<L�h��lݾ������1��Y���kp<\�,=ӄ����5�x�S�9H3����<��Y=" )����<�$�м��:��U�)�޼}�\<�)G��Qϼ6�=yl(�5�;�災)p㼇�ȼ+[=B
�<�9��=���<q2��堼)���#g�H�{=��ܼ6L���0�^N�����<�X���C���E���=/��}$R����<�(��������ɼoЎ�xSY<�Y+�����Gǩ<M�H������Z�;��޻�⼕|���
�d�X��o�<��H������<=Ѽ�q=ݯ��B�<O�&;�)l�)��<�V�pQ�<���=F�<=m�3=T6�<���)�<�����'�:}����&I=�	S�w4���=˼��%���,����Q"="85��$��"M<iP��Ğ=ޕ=�-���=��䣻m�<�TW�o�;;U����=n3=W��;��H�S�d<'=�;��@=��C=s�)=(F�<huv;Q�,�H�*�i¹<�p��3NC=��h���]=� =xz(=V���8g��$���{s=i�i=#�_��XF��Η����<��ټd;�n:4<#�=-.��T����`I�<RAj��ʻ�J��.�l=
�I=j��5E��B���؝��h=�U��C=.gn��9��$�8�	��0&����<����C���C=����G��=kwN=̰�<{a�<��O�N�<s濼�Ŀ<�D���a���l�^=k,=Kh"=�u$=��w���<C�<g��<Po��F1=������=[4����X�䦌<��;=(5�<b�1=��9�S�E=��hd=(mD�6�:�[<��0=a>�3�2�L�мե<�^�<D�;g�K��#���#��I=gґ<�N6�_6�=o[�<`Q�:[[=�%�<�� =hmw��=�j-�S��=��
�,��:
I<�(T:�)c����<[���-!�"C�<��<)ՠ��AW=�K�;z֥<�3���<D &�\����<�ռ�ˑ��j�C�����f=Jw��?�3�[�;=���<�+=�g��e<<�T;�Y =BL<rX�<7Jr�����F���<�3<\�������^�l�5m��m`G=�g�;z0<$X/=��=Al0�C��R�5=�K=�s)=fi�<eW��=�<|~�<̀��>��E�=�I�<O�-��� =�F�<��<��W���<� ��Z<�	`��z[��	=���#�?���=)����<��=oC=M�<Aו<�r�<���<��k��ef=�-�<��2=-�?=�
i�,5�#*�<6f`=�:�;Y<�m<<� �J��9�V�0M>��ң<ޡ+=���<�0�<0`�i�]=��;i,�]���=�=A6��n?:� �}-�<�W���@=
Ww��Ǽ_���o/}��)ۼg�:��<�[=D;��� =�!�,+�<�V<����)�{<�H�;>'G=��缵:�<�w�ᦇ��
ռ�f��G�:����@]��~<�M��M=_X�g��|��<T�F=i��PN=��-=Z?�<��:=��B�-.k=cu=Kϼ��R��(=��lL="��̋<�޼�9�z��O�(���?����Y0A���<c�7='�<�Q"�qJ8��Tż�U	���:���;��;���<�;=�.<=Ʉb����<ԙ���)�^*���������\h=��=ms8�b�u�N9�6 0�<��V<O��D�<�>���Y�*��O��9ݍN=�yG���:�����D5=��=;g��O[W=y$:��vB���J�%������$ʻ�k�� ���-,g<Ws0=���<E̼�x<z�f�=�I���t<-ݏ<�%�֨p=��K��B�� �<7�H=zW<��'<��<W�=0�=��<��<>P����<v=�$�v`�<�DO�)�J=0�<q?l�'?�f ༌��<{�=��I�_�lh�=.��xw��g�ȃ���ϼg�2��߼��<!2��Hv�I�4=�V2�,:L=�l={�<�w=wȆ;﮶<�T	�;%�t=�ad��ř<��Z���G=�;ir=�w}�[���l��<v�Һ~n%<Ҩ<=k^�*��<���==�^��>߼4�f��|���5=o�����=
Z1=��<<K�;�{���{���ڂ�0��<�,�g�"���OB$=tBM���;�Q�F�_=r�7z��=c1���wT���#�Θ�<HH=�E<;�T;MfF=;�=��<����M ��~��PV��s����4�v!�<:+��@ȼt���<i<�X:=��!����[=ao-�*d~���'��o�<̅*�kR=k?�T������.=��]<�,�~���Ԓ;��N�P����O=�Z�o�X;2�-��<�<�������-�<ho=�S�;(���un<=(w��w����<��<��+=h_��S�;��Q=��<���s�ѭ�<G7����X=�P�7�Sֻ;3=�I����b=l�j��<KL�<���K���	��<���<#�F=s��O��ײG�Xn����G�$R=Ψ�`�5�HȘ=m	_=�~4=�|��a��Q,=E�%���C�%H���Ǽ�re=,�:=I����D=�3��?U���׼�*ü&Xл?�U=��=��;�;S��¼��=�%={�Y=�y�<;��9��#:3�=�"�Ns���<4ξ;�`=,-=�9i�'��,hS<�i�������%L��2iP�8R<h�O���0� }���]L=�D���T��[�=���=�i�q��;ѧd�b��<��k��P�<L�=��r�@?ܻ@�<��V��. �T�<�*&�W�E���%��f��'$�������K=*�V��˻�<�zB�j�<�^���	��� ��=�WQ�,�d����<��8=��
=[q=I=DAN=G	W=�<����L�����[:J&F=c�L<���{˘<A_�E�*�'l��˼z<	�<XZ==^��=豢�<$=�����p�<��Q���6�%:=�nK���p=xݰ���7�m,=k�2��&=�M<1�P���<0�O:��n=Dt�<�<�^/=*"���=BG =�l=���<S��;�{��	�1=a!6�J�+=�̈́<e+,;�j/��o���lD=���<huE=>>=����!���a=wO�����N�=��<X�i�/L�<_N#��g�<�T�<Z8<A�<dP=!I<�� ����;�qH=��<�-=��7=�Nz<�vм]� ���<���<!�>�=����B=
��������]�t�,=F0E<�s�<zU/=�#�<ġ�<Ȝ�;��|�I��<�h��Ѝ�ɇ���k���伿4�=�ñ�� ߻)A�oZW�1φ�A��	�^���ϻ��0�K}5<ڢ|�m<EH=��ݼ�i��q<�:غ��I=��;�����6���ܼg�<�0)��=�<���5<���5�;��*<i8�<�n�a�=E,�,PA:q{'��ӱ�1�-�\�<�R=\��<����) P��{T;�M<�_#�];P\�����y�<��������b�<�{ =�z=�X$=*_b=�[O���K��"=տE��ui=� ���td����<M��5��]���T=1m�<e�[��FZ���=�a��v�	=�X%=��<4�q<�2���a�;�l�<�s�6=�Ls���<ϩ=����	�s<�a?�81z���/9%��=��
=SӇ�Xb�gh`�*�D�D܄��� =&~=l�'��f���ӌ<�����J=�3�<�bἔ��J�=��%8-�iBV���^� �9�t}(�0/=�S�4�\=G[l<@*��������^��<��`���#<0�#��H�<�,b=��S�᡹;olQ�{���1�5;�"=�,�<��B�')�n�3�e��<������;.=jt=�M=VZ�OG ��<S�`hݼ9C�*�=�=���<=�<o��a�ͼmcX���ɼ�
y��"��Z�=HY��f<���؉<΍�<J��N���u���;�K'��:��<�<b*�;	:���D�<ۿf=��;�H^=?���$����;ek�;d'�<&e��}�z��; s��(�yY�ລ<�6n�<�H.��Q�Q}[��!;T_(����<6==}�8<?+�;O��<���M����<�
�w���x%-=�c�<0��;G��<p�Z=t�J<�/��zϼd���k<�V@��,s<)�C=U�_;�?<���<�u<�;ѭK��a��j%�<ܐ�v�Z<�x=a�<����9;�h���W��1�89I�uj7==M=!��;�� O��$=��s<�2���"���;�	^�y��<G"�<�^	��Ն=� C=
��<�Ҽ�Za�Itk�bqP=
�T��<C���=�x�<(AE��X�T��p2�<E֮�q7���]'=�H=�r�5U=,�u=�>����������=j@�9+��wi���e"�� V��aK=�鞼��<�i��;->=.�t�7I�<*�f�('g�{h(��#q=4ދ=��2=&vڻ_�I�R;\��Mm=y	ټ
7=��?=4��<�F\=1�n=��`:�9�<~-o=ۤ>:� �;�%;LC;�f����<|� =^`�<2������>tu<�;��=u8w=��4���D=��=�ؼ@_)=���J=��s���<���<��,<��e< ����<N� �r���e
��(���e��2��s�<(RZ�FP%�&�pM=�SB<�_-=H�A�R���F�<�
E<��a=ɠؼ�<h��Z��p-���]=��=m���M�;<:�I=��=j�=��<)�$�lZW=	z=ߤ�����<-�
�pt�<�㵼�Vv��JI=o	�:����Z�w<gA?;�e`=����7j���,=;V��R�b��.=��<�0�=\86�s(����	��Ԇ=��ʼU���$CD�􊁽[*�.� i�<E�!���
�M�<��Ҽ�=�ce<�m���P=l#�a�o����<eN���L-�G�R<�,�1,�<zD�< 
e<J/=R��|�C��=]�p<ay��4�<�����ۼ�ܼ�":����<����|;V=/�CV��P�*�e�'�f�L�xL�<�j�<��}�c^U=9k�[9=Y4=���� =oF=+�C;�~<����:
b%=
�.=̌�<X��<�ٍ�^�K<�l����<���j���� =�pk��x�#D�<]�=�n�<%��<�]E�>�ټ��N�%������7Q�<�Ό<_<�W<��=��<��2���=��:U�<R�=���&�1�6�O;��2�+#6�9?��>�<B�v�`�`=~\Լ��=��?����7D�q��ͫ��c�K��<��>��iǼ/�q���[�����=<��1�l׼&���$�G��=��m=[�a�0ʱ��<~��U�<ĻL���<:ݿ<�H7�'C�;u�K��D=X\K��κ�~n =�1��c�pa<�x�ɜ]<�uu=IA�<�lR<�"�0XZ<.�;:3���G����K�����<��,�f=w9��cT=��F<3��<4Ъ<�E��j)���Gk=D�<(f=�|q=�q3����<y"<t����=�W8�*<8���;�/=��e̼�+�<d���C='P�<��A�Ԙ#���,=��%=�O�;Y�?��m8=(y�[��<�钻��J<��_����b&��P��<��</I��u&C��G0��i58�<7U��q�;2�뼄�Y��!�;��ѻD�=��;=�#����%���E:MPg�?�<�2��q�C=�ꢼkt�2�*N=cR�;��<q�=��-=E^#=��<��=�
�=if�M>:={��h\һ~���/1=l+=�TE��&j��i*��*|�u�B��4f=J�]=Ű;n&�<7s*����<�Q2=�;�y�</s;����W����X<����审<22�\�<��P= �<��<�;{=u���a��Ea=k���)�Q=�>=�����ӹk⼴���Y=������;�5��߻łV��*!=�R�<,��<��Ҽm=�;�=R����ɹ�g�B�ټ�z�<և@��v�<�G�<;ގ�/=��＾��<%[\=�R��O^���7��I�=4�<-Ft=nE�4l<�'Z;E#)�����y�[����`���"�<�޳�;�)˻y��<��9N_=���;�/�T�U��_���2���)=��y�8];-�0=��F��0�9��,=�����̦��z=p _=�Ӽ �\��05=$�ȲO��Bs=��9=j�:=HS��
=�d3��9��=A�<̿A;��<�b&=���;�F�<�Sw�� =f�%��c��J$w=�DU���ռK�K�[���J�><��</0���C=O�=/��<��<�>�<+�g<�r=��H%=}�:<�u)=H��=a��*�<5��<d<$��;=�*�d�����I�i����<<�Ƽ��=�u�<��4��L���<���;ן��Ov�d�C�k�3��E=�X��t*=��T����5�*=�d!=}/�;ٟ)<h�_�Qv�<΁k�N�x=�C<k�˼NN1��ޛ;8�]�)T�<$�P;�=��u�3<l�<�0Q=g���#ꩻ�D�w�ιS%<Xp�U:�R�tD;��;��ۼ��.=3⮼�V=u=r��<+-4�����Q(���ʼ�����u=e2=�`�gOa�|�1<D=�={
K�N��<(��:�@��-�=`aɼ�<�A�8<]�#=�=��(6=��=���S�5jy��؂;)�<(r2=]ͺ�?��&�C�%�>/�<�7?�F��<���<5=�o��=�t����<�ݙ<|O�=��Q�L�=~U��������]��;�._<v���� &9�'&�M�̼$<=� [�ߝԼ�詼b�=�w'=�f7=�Լ�6;)k��Jc;=ޑ�<\��<ϳ\=vx@�N�n=�t�1��UV�(&#�g�=G��<���)<����9������<�P���
.���2<�YZ;��*=7�O����<z�[=e�<�>�<l��<B�=bo�<$�j<�F=����9=�_�a�	=��<�Vy=��q=6qJ;[�X��8���T=;�<"c�;oGn��7Z=�V=&>�:��V=���B�=�琼��)��=��d=3k=5����E�׿Z���5=�N�y0=>@<>l���ɕ�[�<�k�=oT"�kO�<��0�6BE=��L=���<zY�K
4�I�=A��$�7��\�9��Ix��	��<����˖i�p�b��QF�QF�n%���`<E�ж��A�<�4�9F��=��`��ƈ<Y��<�*<1=�\U��绖�0��л���<�F=��������r<�B�<8=��/�yB=;YR<T�:�}Ἃ�u�ʐ�<�Y=?պ��J��EX�7�=��f=�=��<�b=!�ؼ`���u0��=Z!=+�����<�TB����<����#��D(<Tj�<-(/=���y�#��c�E�,�^;��<_~�IVt;mW2�g�"�X�A=`�S=n+=�0=�h0;z�"=F� ��C�p��V�jd0�"t�a�$���<HM��$�B=E�d�4;l�.�R��:`�.�>,;�qG=u,�]�3=NF���H =8�:�/��<��<�r���������O�<��-��f =�<bXi<�w�;�0;��;'ډ<����n���gJ=H~=X���n	�u��<��=�J=����] ܼ�=TYu��մ�p�=IWJ�蘎<#�Y�&�3����^�	��8G�����r�=6��<������@�W*o�t�=�3���<R'
=���:u0J��-�;H��<4�<[��`<j�=�N�<�u��b=���sl1��]M��F/=��a��g]<��=  �=�Qj�1�=��9=�>�=	>��'�<�@�k`�"�:�Q�K�Cs#������Ѽ��O=�f��[>弲[�=N��:�]=}�<���ex�;`N�<?��l��<�n>�Tf&����j�0��9ӁK=��@���;R�=P^⼮U�;��<3_=�<i�ļT��0K�<ш	<��;^�I=�/=�w*�)��<=H=�#<�!=�	l=UCC�%=�<,(��ۼ�vA��\�;�il��<g3=��<��=�{�6=��p�}�ټ6.%���-=�3�Vm���-=���<L�B<oI���3��a=���<�1��F�8�M=d�_<dne��#=������=ϖ�����l�O=�=C�U:�W���
=�@;;�����;р��Ɂ�)鴼C4�� �=�젼/`<�f:=:7C=p�׼�1�;�-\=��<�u=�}V��Ե =�`=�6��^�<�{�<�I=�����=��v�yN���:�ĵn�(>�V'=z^n�/B������6q<#F|<�F-<(�O=��=�l�����<�R<��׼�#=���<���;�����fp<��9������*;��ͼ������FY|<Nmɼ�I���P�j��<s�)=��ʼ�3<�2�;�D=�j=e^����~1�<�gD��(=�d?=��<�c�7~N�x�<��=(�ؼK�x�fƼ�9$�p=FWQ�I�=i�0�h�5;2J2��=����%�V'=WH��/<���nT�G�b=���<(�p=�ը�Է#���S<$W;��=x	=[��<���;xu�AO�<(M�<�7e=�T\<��=�Q�<x��<�+~�犻�N�<�#���W�<�<�d!��aX;V����<ɐ6�����)�<7RM�~sȼiҪ<ZK��a
�;S�='�<7�=Ż+=��=W�:<��μD�[���"����r=�����I+����Ù<��%�\�ϼ�)�,�B���<��<�����
��!�[T�;�:��d0�<$��� ,�<�}<��<�K=��<*)=���;������D�>&����z<��6�?@�=�k,<?�7��o�<��4=��.;I�3�:���f���(�>���ͼ �<��?<�ۻNR=�GԻp�F=j�-�2=�_<:~�����<�c.�)�=�I�<E��� T���޼�z�����=����΅"=�3�;oj~���O�m�=�8���qf={�_<����b*�;��%�G=P���.=�?N���U<�4N���`���"��r���V=H <��;?G��N�s�8=�r2<�K<��=P�=�6»� ���_T=l�=��<���:���mh,=}p;x�=������ �:���Ƽ��\��&I��W�=o��<~m=Y=D	�F�d��\=�Q�<(=�C=�=y8��^�<e)0=��c<�����h�f��B�=��4j�|�<򑀽��μd0=��/=�Id=pgC=B-������̅=+A3�!"=&*�=)f=��<�ּ0P���J�诤��Op�����<��}=ȑ;���3�~��9����<B�.��<�l9=1�r�G�ͼ𸅼��»�rn=�Q���;��<��z��T�:�o��-�=��=��D��U�;5�&�Z�R�;w=`��֚<?M��w�@��Є<ĉ�Yɲ�E���:(=f�7�*��AHS��ݍ;�*%��#ϼ���<�ۦ��2����<r�T=��g��wo��>=*��=
���LD;�ٶ<F@	��Ҽ8!*�;������<��6=�^�a�n=��,<���<K�7=���<�-=)JW=�O=�F;I��<C�U<�ĭ;nG�<%?�\�Z�b�9;=w�j�-��ǿ�'<�f�8�T<JO���"w��8=per�\��< �D=t�U=����=E?���oj=[(���$�;�N���=I<�����S�/�ܻ�g=^�O��E4=�م;K�!=��v��W�<%ǭ�X�<�ʁ=c��;Ib =��3��7�;��\�0�,=���F�'�'X	��U�<'d�<��<����/���v=�=p~8��2*=$���.=`\�r �<m�;���<TR;g6�<����_�<�iU���W<�>��__��m+��������8�w;�����$��#=��]K]�s�<�L^���=�¸�	~~�F�<��i�2��<�Ԓ��Z?�Q�=ʓ�<�j
8�S;��;����=,��^��<buZ�@��;�^r<�����=�2u��Bg<J}�;]�=S؉���i�����A��p :=�V�;��<�ֈ���I=h��<�%t�L3N=]`���=$J,�bI����<�Vp=�@���9�ɨe�
Ɲ:�S0=�s =�2=\)=�
��F�z>=4i<��=VHC�h)Լ_�g=޷=��c�鼡u�����ս;=k9�4��������c���ؼ��0;<\Y=!A$=r��S��;;=g<9�����A=��<3�&��e��GQ;�|$���L�Q{�< �!<�s <	h�	|<�(H<��<��<N=#�<���]=����Yg<�@O����=x�ﻞ����<#e�<�g<�����.<$�<Ksg�?=�-:�-5J=�^���=�.��B�<�(�<u��<F�����G���a=Y��;��=���<�{��<g�e=	��̷=���=��=W|x���<�4W=�懻��3==�<�g<��i<3B`<>��;�O����Z��d�<#���H�,��|=�]��G=�[Z��US�<�+4=J-�=w!g��  =#^v:b���'g
����<�'<�-�c�|��P�������c#�<&'��Z �L���_�D���,�=�����~�[O��(�0<=[�,=M���p��A����=w�׼9�=�<c=ZM��'A�� ��<�짼$����� -=��M;?�r=3T�V�r�NJZ=�d#�F�k�q\�<�`�meY��¯<K��S? <��<|�a;��3=ᗗ;k�'�\_�;;C�;��~�ﰀ��r�;y�\=5ְ�y���-=�gw�rSa���=�Ñ�<�<�y}�=;����:��<�|<=f���%
�3�h<���zc< ^���]�z�(=��~�qg�<�,=�T=��F=��,;e�<�5�<V���GV<���<|����
=#��:?i�<K�H=`��;ۖ��I�@=3���	>Ӽ�BQ=���;�6A���d=���<O
=�+ؼ?�6=�"�y�f=h�<�	�&=�=[U=,�=�=��=����B=Ѩ��鐘��6)�K�^=l�z<4޼o�8���E�}ʈ<� �i�C=��j�c&�;�d�<K��<�h�9�û/�=�.5G�Cq��d`��$gi��}�!=������m�L������:�`-���'=��
=���y7�S@���v<�=�L=K:��	y��=�"�;ݏ�c��<К�;x�6<��/��*�q'R=G���K<�b.
=j�����k���(=�V�<��=Æ=�:�<boS�%5Ｑ>'=.�<��	��'.=��;��5=@�|��QV<:���l��?��
=I
����<�1a<҄=�	��V`����l�8���l=�'����<�dF=���;��q�JXF�,�B�N>O�l�=�s�:Q\=�r��sz��nk=�9=܏���,/���H�&}=�x��`<��F��=�<3i�i��<���<[e�<cU=���q8�<]�$<���UG�@=�- �{u�<I�=`B����;^\=N)w=��<B��LI<�I��#V����c
O<v�6��`.�1���{3:��<� L=���<��ur=�J5�Ё?�+��<xEA�r��=`E=�_{�F��<�x�W�q�Ee <�@�H=�ч��oL��,�< �$=3dƼ���W=F�'<&�+��<�q����<�̀�g�X=��<	�=��$�����,+=y���=�;:��<6K��q��+= Z6�a�Q<��;y�t���J��d�S	������$�G�����*=o56���k�M�<����rWѼ6�'<��:�N��N��i���4���X=���<�_<�'@=��/�Ϊ��S�Y���n�2W��	)��X&�0�8=���f���k��q�<u
=ѽ�qX�<�/:<����L�o;�i	��=�B^=T�&<k�x<�Q�
ն;�0�ߤ3=����,�;<uz=��@���T���<��$��_���Q=bJ5�_�$=_V
�j��f����^���]=������@=�+��(P�B������tq��<�V�
�s�|=�eQ����<����m=b��;��{=������#�%m=%<�C9���=��=�2�����<�@p�)`C=n��<�㕼eMY���@��+��k�;��=2�}<�G��S);�
�<gż�gJ=]B@���/=�_=U�<�B���Ի�T�<�Z׼�:=��,=�d=�=�����=�Hj�;�<��=N�1=��v<��%�ʼ��H;��;Pż+N:�\����<yy�<&*Y�1�}��T���U��ѻ�;g��+���<�C�;��= U.=�w<*q�;���<�����V=C��;@f�~�Y:�j��na��T��|�R�(�D=9�<<3Z��O��~��L$=D	]<��; Hv�=�*;iR�<قG��/��y��<y_=� ���( <���<=���0�-=ql�<�Z#9�'��?+�<��NQa=��<�'8�P	���4�>S�<�����c=QFѼ/UE=���<u�Z��_�p�G��'�<==��c<�|>=��*=�F"���b=vv<�=�V�1�K=�M@=�:h=���<���圁;q�g=z�9Ȧ��I=-Ƽ����S�����U��;�f�<��=��˼��?���#�=�L�<a�]=�����v���:�W�<҅
<�1�16)�07G=˒'=��n<�I5=���kټ�B���㼺j�;4 ���s;+�ѰR���Z<H0�;��<�.r��-�=$�<{�:U~�<��=�=�<p�<��R�6�w=p�;��<�?»���Q���ko=���:��<| ���==~n=�@� p=�g��z=<=�f�Y�C�$�H=�>��\��̶��g5>=���<:"=��>�P���*�o�A%�;�',��؏��몼9O'���K��q=%!	=s��:>&Ӽ�v���y�<.�<_���j/=*F�_HF<�.=U-*=D�N=γU=JN<��<�3=S$=;��kS�μ|�i��#ɼ|gT�a����ٻ�F=�%����WT=��<^��&�M�Jd<Ew�J =�M<�(�=���X�<��:�(m=�����:=��<Bj����;L/���qH�Z۷69�=���v9�p�ϻVS=�Ԟ�l�<�x����<��Z��>=�$7�˘`<���<S�<�=�|/<�.�df<��#��b>=P9	=��+��$=�4�<N�m=-�=��N=<����<=� \=6���gz�;��?b��6-��;K��s��k��<�	�~�u=��n��;�<���<����弗n�<[�Լ/��<��˼�!�:]�f�9=��l<Ӻ�;��D�VU;l9�Չ��"T=��<�1=
�0=,��T���}<�����U	�~�3�9=o�W��z��<(�=����0̼�zT����4�3�ͼ�)='0�<;�g�<H-�ڙ�<�i=�J��Mn+�[@��"���]R�VTy�N]�<Z@�<�-=��=g�Q=S�<q�Q��4��>�@�R�;,�#<��O��q�<��Ҽg�s=�!���s):D��;�~0<R|��M??�����ٵ�<����<��<��<83�"�
��V�@9�<�˲<K�/���Z��~=Xh�<�cM<H E��A2=�0�<��<N�?���=@d?=��,�)�
�d�;`\���ƷM=����-����6<��3=������;�Ȼ���<r�/�<�廸%'=�W)�6O,<��q<�n=Tz�<�3i���<����莴<x�!��m��k�;K��=X�:���=tأ�3�;=��<ۯ�8;=���X�@��D��nT^�͌:��_0=߶�*����	�<�Y���> =��Ѽ���
��z)=#DF�R�м�&��6B=&��ڲ<��J�V���xK�9�ػ�ƪ�{�=6�i=�"=��)�@k�<	����Q��U��$=Q�Ъ8=\TE�bm�<��J<�4=�,h���J=���<����k�y���g<r��<5e3�fMH=�5�;#ͼs��<��
<�M��H
�(K#���.�p���c��n�=]Q�(�]<"��M�~=�++=W[<3D(���mG<I4�����O==��R���0<��-="g����ᖂ��'�Z����՞�u�ؼ%u�;6N-=�\k�	�=�`��^Ė<w����@�ڎ�<F�2=gj�
ɼ⭉;���<d�<� ������=�D=kgQ=+Ԗ;��0�F�=~O������'�g��;��X<H<��X<h�=D�=�>��s�S�3$�M�Ƽ��D=R��<b��9��=|��6#T�;���]�f���=�kX��]��;<�02��=S@�<{��;`%=��2
=��=8dM��k��*_=�
�<����F1��)����q,=y���p��q�B�z�1��M��n40����;x�Լ��ѺZ#��tzY�Zb-�A�d�=%t�����P�<P����R=Z�(��=��Ѽ^�:=Q�J�6�<o�^:��/=X�$�
}M=�j���0�S�8��
��μ̻=v����8�<��;U�3��98���6=�� <[V������<���:<���(���S��\��<�<�;������̼�y+=�KN=FV[<R�=��a�13��ۛv�\;D=qXF�#Z����r=�_}=���Z�X=��)��S�=�;d�G���]�J�7���<X���=��Fx���Q�+~ =%�8=_�<��=� B=%En���r=W��<;�=	=A�==o��Gv�<:%=?"�yR�c��<�7H����t��=�T���W4�K����<=��h=�0�<c|�� �r}ۼZ�\�J	���gl���=@Zd��� �#{��;l=^�<|�]�=Xe<%�#��EؼT�=�uh����9�t�?Ѻ;OZH�Γ���f<@��{�]���@:��=G %:� +��}=�K�~$6=�H$��fG��Mb<�S�󬘼3��;Д<��<��<�j��LV<��/=+9z=��g��"�=I^1;H8�<�P?���==rD=�==@<$=(IA=S�;��X�(mS�W��pU�<�&��Q���X�<�G�<�[�Ղ�j��<��<uX=��<�y1=���<�*߼�<�T0���K=���2(+<����8X=��=�K =���}����1�;$�<.��<ҿ^�����1�!;�� ��[=��４a'=�͠�/�`�V=�o;��CG�Ot����_���X��,���!=R5�<ϕS=x�t=<�ܼL���r��=���F�Y=6;��2=��u��-x=�U9��K��P�6=�,����j�� �B�� /;��h�����ȻF�<��U<�
@�-*"�~����<�Ċ���< rc���<��=}��A0���$���B=�O(=���C{;�7=`�'�*~.�޵��=<�9=m�V������	;=�1<�S�/7<� =���7�9<sq=O���+��<��<R7<<�W��=�ʝ��{�0=K=�6=����a�<��!=�F��v�CvC�}����$=�߼5��<!VX�y�`<�9=�lg�R=�Ļ��m=J��Q���#�<߮*�T	X<��E=�F���I��M�<c*=��-=���u1��i1=�,v���Q<^�6��]��|���==�M\=��=����X�x:=ն�7��;s��<�(�<�I=O-H�n�D=��޼4 Q�DC=t�<�)<=�
=ӛ'=S��Zb�+C��t�;��4ڼ*�=<�4�=�#7=�g�<_����,=��g=r�ɼ�i�<�w�:���ꚋ;��#=�ZK=��_�n�]�s��O?�]�=�{_<�\Ѽ�a =#� =��W=/�������0�⼻y�<��U�s�P�^K�R�$;W�&=���<��j<D�ƻ���@�*=�p��؃�� �<���<�u#==l��5)=�=�=2��G��<^<#=p��<\��<���=6='3H=�k��U�=�Z=�;<��<��1<�f=�Tݼy"�;�<v�8�(=�����K=�~�I� ���,=�xF=y�~��$��;P�/��f�-�=�D����<��<=�]�sY�<Ų�<x�[9�R����W<(���_b�<pU<�n�#»4@=I�D���^��8[<No�;K�k��t=� ?�<d�=�T�<��;5,�)�<��<��_��,=��Q<V��<��B��0���v=˅�=gU=F�;=)��� ���e7<))}�qa=2Y��2!ż�=����L��őe��iO�e�<�>;�خ���<�x=��%�Z�7=�Q==S�B��첼��*:a�r=�
�;Ћm=�T�KS&����k5=���L/�::)���c=��֛�<��A<�#��A��W'�<��ݼ�����#��`Z�P5�A�k8��Ǽ�B-=c���5��;":=��<��{�I�����@һ2�<�nT��e��]��l�0=�ʼ�������ռ'T%��F`=w�p=J�;������B��׻���<�7i�q/W��;��t�Q�;���ػ�x��]�<*^ ����^�<�J�p �"={�Y=�8�;�=�P����_���ür�=���kF=Y��9��=w��P#<#�<�[u=6�-=�y=��P=a�=�X =�=A�K�#�Q�[�}���;[��3�>=(O ;��|<�?~��μHS=b`-�m�R����]y#������	V[<�Nc�^-��;[�Vl�:�qμ1u%=�$<��E����;
U�<k~�<������<=Kح�n.�׬<mB��b_��ay=�WǼ|Q�Xļ����P>�
P�<�z<�+V�Hp�8_�^=�E����=���v�/��;� ���:��ߏ� mf�6��<_��<���<��R=���:1c.��F���c��i��Al=NO�/=��.��#~��#F����ąp=P�&���<7�7=�G��,F=�c/����U:A�*�5=��h�i=Ә<�^H=�.�C]=�e�<���(ב�9PI=��'���u�`m���e�:�6}�A�5/=lɊ<��V�R���'=�6`y<Y>X=���΋�;͞]=��˼ia=o������BŪ<�E���vz<�}d��/���<ȼ]e%=�hh��=.=�-=��;�FG<�������D_�uރ<;�@=�#�-��<�b�<x�f��$�����񁽿}D����4�?�V�l=3k.��)�<'��<�!��*�0�@<�.�<���<�k;��K=W����Z�<�Q=������ �����0�]�tm�C��<�/�<̡<��q���=�\����A[=��=���;%P༕�=�%E�ϙ=)4�<n8=�>��<@H�2�y=��Q<_�<�f=G�b=��;=��<qv�;�L="	=3�=���<2�*�3�=��<Ӯ+����<�#=;m��h-=�����=�E=�e=��</�˼�7�;�U	�z��<7	<�Az=M�=�Y9=��\<��;�.&�� 8�<�F~=�l���;�$ = [�<L�&=�S={�a=ڥX�E�F=_�;�}����O�O���޵;�R �;=66%����<�x5���7�Ʊ%��F$<U�X��$<a�:�hc��V��t�?=f�-�tF�<�A=C:�%�;bUM="�=�1=E�<��ϼ�>><��;�K��Z�=t���M��;�ެ<�i=�ނ=��G=&���<��=��k�?����rs�M��)�<��t���iH�<��0=�u'�p�<��3��/��@=x�P=� ��V�<�ΰ<�B��H�;%�=�Ѵ�)'��j������fҼ���u���<���]<�*��L=G��WrD;��i�)�I8)�kݍ<͡ɼ�wϼH�<��K��><P��<�м�B=����  7=g�<��<�K#�Y�(=�*'�<�P<�ʯ�]洼�&Z�ڮӼ��/:�~D;���<�~=���=�o9�)�=<3�;��o�w8K��"��ڻ�;m�g��<�L0=�L�1�<�2=�
=B�<ж�<J*=�F���O�\|�<X���U�<�l��FZ�� �<Ml����i<ǋ���No�IP��
=����d��@~<=�.�䇦<���v�����k(!=�ȃ<�`2��=�gj;�|�<�d����<3�g�O0��"�2D� �(=7�
=��.��$/<�=E��̀�1��<!`�*�8�~q0=.+;1�1�E����<��Q�P-ʼ'=.�;�PS=AH�<��*��%=+ <���<�*t���S<�[2�1b�X6=��h=��J��E=�b.�T�=�q</G6=�r����P�� ü�X��=��P=��)���D��8=�+Q=|9p=2�<����T-e�"=1��̼��I=Aq�<R�S�Wl���VQ<B�,=��%(�<#��nJ�<�x=Z�6�<�=�c=�
�=��P=��%g<���<Nn�<�˶<�n���=I0=r�X��R?<,򢼃��<�B߻�"�o�u=٭�=��9=��==��:�j���P�>=�ҙ;�HC=��/�?߼<�ۼ �$�U���L=���珥�b].=-N�,��<���<-���;=�#_��V=4�A;]�����8�Z<�^�ϫ�<+�n<J>E�j�Q��]��w�=_�$������;_�<�3V=��=��t�~;K�m�	��<�.<�1��:i=�Z*=mI=�!μZAc������e1�<��=�$�;A�T���<
�;=�g3<���>"=�+Ҽ�(>��-ɼ�}0=g �<�~]=ׇ�J�Z=ԯ�<p95<�I��	�"=���<�Y.=Wp�aI�<�5 �7��<=�<F=Eu=�� ��n����*=X�>=���<�h�<\�#=J)c=��<��<�/�U8<k�'=�:����8�ڜQ=�s����=��J=�'=tq�B�q<���<
��o!�bd�<u>��W���=���!J�<�t��;<=C�Ố�@��0:=�<v����镼ɬl��w���|�y���t��<9��b�:9�E��k�=����_&\�K�	=+2��7k�uj˼)B��U��62���B=�<`r<��8=:!G=Q��;#�==bL�=)=&��;��LjL��5��tB=��p�&Jb���c���ϼ�]�-	���켋cP==��1��O���=��j��2�����=lG=�s$�C#t<ݿm=���<Sp=,i��'=F�'<;`3=��^��ř�4\[<�7�?�f��<��Po�:�;�lC=���<ŋU=�0�<$gt<�<$ac�t ໯�Ѽ�7z�}�y���u�*�x���_���#�lY���<�?=���x<������E���R�*7v<�<�<G�k�#����6�]�<�;=F!]<!�Z=J��<ʬ,��Wd���[�)�{@޻%����
=��_�.�:��m�J�}J�<L>��9�c=ǣؼ �+�?S'��W=L�<���N�y�7���R=�g(�@������+-=�#�o �;�T�Gqi�ve�d�����4=!�_;X���Qw�<��;s�; P<^�<�hN��#�����ޢ2=}���S�:�j\�����I<����5n7�wt4=Et=��q�O<�.�;Ҭ<� <��=<�K��o4=��a_�ӣ�<��W����.=�����%ϼ��m���˻��&=:&Ƽ���<	]�<��O��7�<��S=l��<n��<$�<t�^E<,�U�:!%<Ðl<��"=���<�s���<x����=���<�t=A/'<����nؼ�W���_=�v<)~>=ٽj;�.=��;j�̼��������M=Y���Z-H�U? =iǔ<L=2�����Hf<�׼L����-���d;�&=��ͼ��=�μ�M��<=��<5���Һj=���<j�~v=�=�*������{�<V��|I�����B��"�W<S�I�����=n��:�=t�C=r<3E�������Q�<�ㅼ�+�<·3=�<��n=��L�*q���s�<_b=�GI<�?N�J�S�Z(�g��v���;b�9�^C�<��K�^��<�%���?t<��="1J=��6<<�`=-%=H�;��Z�'�?���,�MR=�k=ϔ�ؿe=��;��=�#�<;�G����!�ӱ �K�<�<͗�<���=�4�'���D/�(T�kn<��|<�=M5=���;�tET��#r���<��ؼH��=��;:�F<Ќ�;���F(���4�݌�<����n�<��`���#�)�:������?�/��8X��wY��!=Jk"<9t=G�='�<��߻ٿ���t*�,�M=��<;���[��\<Y<�9S��%����g&>='�D�_�5��q�K���\���w�#��<��
=0�j�l�"=�0=.ͼ+0=��<��}=��=�5=�c,��1/�?<8���+=�څ�[��i��;�8<��<ŅF<����u�6�MI>=��<,�W�UD�<�1E=�?����W�:9=@ӳ��=�>4��u�<Х�k�;�{W���i�p����L�F�Y=I4D=
<��-0���V�;��=fkU� Aϼhb���=�U\=��<%��<wK�/�J=/\��Q2�=�2��<,�޼0�;=�{=?{r="?���N�>�����9k�:��<���� &�J:+=
�7<{���p�=�k���A<ș��Wp:�a4��e��y+==v�<�I��� #=�rx=��_��X�;_6=���_�/1E=T�<8�1=B=T��;v1W=���:�����؏��'s.����; ;=���q�HX<��r���<B����=<�:~<�b=�� ;,�M#/�|�2=K�|;�=���PZ��7d�	/��&��<��Tּ�6=�ϻ�G�֮�;-Z=8=��K<2):J����׼G=�*<�W5����钭�`����k����<ʝ<�?3=��A9����F�/9=��D��-P�8,�<K�?�ٸ_�%�?㼵ʹ���#��>�<Qjn=�ͽ�O��E�޻�_�;�Q�\�<0!o��߄�Ǣ�<^��G
ؼ��Q=5D��f==RP�`=�t=�&o<&���y<{=~u�=,�*���&<9�;hs�n�n����#��L��O�q<�3������=�<�Q@=�wd=�9�R=���<ƥ<"g�<�ԼG<h6Z<o��0�	=r��<��?��`S�㣁='�1=��=<�M��a��8;����h<v)ۻf�<�g��)# ��6���N��a��;k�Q<Gt~���h<�|����]��J"����=1`�����߼s#=�a�;P0�+@O;��4::&=eߕ���A�ȸK=�7=H���'=Ÿ�<��8��k��`$�<@�=�1<��;k�����=�F<����3,@���<e��ҳ�<��<T���\�<��<�5.=):<���%=�a ��ڍ:�� =ob/�	s�<?���M�(=�@V�U�W�+΄<]���F��<P`���<Uk�����	�ۛT=�D�;�kϼ��%=N��;X�f<��s=/>m=����+=��[;t��Ѝ�;�E=�4Ҽ��&=��T=��<]W�E5����6���F=�G��h=�ܼ�#ܼ��ݼ���<�P�;J����E�Ƽn��$|�@�Q=�g�<�)�<9�K����q_��u�л8�6e��'���$=�nH�|B� ꍼ��2�ʪ7<'J�;O�=;��<ة=�i\��Jo�;4d=,& <N�9���%�¼��
=�2�\};=(\���<�{�:��=��<u�_<�#伜y��]M�7H�+�=<8��j���ޡ<�t�����Ә6=V#Z��b;wP�<ဂ��������U= �ּP�U���=���<��y<�߰<��ܻ��}��DǼ��Z=-M�hA=���;�߼Djq�!U���W���"��D��Α=#F=�B=�%b�簇�x �fs$=+�*=��<-+F<�Ĕ<�kl=Y��=����o!�+o޻�>&<s��<_�;��<&غ�� ����:��@�[Z=�[A�%-;��!�(=k�[=��ڼ�0��4C�����qg�<h�=g�<=(�M�^�Z�0O=o�.=|�+=F�)=�]�<��ۺ�T��7�<zI��:���;;n�<|�M�s��;��=�V�UtS���B�EF�<�:l�̰4<$�E�}q�bo��<1<{�"=������;߹���d<��U:�=�yN<�U��Fj��ܖ<���<�1��Ѫ<7�i�E|�<�؃<Q�5�N��<��e�<�C���+;���<�幼�K =��c=�H�9LD����������<�<xe����8=":=���<��g=$�����["ĻBI鼣տ<E=4�)�-��,4���H�;��f=CH��FKI���z,
="����Ca=�&;���w;^�=5��<6�����I='��;��g<,=}"ü� �:@U���ͻ'�!=Tθ���ݼ����(�:?�(VQ=�(<e&���<�Ǣ<��#�֐D<.���^����<�m4�#�U=b�=��I=l#�<�31��<��%��Y+��\�<Ǥ���6��Z��<FD���4��D�w<�}��n0��ʅ�9����<�%�/ <�Ǽ��a�<�$-=�Ł;�5�63�Z�K�p��;��|��S�s�w�[�F=�.�=�=;@�-Z�=�B<<�=	<�T�&�����<�iP=����żtn�F�=͎�<{�^��/�<�,=J�	��w�N�=�Կ��E��U^��W������S�}���W����&-=g�%=eD���=�3���0=.8�KJ���+<�W����߻��=3� _m<bD�<��k����<��D���櫟;�����^��;3�=(�'��3�U�V=DXW=��=��7=���/��=� ���=�v.��#���a�0P&<a�����B���ɜ<L�=@*�<N��<�]���k��wQH��vQ=|=���w��=C�,��/�<�蝻��F��	)=#�<n\��&�<���;��~=E:��c�<��X���G�O^�=���<e=ƣ�<���;�QJ����<H�.<���%$q��<ϱ5=��$=H=5=�R	<'=��U�8����<��:;;ܐ<'�<)�X��C\<�!��G���w����;.�J=�&Y=��<���Ґ<d$μn0{=� ���Q=�w<��)=Ik��%}; �A��U�=�3F<�fܼ쁦<�4o�{!\�/�/=�8:�4�(�U	u=.nk����';��m�3�"�-�/m�<[�<?���`'��)=. \;W"�<�ͼ�<��=Y��<��C=�O5=��S=&�=@����<xg�<��= �$�b��<OK�RI�;�_I��N9��y|��L��Zw�w<��a=��-=��=Q�����<>�v= ����+���ӼKzO�qI=��4�Д�<ذ�@y=�p��ę<,��0:�yN����;.綼N�ټ��<�� ���?���=�	��b�[=�B^=�-=������W�8K���G���ƕ<#�"��F�<�@��ƨI��!.=���<-���[X����ތƼQu���I������,�<�ļէ��@=�R�=O=�2�;�I"� <��\�N�Y�=Aem��[B�j`n��씻�Ǽ��[�>@ �<�	 ��%�b�$=�L����$�<m*=c;��@���<ӕR;�:K=��� }B���Լ��_��B9=�0�<��K=����m�h� ��<����u3�F��⪴���Ċ��[��g6=�
���k;`��<�JK��O�.�f<,�T<��8�3�-=��K=���<����
A=��9��_�'=a�<~
D=�l=AF�)�= %=�}I<��K=6˩�x�'�=��<�ϼ~�ջN�9=c&j�Jg��j��ᑼ`�Ӽ���;p��<���3/����@4��V=��A=c����+E_=ˬ���}=;@=��r���	�|��;"a<`#�=fT�<3�<i�"��6=REM<f[-��D�;��	=c�;��<9$=&���re=&�2�=�M�|j4=f� �D�c!3<�u�;��<4� =<��=����9��BT�<	]���s=�,���� c*��Kd=��w���7���$�^q=�<!'һ@TX=1�;w�<�狻
w<�U%N=�4
��C�<�:!�$�_��u�<��!��0�A	�5�c��7Ƽ(�q=�f);Yg��:�;�����:����B��jl��+=-%o=̹ܻ{�;�N�:�'`�|P`��L�<hC�ˮI=�+%���<˺,�Ǔ��?)-�l=�m�<-�=�i)=)GK<9'=��<9�F��|j�MX<��"��6ɼ�<�;�<�8Q<��=p���V�<G�e=�-n��_��-�?=��*���)��y�ɹ��SB;u,d�h	��{�l�Ӿ��Y9=���<�S9��]!�;H��W�c�$����o�T=h�J�c3:<	��<���<���,�N���E��M;=$e=;�,��<-GR�O=-vU<�\�>ܐ�l�y;�c�� �<�k=�@�:*J@=I�<6}3�Wu亿̲<��p<[8=~��<�=ا=�����!=0�[=��(�����'̼�㉼�kͼ,J��}��ft��x�_,����;p�=��<��<�`�;se<�`ټ��<o�>�>t�<hyU=ޛ�Dy���
�x�_<5EI=:�{�<w���}��:�<�t����;�c�<�N����=N51���<ᜏ����X��w�(=<�;=�J@��-�<@��:4�9={y����=S,D=��<�/<mͻ�p�<U��;�w����+ȼ��E�M�(=��<�V�<��G�e�=ʲ=_K�����:��<J_?<?�<�ቺd؁<���<������ƻ���O��<�+�l�ֺ
qD���<��D�����������sHѼ���̈�A*J=$I=��M��鞽m =�?��Ws߼+۩=z-&=�Dm=H��;%#n�b��<� ==,4�<��=���%��T=�����5��g`=z�\����<�V=7=��"��j=4�<MOY��i<�=�`�+d!<�=������<�8�1^�<�[>�~y=|j3=���;ێ�=��<Dw׼�sT=�����L��sv��b���58���p=�	��τ<y=�	��]:�PqV=v�=<��g��3&=�1���eǼ0��<�B�<���<ep=��!=��}=��;��'=��<�_�54 <Rj�2F��%�z=�^;�%�<�/�<,��<0V���<=�;�rY���=�F=!E�<��ڼfFr<���<�hʼ�wI=a0�;U��r�#=p��|<<Q�9�|Sd��յ<���Q��D��<�<�. =�h*=-��x��u-=��'=$�=�8�<s?��4=�a<������;�ս�2N�<U�Y;�4?=�=U@ٻ�)�<��<�x`=>x�<��q���8#��p�K=�h�<���=6���Od:=��<�&;r��<���<|�A��e(=�P��m�Z�&=7~��Lg&=�&<� �<q(�<EM$����Y�F={����=Rq�sZh<Ò��HF�Ԍ+=TT�5'4<���<��N=B=o�o=L�==y�C��꼻#=:�$=�#&=#��*wq=�=/tѼ��}<�=i���
�W&Ż�R-�Om|;"���h�<���H�=ڤe���=�8=����D���Ҩ)=U���1�`Q����;}����<͢��6�3=�ĭ< UI=|��<1e8���s��;ϼ6�;��H���b=&��zN�8�,l�4:�<�>=`E��R=�����C=if=���|��vL= �;b�<�K#=s8H=�O��P�&����_[#=���YM̼�v";�,=��U=��o=�j=�ut=������<[ �<����*��<Ԯ�J��M�"�%q�<%6 =4�ϼ!�=CG��0���xM=Сf��H�<|1��];�h<=UTݼmf#��D�PB�<1��<�����<�<�<�=��{;1P��=?���4�*�=n�j�_'�n��<zDX=�"=9�ڻn	�Y1�W�<�1<�9=b���=�r<���iJ��.＆M�<\�<:nԼq��<i1=��8 s=df%:��$�Rh<��A=4�M��H��8�o'���X;E㑻��=e�~�4�ҴR=��<�+���8��%��d��?�O=�Ǯ<�NQ=Tt�<�&��n��<������4<������<X���O<�� =��7��,�;�I�:O<��=�
�[怽%p��d��p�=�.�=���<\%<�b��<J�<�����������<�P��i�*=�m^�L�Z=q�N�W�����v��3�$�QI=��#=�1T���;�����h
�&���=��DV=���;C���=����<�¼JJ=�(�;<.�<cVV�y��<m�<���	��72�[S�<\m\�GYI=�(M=�n�<�LV�-�Ǽ�3�<�9r��6�LF=����J<����I����~=���8�;t�"=bk�O��:d�:9�<��X��� ��[=c�P�N(��H`�����N>���P=���<�&�<�ܻz4�<HѼ�=T��<�&=yL�s�o�IQ_�.�U=��$��R=�S=hJ�<o,5� �Ƽޭ=% =��P=�v�9`3��D��<�X:�0�d?f;������= I�<ƣ��&�q�7:3b<�f��<��� a=A���t���<`�=��U=J�*=�$�<wl��eM�Y-
��2<Q;����ɣ=]�I9N�m<n%?��^=��	���<����|��n�;���Ǡw���%������e��&���=��=BlƺO�5���ļ���<j��iV�F�(�(U=|��9}�t=���<B=�?� q =hx<F�==J4�<eлf('�1˃;�F7��	�?ּ��=qb_=k��������)��3P�����;c{ӻ��q���0��b�<nn�$�Y�S`�ֺuR�;�n$='
1=hk=Z���v����b=�칻��&�e��9�i=�FC;���/i=0��GJ6��᤼k>�<�O�<4�-=����3�L�w0�`=;�3�<q�$;J*;+^N= ���H� 韼aU�<�K=�Z�>q�Ɉ<8��C�<8L��[�<��P=�L�8)�UغQjK���+=�P,=!��;D�g�6s���9H���9;Y�F�@��<t<9�=q@Z;�<}.*���9�ݻ��*�QL)�5�E��gM=-0C<4'�/���4=5�ݼ���<~T�<ܻ�IV���<���<�%\<p�z<0[k�b��<b��<�)�;����{R�<tJ�pK�����<���r�!=ݍ�9��*�q���<�q��o��^�GK=bT=���;�XU=�+/�JF=_� <~V=�[�=��<n�<�I��s���=|�����ؐ-��;�
ϼBF��|���ެ6�[�:��<Ԑ��X=�N�<h��&�<-����:��*=i	(�W�
���`=I���	�Q�'=^ᗼ)_L=��Q��ڼ�r�����<�A�<��l<vO�<���<Sh	=u#�;P<=�f��3�<���.�:��g=g=,�*�W2�3߼�)��Fn�(F=k�<o��O�$�u�J=W��;�:��:�<#־����.�}<���,�;v����2��ŝ���<_�<�?@=�0������<J�V�lBO�r�X�:�3��</<�<��=��;*�<6�4�	�<�����S<S�5=�I����<1w�;���ڐ�;,|�;�Oj�yc=�����J�<g5�<==zA黮�{���g=��Y�/�A=M����9=�@�<�s<�����=.�<�5=���<x�7=�s���`���=i�}<&6=�2r�L�';h�@<�^<��.<k�B<<�';	�-<��R��tw=Z(�<��<m�J<��^6B;�I�;�؆<c��<�N���%=�U&���̼�G�;��5�y8/=/�<��=��z	=�3�=�#<�|�Z<K�:�e+�������$�:��<��M�������<�_�<�-='����+R�Ư�Y�ټw�_�<ه�0�;��;\i7���0���m=�D�q��;W}�-^�<Ø��7�]��	X�11�=1�6;H�H�7z'��]����b�Ѽ�:drZ:G�m��/=�N�<��D���Y=�L伿^/=�d�����<�H'=�p���|��X��<O�<��M��W�<�(�<�F=4,�<�=`����5�w�<D'�;ߴK=�Ѹ<@�*����梼���1����W%��6�3k	�\W7��YY<�ѻ�?���:��j=���qU==�!g=�ݣ�y4��"�Q=J� �Dd�r^�1"����:W^<�d<=X�)�B =p^>���B=�Ӆ�<u�<�4*=��C��HӼx�5=�GI�7}��)�ͼ��6�pT�2r�<J���?�;�1=!�:�ʣ���Ug=��+=�?�5���>��; �=�lg=�	�~U�O��W��'�T��(���傽��5=�+��Ԏ"=��ځ�;�;>�*M��B��<��X=�r�y�-�o<�~��T�;��O��̼���<�IH�:�J=,�P<��m=�#0=R:N=8F=�*̼%�t=�*Ǽ؁e�R���s�<i��f���e��{X=����=K�<���]��^��:�B�;-�=�����|=�7>����n@����<D�L=����.��D%�A�<^�=3F(=B����Q=Ɯ�U�=��&��4���4t<��<����c
=���$
>=�v%=[�s=�0��#ʼ�$S�ί�<�?=c�<��?<L(�&t;�!��=ǟ��E=��?���<ِ�������=���<:�G=�����!=7��<��+=��;�=��%<>����)=&|P;�og���n��=1,:��Tۻ G����>9==&Y�<#\�<4w<o5=WJk=or��Is=l:�<D�;=9w#���F�[=�5==�x�<e =ؐ�<d���4�㧈<�9-��aD<�#}=zcI�}�,=��]��<1r7=D�J=�P��	���<�2��S�&-�<]�E�a]R<�l�<� $=�F�j��<��K=^�C="�w<L�7=��R<>h�=AԄ��h��5 ��z/=�N��a%�;��ΗW=PW�?P=�A=h*�5${={�g�=���=28�*
��ʼ��<�]=o8���߭�G�?={�<=��"U =k;�;�Z=�B<�=>/�;��F�g�;d�r��@�誥��͘<0��<0V�������(�<�+��C��ʂ=�l�YPC="�Q���G=��U�0���^�߼�Y�
"Z=��=���<s���d�<��<��.<�x'��+�:\�;=W��<�rX=c�?��W;��Qa�!�Q��'�S�<i����G�O=���ۢN=�ը<�<�'=Q޼��<0�;�!��/7��J
����8�!�-z�<�h"�ҷ���5�n���}<�]�= (_�ݤV;��:�O���(�<p`,=�+��_����`�#�D:7�=<E_�<��	��C��t����q�_��wP��Н<FA8=�%�x�:�s�"7c��/@���c;?��<�[�7�-�qf	������5��o޼	Q=��U=��?=�IF=��1��<��>;*�=|�6���<$w�=U�t��&ͼd����	�4=A���<�_��6=��H=����Ѽ(�L�)�#��-=�P��M-f�n��<8��<\荻�=FU)=>�_=[<�Yy�߉��j�	��7<�"K�5Uz==�<?I>�1�;=R���|m��/�.Q�<�E6=��L=���s�>�͛g�t:�D<�<�� =-��;�@�<)Q��X:�v���w�;�7ż���Yh���_<z��4<��W<�C?<<�_=�J6�>�p��0=�<����<,ml=�:K=�S��#<y�_=�`�E���]���˨T��<�;|�<ː=�O� ���Hϼ���<k.漂h�<|=��:=w�<�kS=�20=ҮL=�p9�d#=�f�����`@Q���<�7S����;��.<ˆW=��z��"T=��;=]��(�;����(O �nd{���K�L�����<�.=<��$=wk=d�
�?[t�U�,<���<t�a=-�<˴<���X=�Ͷ��k <eY�j���e=��ռ|k=�����3=!8:��mj�<=���Ӏ<����q�z7<6״<�2��T�%�ϊ�<C�n�k7=�\�"q�<@M&�%g�;�w�<�v���|�<�X�;գ�]��<EU�:S�iv�|�d<�n�~��;��w�������"=<��G=�{�e��<�.��;�J�֗�����%���En�<C������<�������h=:Y��S�6=<�~����Q<�<ތ<��ނe=�� ��=;dn=��=�ռD�;�f�����<�0^�L��w؃���$=�D(��=#;����Q=��#=8�!<��h=�ʄ��A�FXO���:5=�<�sM�l�=����A���'=��<y[�<+5����`��� ���һ=E����<s��`�=?=�1�q��<�?[�*'���8��1���C/s���<��-:��=w1$=8md=R��u~=	9��7zB�x�a��]⼗��������<�s@=`��:ԟ����
��5;��¼��5��6��\���H�Y� �˵o�p�]<�OQ��=�T�L1W=�Ἄ�ּ~h�:��;����qq�<�S���n}<r�;܏���+��"�;�5�9�b�K�(=�M���x=ry��K��<wR�<{A!=h�7���9���S=M��s^���n���6=\�� ��<�����G�<؆4�����c�<��Lnۼ�Ƽ��@=�}
�U��_�#=��$��(i��k���=>=���D!=� �;?���K=d�<=�<Y�<v7��@�ʿ7� *=x�:��dt=P��<qQY��{��g!�<A=<��;�.�<\p�<��ܼ��m<�n�<qHK��_=1^�<�I=�����<�q;�ub�� ��ʧ�^[=��|<^�;=�
�<|�-��"=��1<f����>X�M�(=�20��4��� =<���8}���ɼ�$ͼYXi<��0�~;���;8�<�O��\v�<Ĥ�<�5:���?<Q&&���`�;h�"���l��#�G�n�<����u����T���<d��<���ª	=��!�?6<�3d=�j���W<b
輕<�����D<�# ���V���X<1��8hi��^=�����'�=U�f��ջ�h?�թt<0&=S��<� /=��ҼU��<�)�# =����`z�<F�L��>�<7	!=¾3��H9�vO_�m&/��=��S=Ӽ�}��%|=w�D��<@�;=2g;�
�%�B��<��o9�^�Y=*�4=D=�)'=�z5��g+�Z�=�d�b��<M�=p] =�vX=�����v�غ�� �<x�=N#z<�|�;�H��V�k =�x<���{;N V=�:�<��<嵥;�ly<�7�pa4��=ɻ\�Qk,=�/6=J��;��C<:�ϼd�=<������w�?;�-��%(d<M��<@Y��'���'ا<>Z�<Oͺ<�#Z=�� ��}��x*���M��&=0R�m��1��;�� =���;,����-=�Z��o��@�����<4t��-����*�0��;�<_�=�C�;=��,���¼W;�<)�=L>=^=}��������+=2:�<�Q`=o�0���:�Fd����<rL���l=8͘;����y�R{���\[�I,=x���o=dD=т`=���=ք����q�U%��i�����:G��K�<�� �ZY�<�5�<"�=����6Hʼ�zO=t�-�Q���@R=�`K���C�-=܀��*(��T�'��
=,��<��L=��غ��^���]==� ��f=A���'u(=���;�Kl�Ш�;2â<V�X<Y��c���c=J�<?�<�'3=�=�;��:62=��|;d$p�n>�;�q$���==��#�_�=��<=�j��s�A�V���S�i٨<Q������;G<$s��#�޼�hY�Ш2=vVڼ�ļ4~'=�?<<���=���B�W�̼�;�W��{�F�༈C�1�޼����zh/=�W���Y����;��<U1�<H�W=6,B�c�+�i��>@2�[ټ��<���V0G�ZG=��t���J=���<��<V�1��=���;d�(=u�J�,={*��	�;���/=�<l����S��)�;���<-G�<�O�<�ݒ������x޼���<�K�<��<r�=J8=��&<�����~����9��=��+<�D[���<藽%���x=�sy��i:=��<�q<4@2�G����U<���Վ�<����];�f�Uq<?S="�<��<?��=W��t��F�_��n��Y	=�K=K�ϼ7�弆>F=������6���a�XP �	��=F��#��;�q����5=��=:�$����<�B����<^+���|E���R��~���S�<��Ҽ��<�F^=:���I����9�1?�ևM�b�o �<:1�!�.=J� =�L�� S0=�L���@<�'ݼ7����F<���Mc�<���D0=n�<7h�<���<�X�����6�<'O�5��<c�g���<=c�ȼ��<�.��L�7�ɕF����<W���,�p3	=�F=� n����x�&�׷]=��=e��<g,��O���>�c��iW=k�m�3�P�b�H�h:m<�}��S=Pܟ<�?^=��;�!=:�?<��<鋨��gT�S���vX=�D�<,�7=��r��
��	=�����&<!�<1B��+0�<���0=e缡4�:G*�<\��=%�/�?���ӻ�e=�$I���ݼi(ӻ6�<�]ӺU�m=d��4YD�U"=��=���<ॣ� e�3�<��ȼ�+=��<|��`r;={�y=+�^��3Q=�k)=�{j�	ԑ�[��;l�<��\��d=�$B=&b1�Rv�@�
�� ＃ =}G�;��$=]�g�uT�<
R�eR1��k�:Ð�<�.:�QP�; 9�wi;ޣ=�䃽A�]��M��Z��@=;��;WyF�8?��Á��:0���.=��𼫪�����������ڼ3(=��r��-<��S���;��w=x����{�<Ȇ�D�D=�t:��3=!�b=�r�a���@V=`��=�T�<1��L<�y��;��?�$=���S�=��; ��;z�伊O_�)���+�b�֯%�
�������N=7;�`O����>�h;���<�9<DF=jTY;��)��;vw<2����u=�jc�Yl<�'E�My<�u='���]K���<pg�,^/=�»��=<��<C�h<�H��A1�<��"�\=�,=M8E��z<�+=�-�<�+=�j=ePX=��>=�值��һNl�<�TP=��< Y�;�Qļ���c� �W༬�Q�22-� �G�3&Q���*=� =�=��	�lTX�!;ټ%`=#�<���:$���:�������<z���:��	���
�=���큖��x=�ʧ�A)�w�K�8^ռ|��<�W=!�;x�����f=����=�o1=i�=���=�0��W�<i�<��[=��=��<Vm#����Oh�l���q�eF�<�h;��U=B�@=��A�����s��دe��>ڼ�lv�"�i=;M�:B�(=t��+n=}X��iHT��>)��ּ4����V�9�y���>=�s�<Z�=�&:=N����S��&�4�=�v�!�g�zT�bu��.4;wű�NU �:.����>=����u=���;�'���Y�<�i]����<�x<d��<3�=���;��_��)��7N<�������q��3�Ѝ��궼�O���a=�I�$L��G=9x <�����<E}=#��g^������N=B=Wi�;���2`���6�~���=۴}�-�J;s����=Kӷ��|y�dK���:��ۼ�经Gh�k�I<*E1=���<���<�(=0�]�a듻f5_=q����g��w��:�<�w�������<m����z�<�'=�zg=��[o�< K7=O�P��P=�+�'׻�K0<�+����c�r�⼰;=��_���3=h�\<ֺ2=?��=�ּ��3=�L�/C;E7 ���<��T���;����F>�<r�$=×���]<k�1�{hI��Q�O)��z����<�z1�2,�<��<<���\<L�����G�>fq=�Q<ܫ<�˼^����V�<�$=oia�N"=�&�W��<Ϝ�<�0=o���b��;_�<�Xc<F��<�
�<��F�`��,���<�U3�K�>�{:=g��<1������<��=�j���-�C�,=����O߻#&!=�.м��<�;<hD@��t0=���<�+<��<Z��Vv<]:��0��tq<��K;��&;�I.�[<��=%16��� =ۗ=�$=�D2�X�;=� �<KN �VZ!=3�=�����h��qg<u]=?/<2ۖ��@F��D�E�4���n�*<��L=;m����<^�x��tB<ɖ�:��a���
���"=�?=z7=�Y�H�a=��"ܧ<"�:=�=�<��<]�N=�]/�oҼ`�9=\A���K�!� <(+�<�=��<띘��i�������^6�de=M[b�6}:<U�@�c�==k6=���;�*=�~=ʇv<-�:=#u�<p�C��#4�rC׼iC3��+~�"�E<K�=��Q<��;�P��9�i�k<�~>����<.���.�9����G�<v%=�aI��O.���?��<x=�A;à#=��<�|$���\���h=��,=FK�C�*�y���(/<P`����:�0�<�����m:;2�_=���:fn�?I�<��x� =ZK$�Џ
��;�<�qP=`u=s�=b6>=�����J=}����{<�a=��R=�IY<c�;�#��bG@=J(=��J=%{�<3����U=��ٻ�`fۼ����h*=e�=�DQ=Ҵ���v=���:=]�\���w=�tb��M.��3i=�]B=1��>n�n�\=�73���C=�6��5E�&a��ǇM=F��Ə_���Z����k<0�T\��sƼ���xX��e�D=����mqt=z���a@�/G�2�� [�:���<|��:!w=˫P=dT&=�tK=�#���2�==gS��6��<��ļ��s=�PB� �{��8=t��<*҄�Ws��\�+�\y9=�]-=�� ��<�\=C�"�-Ӽ� =��R��\d���<�.K=z_�<�TB=�$ռW-=M��?=�]�t�/;�Q*=k�<�2�t��<ٙ<�)��/_����<��r=���:�F=���]<��7$��q�~����X<�OE�ּ�����j&D=)�<���<�<��E=����ȼE�f�|�=9��g� =E��21S=a�8�\�#��r<��;밚<(�\=գR��i;���S,�<�ܼ8�B=�~�;_��<y?��;�L�:��v�g���պ������3��;6�λʣ$=���Y�<d40<��G��W?=�b�<MP$=���;�4=�(�<�E:�	��<9�Ӽ��V���L�:�!��<=��U����Y�9=���L2��<E�ch;=����j�<�����⮼V��;�Ũ;�{<��Ut<p�<�8�T�C9Yz��!-=���N=Dz�=�伊n<�j�;��N=ٺ�<�l�A�(=�Һ�Vc���=��͹�p��M �=*q&�w<lnB<UJk;UT=V�!�!=��}<Xޕ���"� u�<Bt[�w{�<?`�;�q_����<Q�p�?��<��b�D	�a�*�(�<s ��(=�46������G��������F���VF�D�&=�,���%�;�#�3=��H�H3k�ƀ���;N>><N=�$&=��U���k<��.�j�D==�<8�<��J��:�*W;�����߼�-�u��<IT�O=7`6���: �o�1U=J��<���|	���Cֳ:3����<�:�4�<�W�;��K<K��<��؅<ٚ.�0o=jS=�o���;A�<��+������ <��=.]=�@�<u����=.y5=[s=Z�;��;�!�<�2�f�#=q0¼���<��Y� j+���=p�U�?J+���<H-Q����׼�=�"�<k�q=7��n)�B�Q={G�=�
��(�a=�7���1��;�������E[��X�D�=&H�<+Qh=�c��<Z�;����� 5��nS=%n�<e*$=��.=��ƻT�����4;\�M��:����<�़�'�=�˳<.5ɼ��=���B�A�;�#<�U��ZѼb����� =�u�Z=w:��1�<*j���==�l�%l<�B=��F�<SO��)��x�� �<�����=�(��4�q9u �=��!��:2�dмQ�x�B �<-�]���6<!ڒ<�~5=�
<��J=|����_<��=����L�:W��&�O=�5<���<8�	=���;�2�<�]<�_�ɠ;l�<�K����=�һ��m������0��l���= '<��3-��AI<�ug<p���v���B����=rKf<S0�)֞;q=��5=?2�; ��9���<ì,�;�κ>��Y;=OT�<|�*<E2;K�b=W?4��q�<��t��h�<�V2=eU;G^��O�f�b����2/+��Ӽ�o�;�p��R�u���w�!�����=�=B���g=�k�;sXC=��4=�c<�C=v�<m���<<�4=%>G:�����hټ�f/�oM�<X&�<��><�e^��a=������z�<Ա�<�j=)E9�N�J�0��=j<��������<!�<�-}�|�:�& <���6���cv�6�^��2��Í=4�]=t�G���H��_=��	;�_Q�E#P=�E��`U$�ky�;�x;<��;-c���<M=$b��eb<��\=o�&=K<<z�&�vB�<˅s��f$����b�A=oO�=��X=8���ےE=��=z�=�W�=]�[�Wb����4=@s���o���D=�h�������������:9;�Ԧ<ۯ���J6�����W�=B=4�<�-=E86=E��&�<_tC��+�]c?<D乻��$� O=O!;�%'�g��<Cm�2�<��5��S�s0=��W=[[$=צ����3��;��=�iA�N/`=>�A<"����J�	(�9�F �-r?��Z"=5t=�s,��RɼI���k�;=�M;j,=��!=�[���<v�B���t=��}=�'�~��WG=��M=�Q= &7�p!�T���NH�uT�<Q�b=&�=&��<�GqD;u�8�t�M=�;��<xo�
aU=CQ��J%�J%=�<{���bإ� @|<w��!>��/I=�<�	 =�N�:�=C�b������s�<���<^��<��V��k>��*0<��y���.=C��<Q(=9�׼����Z��K8��9=;c=�.<3�Ԥ/����<'z�<M
5����<��<��s��J���	_=?mQ==��;��u=��)�j��<aI���P������p=<k�};SY}<�J�Z����+�df+��
=�=yⱼ�%�<���<t�'�8=<q��Z=�������!��	=ݓ�:8+��$�C��� ;����.�<%�:�j=(P�<
1`����� ����=���qO����%��L��<�ȼ���<͌H:lW��Ry<�/=a)l�h�<<��<Ù�<�ܙ<��<WN$<��Y��=�� ��r_=ˇ;����q)�*$��r���<��:����h�5;,=*Z�;-w����N�b�Z=<Y�)��U�=��m�ɼB]��)K�B�=k>1=�(;켼D#=A+�:㉹{���<��[h;�c=�2�	�M����;�"������C =!���+B�N=�B��+= Ҽ;��N�|ב<�h=�XO=Y1�����(�c=7�<C��p'��@����G<`��_�� ��G�<�W+;j=²��,���(=͇�g�1�=p\��Ym=�9�<�ad��Ω<��B=9�<Ex���hm?�fIw�TKE�3�='3w�V�����Ⴇ< �,�>��"����2;��ּQG�i��;���o�<���'D���g<��3=���ƽM<���;���#Y��l�#=
�+��y�)��:))\=c��9�v���-�<� ����C=��"=h�=,oH�ʩ8��_�n��H�<�Ļoc�<`��Dٮ<��.��D��=7պfaE<U�*�����
�;H@��V�Y���B��)�<@���8uG�
�=�G@=!8=�0��	=��c;��,=8�2�X�$��#��V�<��`�_����7�,	F���L=%,=��"<�м��=�m=���</4=H�{j@=6&	=��R=<��ٻ4U�J�<n�g=�4\=l�����^�=��=&O#=�͛��0=�鉼k�=���	ټ�*!=q��BJ=��� ��Hґ<�В=HY*=%}=��J���q9�;�n�]=��%9�T��5G�c�:Շ�pD����ٻ B�<��@��_<+@�<}� ���B����<vz��-���h;q�}�5=K��=�ڻ��A<H�����
=��\�R~�<�=��0��?=y���p�<�T=3��<�k�����������x�4�y;��;�z=z�3<��X<����t</B�FLF;na =vV��o���;��= �,=�ͪ<Ð��	�<bؕ�B�>;f�;�6�D<�[C�7�X�?�!=������<�U=���<�9)��$���v���=��~<��=A��u�1�<|�C���3�.�;��ݐ%��m�I�7<�A]��@��Z7q�Q0=R�?=�h��j���{��D�1:��8�,�L=L��<{���8�<�5m=��|�)Z��B;�W?G�<0\=EG�<k1� H�<�����ʼ�N��!6���=��H=Oŭ��= �r�S<��=o�=9pS�Vن��͌�P��;�y<�A���`=?Y�����ZE�<'c�=�&B�um��������<?��$-�(ѓ<`���=%=;�K9L=���
Ă=�5!��^/�N���g���p=K�Ҽ�����b��Yμ	�;�AƼi�K=?�o<�d=,D�;�=�d��U��<�u=�=�G��xx;-Z�<c�=�w�<��a�-���ܼő�����Ӟ��I��E��x�<��̼�[F�׵����<��߼� +<`ϼ�I�<�lȻ*�;#�/=��.�U�2��"t�Hq�<T��<�=�=��K�8:_=��[<Y��&s�~�<��M����<j��.�=�w�<��������,�<�=m�9�O�3�)���>��ץB=0��:� ;֑q=~O�\�ټ׾�<�S޼0	���(�?��<��Z=�2j=؍�<��O=�c=VDM�7��漏�=�u���<�Wb��f��q<]\<rޞ�&�4�CL�<�ݼ� r���>=+/�D�=C��<'{���9��z���
�\�U�f=�<_��k�g�p׼8�3��\"=G�9���G=]�p<%��fdg=R��<��0�f7m=�Kp<ta��x=��<�"�<�n�:���;?ef=�j=@�G;x�R=��=�[~<�ʶ;9�&=ݸ}�V8N�2�&=%݉<v�#=�Os��Ǽ;4Χ�
�=p�R�K�6�V���k(<�=�6*��������&�=�y��M�d=0�/=��=q�J=6�;4)3=������<�#�;�$=��<�v���=�-�>R��=b��� ������)=<�ڑ���!=��(=��l:14��W'���=�4D=�m<�;X���=�E���o�<q���׬
=¢)�*����=2��f����]��a���U=��u�/�;c�<}�	<�"=tc@�٬�<��<��;i�=���=�Q�:#��<9�����&=�p"=_��:9=�%��Q=��<+{;Q�P������o@���S��ܼdRV����<�n(=@X&=�TG<���<�=�N�l�Y���*B���=�>^�;m$X=�k=q�����; ��<O�<w�C=eﳼ���<z;�<7��<�G�<F� �_<<��/=k
�<�υ=�N�B����J�;q���`�ʼf/�9�;-��<t��w9
<��$�<�(�|��<��G=�鴼�=�z-��6_��� ��\T�ۉ?��1)=��M�;k����P�ټ�����b�<�/����L=T�:�+j���N�X6���,��6�<ڔ��y&=v�"���=��.�K���k�>=g���=0�<�6=;sϘ<7����
T=9J�;/d��K�<;\=�-���gK=��켙C+� K�<��< O=����2=��;X�6�����`�:�������:�6<Q/��2gg<�g]��?�<Tzy���V<3�=�<�I�l;��.�Wn�<o�b=�YμgQ��뽫�������u<�M=g�F<-�<�=X�;D�N���==��<�Er��>��"�/���q;'��%K�����9(Z=p�<el!=�f7=��_;K�����v;b�1<@�#=e��<_�����=�N�p<�;8$�<.���=|[=P��b�!��8�<Č;v���@�w	<�d7�&`����M�JN�-"*��<��?=��F<ď=8 ~<��%=�w#���=s�<�~�;Ӥ�<�{���� <�@�<�F��b�<B(¼a�f�&��;�2��}=��=	x�=�m¼�'�����<\Z=��Q�S=צ<�HM�l�<�B�<�u�<��m<�g���1�;�=Ӌ���K�<��8<�Lo��~D;R7�=���u}=ߚ����K=�d��`==��2�u�'=�^j���j�r<\�l��7#�᛾�W) �t��<�_(�kG=B�ϻ�>����ѡ�<$�~���=,��<//=?{=�>=zv�jBd=��;��U=�����3R=2�G=R4#����[�K=B�=X���� ����h9d��ۺ[|���
<͖�<,�����G4/��=�Ɓ��<7=M�.�)!<�F�<���<�<;ƩK���J;	�~�w�-唼�@�<e.�����p�=���;=�-��$7�z� ��3W�<!T{���;S5��/��rR;ύ�<��;��m�/6�<�t��:܅<,�<7.;������<�8<iU��S>�31��뼇�%�Ί?<d�n<�(P��=lpo�-ap�pv�<�=��=m麺��<�����g<t���R�r�ez�����<D���V�ͺS��
<@'8�>��;�9=DKۼ1��<z�s<��:�-=}�?��f*=��y<�,�=ս��h%��H,��p���B�% =)��<>�B����;�=�<N�;cf�;�|2<�=����<��j����9O4I=��l�tV�<Yc�<�~�<�=��<ϋ�<�X<&X=_��� �<�:�[�><��=q9=�������^�Q��;�=\7�{��� zb=˙<BD�rid=��a����<N.�<�S<=�.K=�$�<�}V��M=��y=x��<^D��V�<$���O��!&��[��P6=<�je�x����z=R/��)��e<��]������E��٩����b�=)"�<G�
�"�A=2�.=���<��������XF�۾�<s��;�+<`�s�N͕<_D=�����O;	g�;�2�K3
=���t��<��=�;�"���z�\�T="�/�ͣ7=(�*��R8=G�q='�0< ϻ�����G���Z�����K�<:|�<f�c=����=�Z�A���+<Û"=o�����0�=�1
���L=(�=��g<`߬�#�C=��<��!=}�X�90���%�|6��܊����<���<���<���=�n)=T�^��̓�:\p�� ��QW��c�����.Q�����<o��<I�=��
��a�1UW=J��H%`���<u=.߻L˂<,���<"��w�.=��%=�!�<_��w�o���F<pf<^����N�^�
��d �)>��%�Z�2ے�t՘��AW�����u����<��2��&N<B���k�<�K=6t~;��x<lA!=0����$=�Ǽ�+=ֈ�;�k��
�=��5<�=���:Pͯ<1���m�.<��<w�˼v�U=�U=$Z�����;Ot=2��(s�<�D�C��;�4мQ.�<v�P�h=4�1=j����=�g�<���;.nռ��o�ɲ\������=�V0<�
=w:����\=̄����^�F�o<�����M��	=Z�=��#�)�<��v�n{G���R<6����;96�<;4���6=�'���b��J�)����11=��:�)=��л�3%;A�A<�^�<�Xc='{�<U�W=�)="(���#��Y=����	�l�#�`�;��I=�I�����<�Ѽ��%��~=��=c�6�D�=v�d���Z�<k������M���H��cʼ��=�"��/<_�b<T�<W����T��������<�Q�[��:�
<�"ߺ����d��6f=%���s%�H.��@����<�j��&��,^<��<�iP=��=}�L�J�y���=�jx<p���.�=�}�<��.=Mֻ�(;"��-?�<$��<p�<�L5=�ֆ�뙴�t���=נ(<��z����/:�� �dy�;<J=����>=ʗ�b:7:m�!=����1=T�\=.���H�[#�<a��<�7E=M��:��<M �<e6;éK=<X���+=��J=ca�� �*=]ϔ�-P�<t�x�JM=�i��z'���=�	Ş<�M=J [�� !��ZO=�ǲ<ߵO���Ҽ�P߼�=m�
��|��<_�V=`cG��`=�;�X�9�@=1WB�8O]=u��<w}U��A�t8�¡�;���<ؑ�cOR�L<ѴU;���<�qc:�AB�b��%�B2=��� �m=z)<>K�;Y)=�/;`=B���
�5�	�N<-�B;�Ի��<��{�<���ó?��,G<��&���O�-��<�Z��k= .ļ� ����<�����D�<�sE�e���y1�<��� ���$	�9��<R%&�.}�<��:=�2��]d��C=|�G�=�4Y=�ޅ<� ����4=��&��`�<?T:= �6��K���L�R*L=F����l=>)�P<7@����r;�(�<nF �ճa�ra@���{<�=���5=B��R�S<F��<��=�}#��(\��T��4�˼��<����/�P<>��<��J={`⼹m�<�r�<�`=�6=�2'��-����3�&���9���ܻ��?��!�ngr��Iq��,;=��[����^�M� �&=�=$��<s��<�7.�m7o�u����@k<W (�P�=EG=(�<[��� +���>"��~���.���O�<gx�+��<SuD��Ƅ�+>��f��=	-l�m���C�;J�<��=H�Q=�5=\�?=?��;�?���4�	�8�SW=뱪<�!�<rQ�<<8���^<�=�n+=�(T�a�,�R�G#�<+�I={�0�u�<e�D���G=I�)=����0\g;��6���O��f8=�<���<:<�0=�wV�B�`�(��:?����[��B�<\�9;�<��K=���#/��[��x��}�O=h�^;��<��j;�@м#Tx�N�޼��=\|Ȼ0�B�q�ֻ�G��$����/T=�K��6"��<2���*|��XM��=��G=mt�<��'�Zż��/=�]�FWJ=�c4=����:.<�&<�	��[^=M�d;�=!@�z��<�'�<�7���$��v<Ê	=��=	t����s=�T伭[�|��z,L=+i�,��%=W�M=<�K;����*/=?���W�<��'=``���JL���<l-0=�x�.)�V�����Ǡ.���>�7X�Y�3��;y���-=]ai=(��p��pI�=��a��g�<qVi=-!;=��=Q+;S=�;�<��
=t0���E=v#��<="G�$��<�C�=�yѼ�ï<����FF� �@=k=;$���F��	a�d4z<�(<��2=��<r��<�n�<�h�i�G��,h:T�9�0��Ϻ�# ��A%�b��Հ%<٭ۻ+�n=�8��9V뻃��=�6e=�����i</��<�tw�frE��T���w�<�%=�����%=�<�<��;������<C�c�XN)���D=�_L�(w4=BݼSd���A*��b@�{i����>�a<�R���<��8=�����6�<��;��<��pn*<T�˻e�t=�=�C=�ȼ���;��L��c�<R�+�uPj���ټ�ʼz�V;�(�Xm�<(��<y�=��e<�b'=#�e=�z��wK=s����'>=�#$;�3=��	��  ���K<#nD��QH=��5=��F���5=�H�;S�-=�A<=�p=;��<jʔ�aŹ��!<�턼J�<M�<��N�ۄ"<��=ZQ��=�}n<�
���	;Q�'<����:�<���<����0����=|��<�-��lQ=��,��=7b=oNܼ�6;<N�;�gm=��=3ߣ=������;�<@�<����|���<��0=�3T<�V����<�:�F{׼*b)��9 �/a��<�m7=*f=9 f=Y��;���Bѓ�3 =JP&��=A�{�ļ��C=R]ӻ|��<�%�:6�"=ϻF����y���:��5E=S��:w�ϼA^���� =��=z���=�O�/����[=�}�<t�+=kS�<�e���/I�H'�b_/�O_r��*Ļ��d��2<���;�������()�h@%=�=l�J<����|T=�=W)�剠<�d8?�����<j�`=��	���Z=c���7=�(�<'�D�ߘ<��)������'�v�";	�'=W� =� �� *r=n9�<Rk:=tރ<�l���k�< D�<פ���u���ꌽ�Ə����	uh<��q=��=�vm����owŻ$k��O�W	�<��b��<�w��ټ�h�<R�E=G���'�<�4[<ܘ=�I���g%=s�;c�=X[=f0}��6��n���<�=$*w<\���"��׿+���=�\��ߏ=#�><ћ��A(� ����Kc��x�A��<o�E���<��<sJ�<�0ɻ<�-<T�<0{5� �<_�:�6�=�WQ�<	
=��M9}0=��<�/k�<PP-�z�<l���=`�������ܻ˵Ǽ" �R_�`�=޴Լ�����lK<B���=���2�=u���s��<��%<A�<�(E<����Yp=�=��$�߲�r���k�@��k;�6���49<:`_��/�<�4=�	�<��=[vT<�u�<k�b=@ļ�hu=�)�<�D�:b�$��Y`<�=��j���A�]:<�T*=Ə�9�F=��ҭ̼�8<�q	=�^=�6��#=i,��K�C=x�u��v�<�/=���1r}=d�V=)�O��9�ldd=_��sY<�ӄ�ZB�j	��~���c٤�E[<��Ӽ�:��h�;�p!��6=�z6=��
�=�J���;D����m =Y<�_-��&=RI�O
�� ����qG�ؼ��VSI�ұ=Gb��%;��������=���J�_���P��i�O���5;��/<n�=W�O;�{�<R���U�<,�����=�ɽ<�8L=cd�<���� =D.w=�rg=H�μkN�7Y<a���
�0=�w�;L�r<xF.=$�=�@�<�/�;��<�g=��o<��2=A�f=-�G=c2T=;=�Eɻ��t=��W�7�����<��|���O�"^n�΍=�/=�1^ݼ���;``=�==���I�=g=�[9��E��;k�ao5<��=�s��K<��<�j߻��0=�P�;�ľ�_�=��.=9��<L�<1�<M;=}Z�</%<l�ܻ����I-�;��5=�?l��`��71��%Z:�$�����<x	<=u�L�e��;I���y��8�,���<��1���=B�ۻ��B;`@=N��<DRb<x�g��}�<�}�;:�Q=l0u��u%=�H=��<����\���V��8���]=��8�b���S=��k;�iD���t!=	�ͼ�[7=/H�x>S�B��vܨ�>�S<l��u�!�,�<=�=���=)�K=3)[�!�<db6=R�����=�!=Y�2=�s��V���=!u7<w�	=_p��2c1�̧5��?�ѷE����<}<U�|<*�r;�G<��<��,=r��=�;�oW��@���)�UU=��C��	һ.q���7=y��<�M/<|�}e��yh�p�P=C���7=U�=�3=��u=�l<=qO|���=�! =��6�� ��jü刐<^(=�:O��ü̰�օq<X�6<Q=�-��G��9�{f]<�N��<H��<༡�l�p<	b�<P���0����5�!=�:<S�G<@�W���\�1��$�E<�%=m�z^�<a*�k"�=>w>=M	�<�S�7=��Q=#�A��C=���<gR�T����5c�q�#==J�g줼խ$���).P=�r�v ��g�a=�^=v 鼇��<fGq<�B�;�,=i�]��t=�2k��w\8�W���z����<�Sn<̬�<?��<}6=LF��H�< ���/�<q�$��[=JW��=��������ほ�Bh��Jr�h$<#��;Z"�<��=�ͼ�G�<,Bܻ]q�<H�
=ġ�< �L�<A=��M=y�=fHH=�q�;��4=.��!@���<�\2^<�)��i�j�<=���pie���=4?	�6@�<sB<�.=�ey=i?1�芺;uW�9==1g:��*�=ǩ�<�劼!8�<[�{��p<��Y5�ͯ�<�#���J��LE<QN8��b�;v5��G�<�X$���ϼE�=tI=q(O����;�r;>�.=%��<Q4R=��`�
�ɻ�u�<��@��x�9���l�f=����I�v<�	м0[q�=<����_�Q�a�I^?�_������ԡc���s<��3=q�<4�b�V7Լ��S=��!�_t<(e��+ s�(q8�YΧ:�E=�.v��i=��?=caͼ��!=AL��G=6׼�C��Ŗ7=�1�l�U��0���Y=(Ֆ=��)=����F��=,~�=x�A���W��*<�I-=��<,��yx����;W�p={� ���9���2��,5=]�L=�6Q���N���g��1�ċ�<e;ɼr9�<#��g
=U��[��=�$��E5<�jj=15�=q��<=P�5���̼&0���=L��~��e|�*�<m�������~��W5�Iϊ�L�\�'
=yj�:�_�Fq=��4=m�s��&c=��:t&�����<�ۗ��W�=&�5��=�<�r@=Qh�<��S=hz��v���6���=�5�����WH<0���6��:�^=�N<=��=
�;Ca=�0�<k��g0=)J���ü�
=}o=�0"=���i-���S�d�8=��_=5Zl;�!���J����3b���=�U=��+�+�tS��+�*���)�B}=��K=J)¼���<������!��L6<��P=��T=��t�n�L=�=�΍P��-=Or;�,���E��?/s��Q;��;L��<�e<�����$=.c�=����g=�{N���,<�ꈼn�y<��-�1�1=�����<�e^=��<6�Y<��r���Q����缷�<�m�<"���R�<��6��k=rv<��N=���<�����q�<�!6�(9���?��5<�d��$D=(�e���wH=�kڼ��0�˳�<���:��=�v5�d�C�0;Ҽ���;�զ<M"L�]*���H����[�>�7�>=�'�<
6���1�`��:#���i`�<��?<�W=�5i;�c<!Y������I0�?��LҼ� =�l=�s<��t=d8�</x(���u=mW)���8���<��e<$*!==��&�a=���a=SFT;�h�<%�<�H=�Y�<���U|ǻ�Hn=������� ���c�X�J��)=K�_���w���<4츼Q�¼z��;̦=�=oPG=K��<�;���< �<�����:=)������^�<���䢼#�U=ţ=�0C=�����F�m�%/�<���3=�'P;+hg=Y�=��<?����b����d�=PO=�`)��CY��������Z=�*H=.��g�D���_�������<g;=�v[����8<�W���=ca���=��#�;��q�x<��� <�
]�bT�מD��t�C�W�=+m���R=�X�<��X�M�����;�P%���[=9<B=߬��@J��=4�w<Tt=u�+=�ҽ�ֽ	���X=I:=o�b<�H=a�:ڼ���=x3;d���������ݯ<��q<��;ã%�f̌<6!2�kH<��4=��(���<��s�O#���D��򷻧en��ka�Q�B<L=��(�9�_'=�<<l��H뻴�;�w�<�:=57��R~<�;ۼ�$(<߀�L��<��+=5�<9b���M��r�<�|����<�b=�;�L'�����S=��Ｆ��<i���oT=�N|���<���<�	�<�]?���<Q��0*t���R��1=<�q�&0�$HK=g�^=>k<��t�23=�=����,���jX�i��}<�F<��?=Y�¼�	<4�h�p�OA�<�����=P��<D#�<k�'��(�� �<���;Ч�V�<Z_���k���=%ch����+<���-<�=#b�<J�
��X���?�� v�<7WT�,�<�V�����<\�<�%��_l��9#=Z�;O�F=�ü��1=��=��;� s��(G< K�<'�j��,i��NX=[r�<�Ʌ=�W�n�`=�B�K٨��<|�&=/��;�	����Wv?�P|k=��-������Q�[�7��jX���@H���ѻ�} �"��!P=��	��I��G�������7� p�<I�'=�-5=��J��Cv��H���p<P�������Dd=�F=���<���;$�ؼ
��Ź��������D�<~�׻fA��Ƚ�R3��!==
�����,��7@<W歼�\���6���	�9����];H�5��[�<���;�A<�=�<_#}=ްd�%�<��߼}	=-�/= *��?�����1=F�b=<S�|�%j;��?�� ��Bl�Z�<���<A=��:8&<�����o�m�l�_=j��<��<���}�$��]=�b7=�2�;s��;�k�]���ܵ<<��;,��;֫Լ�%�$�d�]d=�Mֻ�e�����(�ܻp�]���<����+M<(=U�������]���*Ps��-�X}J=��;���<M�j=%�0<��缬V��:���5=�W<[TF=$(ȼz#n;��ּFBV�b6/����p��[���@�:=T*1=�1%=@_=Ǎ<�8!=��[;s�<��x�hj]=��<�#㼰��;�3���=�^���� =�!F��I�=�%ؼ/�%;� ׻S�ɼĎS�G�l�M�V��隼�(=Y����l[=��+=
+���<��-�N���<"D�ۅ޼9-=K%s=F�.���K<i\;;�X=��p=�����:��<��6��'��I��8f���ֺ�X�w�r<��=��o70=T>���N�I^�<�P==|=,H�:�\��M/=?c=`�<f<^��;3��<T�$<a��<<c=��J�x�	<�*��|��F��¢<l,�<�>=�.S��$�<�|λ���<�x�<�U;��O=� N=Wʼ�#G���= ���P�N= �4�f���B[L=Ĭ<=C�*�-��=�>=$�c=;���������g�A=�FY��鄽	��wL��pe=ه���:n<t8�=�h*�T��z�5H��3�9��S=m��<":�8�K/���;\2!<�K�����bK��x"���R��~ =��5�p�F��R�; �K=�c��(pL<���l�;�d��;<o3�Y�;�P&�|�>��'�39K��U�����<�/�<�H˺d�>�����ļ3�Q=^8=�y;��Z��Cr;ϒ=�>���J��j���c�a=z��_=��v<]�D=j���r����������<鞕<URU=S0�=G��<�/ּ��-�;��+�©�<�@==IG<j�'����E�%��3s< a�.�G<��;��A��
�<��<^�<���;���<�Jļ�ߪ����;;�üy��<J>!=᷐<O�<�_���ļH�=M'��h���8=�D�<�{��Gμ��="k�=�'�$b<�=4~D�}~7��t��+�$=��^=`��}#i=oƐ�lL��;U=g:����H=�)�=��s=)�=�~���B��K{�C|<���<����ͬ7�Ӻ�;ߛ�<�۞�+�<�T=�M4<#�5=yڼ	�@=�?=�N�����B���ē<f���l;Čt<�h/=�!a<1i��xʅ<xq=����}�<B�<�M�Q��I!I=ݧI=�� =������%=O�P<��P=qAU�(5����<��мn��<m��<��t<HY5�1�L='����d��C�x��=���<hC�<	�@�b= �D<�	���S�<����֑��=����3����<=��;o��S�\H���6=��pLg=b�w�s[W=__D=�a<�'μ�O&����;Q.�=b.=��w��m�8=�񳼱��<�3��w��B'=͝��m�<9hF<έ1��TؼL���T���:?=��8�t�x�)�	��<��'��}��*��SY=Z}��'N�{��<TJ�<&qU�o��<K=2zK<��W��`ּ�!��JD<-�Y������n���9=���<���<��=��S�=�ģ���==�p�<q�!��ɢ<C�="�p�L=ᭋ<)�73���65'<�� =F���f�7>g=W�=0�ҷJ�,'@��5���N���ۺYYB���G=�\1=�N�+��ɯ�s?�����R=v��6�qe�@Q�<z���C��_C=Z�u����El�,�k;`kȼ]-��A<�>������<�����;�lN�<=Q޼]�<��?����t=�'�<~`<�h=C2[�C�<�X<�t�*�<E7=D'O�&�<]�a�@��u��<H�ZF�uP=Gڭ<��9=�L�<�d1=�<��#=�.=���<i�=�I=��(=���%�<���;��ۺ3�*;{/Z<��û��ـW���3=T?A<R79���y�e<�T�.���[��<P��<7� �ڟS=�z=�/[�I�;�y�<���m+
=|��0�:=	�=��sμ�ũ:��<#
=����vTW<>7=���N�e=�@Y��9��e/=��Ǽ��@=�پ��x2=�{�����fPP�g�2=hJ���"; @7=��.���(=`����6⼿b߼��<���<��v<�H]�"�< ~�Ϡ�m�;<����C==�y��(D��仐�=���<�3���5=���+���';c�:��X�<l�>�I��#�������X=�rû�=��� =jǭ��̑�q����u=Jy_=����}��<9�`�<==:��"=���;(�պJ�k=��2��=�G�M><�h<���<��/�)����n<.S�<6n<��<���<�^ǻ�C;� =���<�(=�iV���=�Z	��Y��r�U��=�;*佼aܼ�{,=�	_��g���!�=4Y=��y;���g��<�"��|��o�Bh�<I��;>�<t����}�<\%�����Z(�$�=�{��\��� 8=�S=F�1��)�<�Z�<������|����;�߼�C��8��<�-��^�=�^�<4G<=x9I��(�S��eû��<N=O]�<�"=�����25=�O�< �<�c�<���;o���OF��k0=����[׼S�+=MI=�=|�ڼ#Ր��C� U��]<���<p��_�i��< �꼫=���;��:���|��g=*�;%��~�����)�G%=��*R弸{���H<1�?�}u8�򘻼��,=)Fʼ�<KR�<�&;��&�<wHY��n<���G4=�E�c�A=;]�~2�����+��<�o���=��ER������`��>���+��6��<=����n<���LK����?�<��=�8;o�L=!��<��&=��E�C�=���Jm�<�C�����5�k�=��>=^��<��[��^G=5v�<A;�D�` I���;�g��#o����<?<_�R���=Qd}=r��<-���f��YW�<Z�<B�;����L8�M�=~��:�=Y��bs,��ȼG=��<�5<��A����U=��(��sh<ʵG�iV�Rt��g1<�S=L\���򯼘���$�;P���p�v�м�=��TN��@�j���(�<�N�<t�<JF���v�=/�=_��:� ˺�[8=��<�
	�#o�<��<~Y＀�G��-G=#倽�޻72z�=�m�0=c�0Y�R��<r���p-�)qZ���<tH%��ob=a��M���X�O��B�������1<8�2�Ӷ_=�<S���M<�2<�dϼ!,w����N���W��/=C ��G�9�>.K�Ǯ�=l�B=ȉ>�1V�����<.$=�N�2�:HnB����<#��< /�!�T�]i=o|���EɼY[P���]���`=�G�����<�:�<kּRmy�3:�<�db=�F���<��;?�<�W�<���<���<�q=�� �1�=yD��[�fe{��һ'򹼪��<���������<�JH=|Q����8�ap�'+{�%��<�p�<�S=��<;\=��f�J���<�G��	=d�==Ȧ<�ש<��L;�ܼ<P �<���<Gn1=���^=e[2�#�L����	�=g�	�PGB�R=b�<��#=���=�X<5��;K일X;k���<鉽�`%=ž����2=�۷���{��	������X��)��;&�����@=��=�<'�"=�:"�b�.��y=�7?��0��YF�;�;��/��<�s<{^ ��b�W=2�=��A�N���uO�<?1=���<j9I��Y<9rT=C��h=I�f�E��aZ��I6��Y���U=b����V��Ɠ<�m;�D >=��E=��R=�D7=D+��Z�8���<��/=W�7=w�0��<a	^�J�=Ó��������
=��"=��V�)�U=������;d��<�y�L�'���b�%T��96���=�F��y�<a�B�ټIo�<,V;*���Z=�V�<��Y���'=��=�7���n�)��<�I���P��oz��&� h=u�K=�Fe�Ć�~O!=f�V<���8��<,��_\:��׭� r=����{�\o����� �W�w�ټ<�O=��u��"���o�С�:�n��d��<�p��΃�-�M=0�*��<d<H��:V=���;��<�O�:�<׀��R�4�ʪw=��=Wo�<g(�<b���@�o�����0�^��<{U�;�U:=�p���x�<l�"��^�<�@��_?�]�B�5���$�<�`�;C��<�C=��a���<��1��^6=hŻv�~<i<B=���<d��	�<�%��.�6��OҼ6Z]��Co���#=p�6< ̘<
�<��<-o\���q�}=tp=e�,�wa=}#�h�O��6K='=7��u��ȿ�<I�:��c1��w�� ʼ��T�q�L�޼W�=�X��4��{:�;/ּ��<��ʻq0=�KN��5��9�k�\�=Ì�tm�:U���y�.<�Jm<�:e��
$�_Q��닼�]���弫�=�b<&����M��="��<���6-`���t��,�����<�&!��&�ǖ �����P�;�6=��2�$�C'�<�Î<2 ����c�#漹X�o�&��$=A3��L�?ש;"@Y�!�k�=�ҥ�~���=�kk��Z-=FF�Aj�!"1�gE 9�㚼�i��� ��o����|��2�ȻD��_�j��Q9��j#���Q�p|;_��=C�U�y=<WE=���*�#�z���s̘���0��<�T;��'���/��&�*�3�P,=;i���+��"B=h��7	=quC�`�c���&��W���;!��;�qO=ʉ��ŧ��<��<��9=1�7=:��<���<��`=J�2���<4��8��� =]V���M=c��_-�;5\1��~4�*�=}��GR�H�g�2U)<�79<f������EO���t�<ї6��.=��ѻ�('=)�<��=L�ݺ�~�8t���N���=�ڢ�-h�<�=R=F�o<�'�W`h��aW=���a,�����U��i�'=��i�lY�<%�����<��'��>��/��{���(=��<��0���T=�9��5ɩ�%X���p� �=]�F���b��X3o�M�;<�5=EjF���=��E��p=@�<:��	��żLT�9��;�?�<�j�<�*;S�]�S�<��X=ş������|�"�I=oI�;�7W=���<����<=��1�W��<֍�<���<�k=�.��簼u�E��n*%������<0n���}� O�</����Nc=H �;��0<��bWp<K�U��'j=��=x�����Z��#ݼ6	b�
vO=럋<��=ȣ�I�=��q��
<��<<���Yn����:�T@=r�o��c �,�:�:=[���%9��S�<6�[<��:p�j��I��;�<��=E�=����Ψ<�L=V�:
˨;T��=�I=j��<�K=;�<s�ƻ+��<�3<:l=7����J=�&0�D,���+��J�"����D4=���&�e�C���֔$=��<$d��C��I�<j=�XG�<��I�4�F�v��<���X#�<_I����㼏�S=��P�	���D	��B==�L��T�P���'<�a�2/�;��<$������iP�<>~3="`ۼ���<ŗ#�FK��мyM=A�+�4���i�<��=��E�Ӻ�=%���2�^2?���<~�<c��@�<�n�p�<,��O��;��T=xPQ=��<�#� ��<f$�<���<��/����<W���A���>T����:�TR�Ze�;��
��U�<7�K=�0Ժ�<�<�E��K�<���-<_^�>^�D����:F���cC�7|<]_q=�	��#k��44�~�D�qIR��n�<iuJ�C��ǋ�<V}=�-'="����=��a�����P=��Y=��A�n>:+�[<wp�<�Q=F���� =k@S=r�H���/=��K��m<��<й�F�%<���;1�G��*�<�9��N����!� y=_�D=H�<�<�{��Sh��e=�-�<`�=G <��0�>R]=k��9�3�D��;&�����j=�x1<q	�<5�H�9�=�/��^�B=�(���oU�<u;��<�w2=�Af�8��<��<�n<W&<�7:�˲���r�[��͙s9�{�<�Ku<��m=��vq��y<<n<i�\����0�<�3�<�Z�hsY�OQ��#�m<��:b�+=U.��\�T��/i��H<��!=e5<��<���+'���<X}�U�%�C�7��H#=0����<H�_�)~1�M��t� ��c�<� 5;`jǼLO��S�����$�̼H�E�zO�=R����漯�=;�V=�)?���7�A'�:�#=��
��ː�uQ><���q�<,L#=�=����`�/���Y~���m=�[	;�A_���=�]O�Vkn=�q�l��=�<F .��^��$�0�<?(��(a�cܼf���wn=ƻ�;`��&�!�!�����҂�<O�N�sB��G�v��=	iռӻ�sҰ<�/=�}����ۼu�=�C��`6=��;��$��0���r�pd&<P�=��˼��=�Yf��h"=8v6�-^?�#u'=����<��ܼ���;y�<��<�hƼ?2��<�<Up���u9=�J�<�(&<}��:0S�;��<[����&�#M<<����h�<U�c< ��t�7=5����U\�%R��*t�=�,%��=@��;xB�ح<%<���=�5�<�o0<� �z�g<�S�;�d�J�!��Wo=�q�<q.�<nTL=o�]=F,�4��$��ȉ4�+�m�4=I[���lf�ҏ��ۼ�n;�p��=�]�<z�;w@�ۤT=���ٵ��S���̼���<���${!=���O�S��G(�������������KP��0=t��\K9=�xP�-W��D*���=��A=��i�
P$���Z����<�I�V!=�}<C�P����<�BG�O��<�x�<�
k���㼻t=�'=�e�<ł���K=Oj�;eT��ԟ&���6��!=8> ��"N=�2K��=��<:YL=ʷD�.u<��C=��4=�H=q=��F=/��Ng8=��Ƽ(<E�U=�;\��+	��Nz��=�q?=E4��B��<�#=�-�<b`ü{nv��;c=A�/��얻\8�<�7��̎<�ƥ�4Χ<�'��f�<�#=����4�=�A=}�ټ�"���$=�=ji=BH���<�z��3蛼^�}<�~�1�6��+<l1�<ʟ4�W˷;P4���p<iU2��ё���{�هX����T�"�
2��A��\*;(����u�<e��<L<@�%�����c�5=�2�<���<~k�<��=Eɼ��ؼ|�;�%�<�5��S0=�u�<�{V=��<��;=��=�!"=�I��m$+��@.=�p=���<8Wa�d��=���5<@�<:BV=�I=��&��jM=,�f���r���μ���<�[^���<�^ɼ0�="9:=��<|��<��-=�S*��޼��=�¦<��a=�
ɼ�����=a�<����|�<��伭��������w=*8j�B&)��2�<�d�RL�A鸼EU�;��<(k���;�5=\�9�^y�����M=
�E��Q]��#{��۝���=��<��,�<c<���z����=��\=�f#=sk���_�S◼���<�SJ=w�(<���nD9�d�ͼ;e&�L��;%=*0=l6�<o7>����<�E���x�<h�Y<>`5=%P,��+=�v�!���<j =7cW=wK<=��B��c�</�μ��o=�e��*��</R2=�=��z<%BX�Ꟗ�L�=GH5=�z=��=%�=��z=�׹��j�U�M�����{�;}=�H���Bg����������Z�!��<1�<�ⰻ��8<��#�2�D=
�<Tͳ�2H���g�~�2��ȇ�	�i<v���=�<�=F�@=g-=�P���:=N�=ϰ�<��=bG������=&*;�s�<����P"�'�x�*o����<W�9��vm���<|��<��'=�`r<��Hp���y^<>v����;f��%p=�,�<Ȱ:<�S=�g$�}�5��V2= V�<���I�<��C�7�'��nX�h<�X�C��B	:��!s����<����?=2pP=�O����B<�J=Y����f��z-��>�<VY���q=��;�Φ�H�=]ɭ�����J=mtO�y�;U%5=r��p=/�/=[?!�j	���y:�9��y=������J=vq@=7�Л~���+=�I<#m�h=�r��췘<ҡ�<�M=\�ټ ��=�ɻ}�k�����S�7�S0=֘m��ɷ<Z���|�_�f��:=>�<1q~<��J��<|��<s����<O�d�$=Z;�<�s)�;~<�:[����ZNo�/4=���GC��]�;I�X�-f����tM�#%D���@=�Dd=c=N�#���<�#
�>Y�=�@�<)�e�ϊ�<⽝������C=[^=�П<OO�<i��X��IM<��h�V�<ţ@��������`�<�S9�3�S+=ӎA=�S;=�Nc=?����A��;8a=H��о��Z^C�K��<4:=��9=�	9�x�1=�V�<��_�Q0U����<_�4��H=�"��E�ك;��2�����5�[�4��¼`�5�A;0f_��a�=(~'=�D��5�<PEU��=D�;Y��<�+�<�F�<��~�J�7���t=[��<V�#����<��<J<_�d%�,�.=M;<�+=)�<�������$�a@+�X�6=:3i���=�@�;=(�=,�9ͫ=�׮<��{�nm��q�'=��;~�<���:�����<��ڼ��F��2a=�נ;��2�Qm�<K݁���=*�N�@�=ǈ=\~<��&�=��<�'�y�A��: ��=�A�I=&���[���	�����; W/<Փ"�r[]� ���-B=[�,=1V����=���;mͯ�B1"��;<<�&<������<h�:=�(����!=��-=]�T��<��L�< �Q;���1w:=�L�]󻌉;<��y6�;��=�jc;m�, P�}���D�u��m$=6p�=au�<j�/�`]1����<I)<��r��n3�TO�rd><T�����J=�	K�]�g;�9<��S=@��TG;���M/w=��X�Z=��<gx3���%�Hw�M�
�]��<g@��P�a<�K=Cjü�3���<U��<�i;��0�;`HZ�S7�<�x���
=t;�[�<ˮ<]ǁ�Ï��,��:�<�w\�����fG��2���<�6׼B�={�-��0��R�<��=\3�; ��<�@<�SE=�c|<�#�;��'=ֺ֮��xɀ9K�N<�(����<�'��>�������<��>=j-<8���&��<�YO�����@w�;&y�;�<WTW=�l=���=P_��q���)B��}7������úFc<�bz=l�<UAq=���Y�/�%k�<�z1�c,�<�W���C=Ix�KdV=������Q�l(�<2�n=�&�<N��s2�<�g&=;_O�6��<��X;�3�����ʉ��I��)z<�P<O�!��>��.����{���<ɿǼ𠡻���<����|?�m1�<�pܼJ#�<	V*=��W=6;���f�`��+�j���L=;�`��+T=%T�<݈�����<Fz�<\՜�� =�����b<9��\bz�=oB�X�;�[��}x<l�c=]���Z;��=)��� =�3(���(��_��sԺ<����<\k[=�'=��G�i�N�� ޺ϛF=����}^=����ގ[��s�"�$�YZ>�2�#<���� 	=��&�rJ�<,�����`���T��=�Y<.`U;iA��N3�<�!�<�f����"=�Kb�R<���⮼-�+�����d<��<��<���<���<vr <W^�<qU����23=/�<�G9���</%�<�G.<��Y�dFY��o�8���V��;�3j�?-=��;��<<�W�̓�;��Y����<(��&}=𘉽�;2K+<ȋ.�#Ѫ�r=�7�;Om=�T
;�_Q<��ռܯ=ԘJ=��E��I/=�"���P=��*<��jɐ���%��,.=0,K����<X[� uZ=�F��7=Q����3=5�=�|��t==�0q����;���I�%�6B=��E<��<	�o<�W<�V,���<�=��s�h8B�؀�<CW���?�H��<��=8�h=:xt��S=�p=4������D�#�ܼޙh=<�J��:=�SS=�If�id���H�<x�;*������Z���i����M=�����<˩��V��=�;Т�����s<#�5����[<���<��Ҽ�T�����0J_<i^Y<-C�;m`�:�	�p��:&������#=x��"��j= Jr=� =>\�;Qi���	꼙������r5h=�b=���r-�3u%����<��&;��l�u��O���=��1���t<��i<�p@�v&����;v�=��;{�1=WK�;Hp{=�� =����6=L��;v�g��<�"��̼N"=m�<X�<�sJ=�?=�ݼQ����;!?ԼG@ =�ϋ<�+����=�	�EV�Rk�<tOa���=��"=������y<��r�$�@���=V������C�(���9��"�#��;�n=�=�4=�11��F=i�*�M=3�K�l�t=�W==��<�\�|e�<�����`U<$2f;�t�Ҍ�1��<%h�zw)=�Fq:��<#<��;4k��j�}�B��&r�	�q��kA<i�G�1��A��<\=_ożW�=_nL�zm�;� =j��<�E��4I��'���G= :鼢3d=��:):<&�=�I:+���<D%�=�n��{E�<]/R=2��<��)����<��O=��\=_�<��v�NûK{=��<7�=��p�4���.<�$�<�\�=�O�0ug<�܏<3�N=� s=��2���<�ϡ;I�|����<�9�\�/���T��&��@4��N	<��V�h0!;�H=I���Ǽ<
�"�%=��S�"���<�����9�%f=ЩC=�)<�|���<+���\�='j
���<�M}j�z�w��]�0�Q��h0��[n<L>u���.��)=�Je<��=��#�;ށ<V�ż���=���<0�o���F�?����y<�\��:>=K>��/~c��`ͼ�ǿ�弳�l<�=4�\G� �8�{���B0<����i:O�K=��W�<l=�N����ʼ_�~����=�|<����`��6:{*��8�;=U�ؼ�0�<�ڻ<�ɜ<ƌ=��I=�܌�O8���}<��ϻ��6����y��<Y "�~����p8=&�E=f�м# =�R�lu�="3�<^��<`h༢7V;�`=��x�&ͼh��<!kz<�׀=�y��\�<;�=�|=�i���<��k<Q�H=|�=�y=�LC��<�흻�I�Qˋ�'!�<�Z�RK�:,�=s��Wl�;�<S,�����(?�9\�(�оK=;?�;�}e=��Z;2g= ���u���>��*=��!=C���H�<_د<�UR=G[�<S=��3�q�f��
w�k4=�8C=��ļE�����6=�F�<=�<�b�:�y=�M2��ή��I�<�����x�*g>���6=f�<T�;_�%<b�'=-*�<F�<!��0�=2:w=Os2�G�f<���<���<��=f���M�=�y�<M�k<5#�;�o�L�8�]"���<��Jn���a����C=!Ͻ;B�*���=���gm����0�ު"=�LN=iE���3���E�:4;�S;=ԥ;K�#=<����t��g��Ң����<�y��F�V<o�<+=���Pu8�w��DE�*��<4<(�F�9�os�=�u�����.�=�4=~����m�M<���m=<m��Xۼ�HP=�]=����3d6=H#-�F�<
}Լ��):��Ѽ�G���<a`�;��<=f�P:E�ӻ�]�ԦP�6r5<��<L�̼x6�%��sC�<^�<Rn�5ƃ�<q����(��,�<�OM��9���-<�~����<'��<�{�;��,<��i�P9=#�v�Y`����<래��2=01W<��e����c{�K��<���<0@='@=Is��������;ҠK�sf�<�a�<ml1=�;K�;�ͼ"`�<���<Y
���<N=���NG=]"���2��~�<��Y=(�j��U��<�aB�� �;tB/��M.=�VP=�5=QyK�-Q=X�H�?���ss�����K��<{���;�Jw=�&/=�7�<P�<hU�<W����vf�0Q=7��S[�����>L<3��<��;�꠼�ӌ��\�Ҍ/=�eU�҃��߁=��O=��@<�����u=�t=,�g��\�ڕ�<b=6��<��V�K=�<�֌�H�g���>��椼�4�e�v���{<�0���S<�\�<!�9�wo��H��Au=��ɻi�
��Q=Ei�4�@�[����<�r=bW���y':�l/�)33���S<{a�<�$B���b��Ι�����;R�ؼys;U�]�/ .=c'[�R2w�0���׼%=ʹ0=�Mn=<�=��¼M��;%YD=��;���N��/�f��<80=�BE<�|���Z��im<�<�:P<$�P={?��~� �� f;z�����-�[�<#��<u=��<|=N��1#=�f�<S�s<�t]=k�;č�N
���[�<rL�;[q�9��5=��]���yp==��<ؕ<��<���X��=n�4=m��Ck��wjC=�*�ap�0��<�<�w<֦�_W<�JK=!:��]p"�M �v�m��Q�9SE���p=4� <׮�<آ0���	��\�<Q�O��^��^8����4=9>�;q�;�1'�<��8=�\�<\���{�wA<�0���̡4=A���X(%���	=@�o;DH=�l�ɩ��B弉%=�׷<R׼��N���H=�[�<Oͼ`�&=��8=}�U<�L��ܱ���=��S�Cߣ��Y;�m,=3��w��}E�#<���<��4���<��˼�K=pH=1�=	�=;�!=�C�YR��,g�<`=^�g<2ؘ�-D˼��<4�F���U��%/=�g�;��<c���ӌ<2���$���;=�Af�l�s� �,=��U�����h��>��_�&<��a��KE����;�6H����,�6�ky�=g�u=�=�2<��<RW�<-E�<O�`<���<;� =`ґ;� �<UC�<��1���d=`����=�<�4w=��2=� ,<o��<I�=%j�<��<=%��I,��]��<���z�<�A =� ��=�-=��-K<ӏ�<��lҼ8��<�>
�G�3�KD���F��U�~=���<��'=�����L=`�P�-H=�D=�?<gFK����;WK�r� <�zA<ki=y&�;�A��Bw<P~�;Vհ�K*��A:>7<��+=��<��s��&<;T�<Ƴ���<�ˀ��2���S=���/�
���=$e�:%ԃ����<Q�"<VB�<��G��E<�����<�;�OӼ�!��D�<��N����\�y�s=N�Q=�	_�j�x=wp������	���G<��<`j&=S�8=6�M�����)<<�n;S�Q���<<��՝ݼp�<���z�^=�jV��`�޴�S�q�^�b<]�)��R=*@o�d��<�P5=����K끼9YT=�z
=x�㼝��<�}Z=Q�G���g�s=8<����8����HM�-;1�".�:�~Z��H=X��;�D�<c����L=��<|�4=��*=`M=�����0S=���_p=�j������;�<��ļ��/=���<a%�<JGE�>R=`�<<R��<S '=����ΆI����8�S�J\޼�
>�I���^=��&=s\�d="���B=�P=��
��H���
[�t���K$�!��;}+=������;[��<!�8<=O�8=�.���a<�z��󖡼�?d�T����kq<��4��M�<ǲ�E���KOd���;r�-=H�<l*�<;��x�<:A���U=����<���<�\=4�9���<cB�<}��xq"=�0�=�h���?=Id�;��H[6=�x=�PY��)=��/�6{)��V��
8��Vo=��Q��I(=|��9��s�]<���:�W.���ɼ7��<���<�)6=&U���J����<΂=5�$�{[�<z�O���\�>��<�UD�?�r=���q���8�i޼���<�]ź?-����U�$=v��{��<R ,��v�;���}"�:�$=��\<#�8=��C���F�T�?S��'�<B2=�� �\��R����;gQ���i=�����;�P=-�����<�<�����S=�a=o��BF�V�=��=��	��e(�p �"��2�����<E?���L2<�~;��� =�	V<�%/=�P��@�(�O<I��<�//�N���U=~C�<o�W�t<��)�� B<=DG��Ѽ�K<��l=k�/=�V
=�揻'�<�Kz<�4=&��;ϔ�<�wϼ�2:�p�;��<O�%�/Q=��&=��<{B�<��Q��0��l=�]=�J=d��.�����@��_���z�;�f�<��<w������<W	��v�#=��X=nμ�Д�g3=K�~�2�m=�ΐ�l1���$=�$S���AT��j����</$0=&��<d1k=k��LDL�9�G�G�������;��=��ܼ�^��H��;�s;=ռ�l�<��9vd�CJ<�x���������<]t��7m7������<��+����<&�<;���3��<��2��h����<�y_��,J�	Pϼ�yD�%�S=�U�<�:G=��M�VE<��;���<�#���T<f-<�{�<�x/;ߟ���N�<�B��Ahn<�"=<��F��<�c�����<Q0�;�*=^*=���<��^=�4b��40<�p��<�W��`.�+�ռ�Q`�!��;c=�&B�_f��@黬IO=�D�<�Y=� ,�dI<#�2���&��ƥ<TȠ<]8�=Z�=��=�:[�#���sC��5P<��;5�<Tqk=Ve2�?0=^�g�({�<�o�<AC����=�>
=�y��Kb_��ۼ?t��'Rؼ@�O=2�=�==�/E;rX�<5+8=��.��v�<đ+=����y�����W�T%!���[9��_!�	'$��;<��ۼ���;� <��A=5>=���<��3=��;�p=�H<����N��U=>�;M�<�<�	<�P?=�Щ<s��<�K���=<XԎ��P�(˖�D�r<-���7,=L���:��<�=�q�<���<_k=���\�*�cK��q<c��<��2�9�[=
�T�xһ�޼�=x^�k,="�W��H�<G0��;<W٨;�d��MZ8��[n�8LB��n��ގ4=G}�;y�=�d[=��~<�����U�a�����ݻ����lt�-Jl=�	�b��<i�H=��߼|��<�殼��:"z(=�		=�:<s�N=Y�b=0M�;i�Q�n�=�V<]�C<qx"���#=��=���Rm�:�1�<�V=��ix�;FD��
��ͨ�
?���Y<s��!��hh�<y*�:�E�N9��J=�"���})=#�l<�$�<yTZ<�^�����Gh=3~�<_Eo<��<�K+=V*'���<�n=�-=� ����:����Υ�9!�-<���<+3;=F^h��U�J�e��YL=��O=P�=��E=�O���a�<�V��M��<�K�C%6��Q�k�<nG������%=��+��E�=��O=���x=f\*�k�<�%9PA�8nG=��:�}��d��<!sܻ�M3��΀�}�=g��<��7<MD�<��Q���=����X��^J���~=�蚼ۮ�;��L<���y�R�|�9�6#=�ݜ<�S�Ti�<�����^�<����I=(v�a��;�^��$�O,m�.�	<�1�/��{=V>B=Z�|��`<�c<-nλ��d�{M=�=B�i�x�I=�x<�7���=M=��Z�p�5<Ap�B6L�h�<.FL�#�A��#���/<ڼ���������L�<Ŋ���jݼmfW=���<��޼����c�0��d=oO=��p=rܾ<���<�H��0B�m��L�z�U��W�0=||�<,���������#�U���I|�1�=��b��-�<}C�<8Y�<��#�Χ'�(s=4�*����<��$=��$<�2�.ß�A�<K�y�$m�<]p�;�ɷ<�y���=�L�<K��<J�<>�e=B��������i<�xM;�y<8�ܼ�u��=ȼ~�<(��<��=� �;�9<��;=��[=�����=&�=�=нI=��3�<��<��<F� =���;��V���C=�:����O�j��>�<��=��G=��r�
�e<J@�c�F��c�:�����&;G��0xP�%��<dw�<n������h��p3=:N#���<lj<g��<U=(=�X�<��e<��Ż�購�F7=��������2�6�<��L�2�=k�T<�%�G�L�-_=4�<k�<y�V=^���:�<EY�<��-���Ѽ��K=Ȫ<�k<-�<U�Ҽ�|=טj���?���`=�5��&v0=�6=���h�D�1=i�!<���<d�=�y�<��	�>�Ȼ�_�/�<��r=�[�9).=������6����;.�L=�^=�G5=��P<��=Y�<<�<q����=����e�<�B�:'��<c0U�x�;���b;��;�
)=��ռM��;��"��L=#mļ~*�w�/=x��;�<���(>A����m��?<�=ȲW=�����<̉�� �-;���<ޫ9=0� �[�Y=]qڼ����yq�"�T=0�U�Ɗ�<�<~�g�)�|=�+��UW<h�6=�=w*<��U7=�=�	W��Μ;��#��^J<[m�<xr<�;Ӽ4�z�w����<;N
���_��3�8Jzü���-9����<dG='g=�����=�Q��^��<	����;��f;� �߄�Bc�;E�6=i�]=�(c<�<=�	=!��F�<-1h�"I<<p���\�����r'=.<��R=������<�{Z<�K=Ɖ]�ī�g�ڼ:+���_�<Ă=��;�ɼ�4<���DR����;"=H�K���&�\�׻D�]����<Ȇ��b�<��Q�݁�;����
e�B�P=�*����<)��2��ğ���XQ��`=s8V�RU=�i�ٹ��3���<�/O���h�3-�)�o�WJ������[Ǻ��G�J=�Sy���
=�p�<�/��:Ɏ�=���G�=�!1��C̻h��]-=<�=[����ɥ�j=����q�@�E4ż�?�< �<‼��s��x$�;�����<ߵ�;��Q=X�ټ�f�y�</K�>G=��}=a�,��A�*��<�����0:����|�!=�-\�7��;ؼ�]�=Լ)��_],�����<��=�������[O=� �<qi����\<�)S=�i==�N='=Լ�^W���F<��5�<<U�o<��&:\�+��껂�W��K<�-4��ة�;E���p<"<��8&�<�������;������ɼ�j4=�G;jE�<>�3�ܚ|;���<�-<�
 .��Iؼ�I.�>��U��<깆=�0�=蜄�O�g(�<�(�ސ�<���;�_'�%(><��B���5=�n�<�Z<S�A�Wc��R<�{�<?j�u�r�@l(=�
�<��1<T��<��<m��<���U���o<2�k|=n	�;0)=n�ؾ=�.8=��μ�f=��"��-�<��_<j�缛=�>����<'x�<���;��ݼp������iT�����W���;��<��˼�rw�t�=0m�+����&T;�=�b���̼��м�\<�=a����|�=�Bk<q\����͡����n���<K�<l�v<���<}L��=���;�<��b=�� �*�<!�r<Tn�<xe4=-_��������@@Z��#���Ѻ<�󕻞�V����=��_s�<Qżvl��@O
��GV������`<��<���9&��e���,�#x�<��ݼVH=�}�<�ٙ���C=~��; ��;�μ�
=���:h�<54�<>'>=$E=m��(��F����X���c�B���,0=�3=Ն�s�N:��U���:�:*=��O<��H��/?=5��<?a=�oX���M=�[=x��<��T���X=�;!:]� �<�߼ben=��<\�*=�U��m�<7Wd���F�w�&=�<���׼��<�ꑼ&<��+=���=���� � =���a4
=��9D���wK=�l=s=�����8"�ѼQhh=�@<>�d��güc�L���Q������m�<t\K���7(���?��C6�?O�=ݟu�ڠ:��j��I�2,���h�=aW*=� �W�<J0=���=�=)@w=���B����;{[��e[b=G��=%�T<d��`�컑<�<�.����/=aC�<�L=g�D�;�#=��h=��.=z��pNO��9��nͼn�)�M�i=�W� �I=	�"=5�e��̌���¹�t�;����S1� �9�s�=�F=t�<J:��r<=9(i6�2O��J(=>3=F{��BB���<=i4��Mv����<#�w����m�&�_�<��8<<@`��G��:(=�=�\��	��iy=�B�;�e=A��G����<���;OU9�ٶ���~����;vqj=���ơ��M%=�3Z����H��Q��y��<�FE=�A\=�Ｑ���C����=�R=H�n��z�j�5=X3"���=�03���'=��< �7< 2��al=��T<�\8�?�Y��~<�������g=�'��b"�<�H��>��<�A��i��m��;�)����<L�G���<��<2�N�b=!�E�k��<��t�[�����u��{�;�1C=Q�<������<��K=@�'��X��$=CN�����%��bI�R==����&��䃗<j��;���F7=�j�a�t=��4=���8��<K�+=��<j"����<��:��?9�(<�A&=w�;Z��<I��<�z�G�<<��<"&k=3�7=��=��:�~A����'_�<�b5��S
��p �h�^<�R=u�<�J=���51=�#q=�9=�%;<�^��㼴���9��nB������[
��"��_����an<^�ͼ�7l���=�8�켤�A����<�Ĉ�4q=���;�q��������<�����P�;��ڻ#�&<����E�����o�;O{ɺyaY�~p�<���<'pW=�o<��M=��C�b8	��t.=��v����X�R=���981����<gW�<�:!�q�����;R<�qj�0T�<x�h�Qtȼ��/=ޤ�<C�=�e�<��<;�;��ڼ����'�<��=W�4�����J0�<C�<d1���e��cu����<?��r޼er�0�F��3q�Q��<�j(�rb=gK�UCq�#�<	tW=�D��/��;�����B��<��Z=�O#=����S��N��;!��:�{�)�<�E6=q�Q��,�(���r =��8��ފ=�Y���ټ�ʘ<��Ƽs�D�
;���}��/ӻ.L��^=Y�"<A�t�&�'�c=�E�<J�-=�Ɔ��=���<�3;��3�<a|V=�d=��=y�<��
=�(���g���=���<��$=RPY�[�弮��<�ê<�ۥ�z�<E��<ĳ3=��G=��b=uE��[w�<���� �fR<@/�<��`<^M��l��^��;�Q`��fn=ƏμnL<=d�"�[I ���;�Dۼ���<��<;xlG=])�<7G��H˼g�=<o�<`M�ʝ�ƀ�;��ǻ�V�<��z�<<ӓH�!�f�,!�y�Y�9Є�f����c=�U=\�<�&d��W�<� =I�4=����@���7���8�<F찼2$�<�'=8�R=�K���Z�#.��3�!=���$�m�ͼP��Zp}<M����n$<�tL��)"�j=o:A<�������]
��'�;�==E�<�D�l�=b���0=��m���=��<i[�;	�u:�Q�'�3��h��l|�����WXO���M���-���м&��;
 2�#�	�k׳<�I���vV�r Q=Y~�RB�<V��G���p[=Ȁ�m.1=
a��e���q/=�"�Ѽ~n��z������u1V=<���/y=��<��ʻ(m�=�+P��u�`o6=��<=s�k����;鎂���6��;�<���;o�ڼ��<�	�]ɂ�9�I�y�M<�Q���/=;�+<% �̈�<E�<��S��V�:�K�@�(��_9���ú��U<̒Q<g�	=
s�{�(��+Z��t�;��캺�N��L��9*�<{��;�n:�`'@=\R�=���5�<��}��+u�������<;�<���*�<[!����߻�bȻ��J<�PQ<f�:�v�F/���G=�OU��w���^�\@(����R:�<�=�tk�<�^�;�qc;�'�<c����[�C=�R��4I=�<����(�f����oG	=rf=`q�j6ǻh�<Z�=�E<���;�k�<����z=�s9e�ڼ�l���<����k<���thw�UQ=J7�<��<u��<�\���J�i�=Q�Q��䢼�=�<:���$�ii���S�;{�;<��k=~�V=���B��m.����<�ḼGH���!�<���^�;�(H�EDL=-M=���<����ͼ���<�k,�ˉ9�0�-��I�<x�7=ɵ=��;�w���I�<(�f���Y���C=�T�;f�;��������U�<��< ,��X�1<�Q�J�
=��:=b�#=�4��gnc=�m��|=��ʧ��"ռ�iR<$�,:�(ü�|Լ1��g�\<��
��+�;�
�
=�<�Ӿ�G^8=�N�<�h|=Sr�ZL	=�Z=�!}�C戼�F4=�⺼B�=g��<EL���ؼKQ~=���3X���e���p=�1�?��<��λ�/��k�'=�H�;�h=��؊.<x������5��/_��0��_B��b���~�
D=j�k�c�1=l,��n�
��ʼ��=�=��#� =�< (�<�=��<jj���617=�bF<�7=i}1�
�༾�&<��<l�=��g=��\<�o���/�<7x���&���A�tms�,��3���H�<@N3����t�t�n=L:�P� �,φ��Yj<��<�E=��=�`U��\�<j���s�a=M6=K0"=
��<8�=&=I=�#=�\ڼ!7���Gw�Gڭ������	��?=��)�<�/���i=wJ�<1��<Ɨɼ������<^-=�<�=���<]"���,��\�<S�!=O�X�T;uk�<;��9ټ،;c��~�~�H<�JE=�kO=Qֹ<5��<l�������iɻdq˺'R��-�X�7=Y����iʼ��-=�^/=����=b�:���<�J�<���$<TR#=�������%�F��;�ȴ0=��<��[�� :<�J���Z;����}����;��;=|;��>=͜M��+=�*���XI��j�<��	�l�3�Y�W���%�����6<<׎���L=E?<��9�D�}<SZ$�ݷ,==�!;>�`�� L=2=�;��4=F3��3�;s=�������u=�i���^���]=`X�<���V�;�6��.�,�4�T��mZ;��;N5˼�ٴ<��.����<Z=4�D��f��ð�z��<���Z��=1��:@�ZI6="'?��}�=^RۼdF�����%=��m=� v��+N�V.�-("�Z� �P �;7�<fa;9P=-�D��H��=�̹�˛��ۼi�<1n��gj2=��ü�D���SX<^0:O�5�ʣI���2='���+������<�T�<�~�\�
=�7k�-�c��h_<�j,�$J��=�e���Ƽ�� =�02=���;U=�4<���ly=�R��}�s���3<��C<%=�_�?�=�)��88j<U�ѹ;H~<Y\��� r�9����F<	6k=��A�����!=�7�<�:]j==&^=@�=۳�<Gp<��3��2R�O��<Y]�$J��P�<J�<<�🼫�r��
ּ�U=Jk5��:��=�D`A���I���y������*y���-==�K-�$��^9;�L)=�-�;	.=z* �?�0=>$��8��hf=�;��=D��<�==�0�����>���m�R=o�>;��<r��<�>C=�>=}E�<�D��t�;z�)��9�Ep�z����Ϥ;��E<�;���V�<8Y�<��~<��'��#��N<��=�q�;u�>9>=N��;��E��]=�p=��=�`�<a��<�o� F=ͩ;̽����x��/��Y&�Қ�quD<�&b�Cy��'<3S=X޹��5a���~=q<"=3=�ih=e<�A#1�«�<V�Ƽm,=��	=lj=L�<1>.���a�wd��ߌ���L���-e��W=Sp=�^���N�)��<�7=�1A=w�Ǽ�u�<nwC=T.���\<��"�,M=�HG=���<��<�A=
t�<=!V��<K L�h����<J=�1�b�C��.�<M�;=|�<�=��/��M'�$=M�,=~45��9A=_nƼ�e`��-=Iwg=��G={{�����oe��ѹ�'P2<�S=�.ټ~aD��_���;��/=@��������K�<R��6z�=�J=d�J=�+�<:T;��<;D<��;μ>�=�8�<H�=��j;A)�~ �<<+	=�f��-b<�&O=�O>�V'<�vμ��7=%�Q���˻�1�����}(U=Ǟ�Ƃ�<�lk<�z�ڥ
��b��:n�p�^��@�C)=a#=�@�j��h�g��p����3�μ�r��eG$;�=���;�
�</d=xT��ۤ�;�� ����|���?�w*���?�<;�<�P�;�9�: �9=�?�;*Lc��p>=D=����:�=H<�t�<X�G=G�c<}���==?]x��>"����4h-����<���0�<1�<���<�?1<�F=�N�O9'���<|��.#=�G���"���=��Q�G"�4�=
�:�B�`K��
����9�:�e��h=�Z=�E=��C<\�;�V<v��;{�5�]����a;1���;=���<9�^=�}e=o�ݻ5�K�#���'=�]T=�ݼ+�X���=��<䂘;e��<n�*��۾;��1=`��<Ħ�;.}^<	(<��*��%�$�f<#i�<p2̼وƼP���]�=�m���	=��s�0����e�z�<��]8�ϲ==��3dﻎ

��b^<�ݙ<Ԥ=�mX=Z�ļ���<�P�=	�	����g�<`�<:Ƕ;kq�<�u<]X*=n���xYx=�zS���<d-�q:� =^�:T:�↌=���<��):�Ww���s�&S�t�)<��G�	P���3��$�<,*=%p=I�<O4���<��<��D��?I�:��<�p����$<~1�<�B�<��i�43�J��%%U;x�D=N���=��P���w=N�a��W��2p�#i���Y�B!=��=G8=O���/:J:g=g'd��j�<����{�<F�1�����=��{=�ҝ��D=T�ȼO�Ҽ}�'��;F=%+μ�uq=/J����½���S<�֒�	����<K=�̾�̱C=�t�<ֹ%:*=�i!��C=;N,=�~��_��T�ٙ�< �D=��^=�'=?T=,�D=E�n���������ȼ��_��|Q���_=�5==�9���r*�?��<��̻�e���<��=����V��\=���<wc����b�[����ż)ZԼ_�$����R��ƫ�ӛ"=:K�$o2��r	=\�<�[�'i󼙔>���<���d%��¾;�������=@R@=A����-�`2�AM��� �	�����;�%ô��	�P�=B =eF^�C7���Z�-�|<���C]=\"�:=Y��/_�<��<�{�<�g��<g㞼r�K�&��B����;��5�]���*�I=��<EGb<�;(=r��W�=���<��=_��<]	��������ټF
*=��H<Z�f��:���=b9Q�S� =�I��7�?��_��Q�;��P�	���	���F��CG@=�GX<Rћ;'��B>Y<��r@�=X��5h<4V���+$:Tg{<�w�v�X�����f=&�+���=�0=ࣂ=X8)��Q4=��<P<�I*��E�<d_��fd��y�B�EP����������U�"yA��D�${��v=�s�W�]=/��J&=���<�����Y�v�=��"=�)�=ܝ�<\�ڼ¯����<�K-=xDX<�U��a<{��<��<�Tg<AlB��/=jV��Œy�}�w�'=��p�fP�<�jd��"�<t	=��<�Z=�q����<u�
��s�TԆ��p�/n�}W-���������H�����!7�<��7=�5�=�f�I\$�
:=Ѯﻅ����@=�j=j
;��M=����%��`�<	�����=\�=7�8=��=��{�m�]=��y�ɫ�<В����;�x�<�\!<�e<�n�_=�H"=P�ȉ.=�[=�AҼ�?=�p��ď��:�)<��U=�<���;�j�'!��U=���<�2�<� �;&t˼��p<�O�<��z��o�Yf���F�;�~�
�e� ='��<�u�<>Ea=��y=��9=<�=�07��5b=e�R=�5�67=e��<.~�&�"<=�q<dD|=G��<a�6��)ںP��<.�'d�[7ͻn�j=��@L�<������Kj<25y;wOs=j��<�Z��ćC=Y�;<��'=�4:6���k<r�u��<��˼�����D����=�ˍ���1�e�w;lم�g��= =G�2=EjϺ�B�;�Z��m�^=�:Y=�*K=xJ�a���x��ߩ��I=&N�<�+�sj2���<uJ�\ Ǽ��@�{�&�!�*:oR�|+!=J멻=I�<����N��+h�3���Jp»v�;����=�gۼ�Q<����X���5�C�;�Ő�=��̼#V��A�;��b;��`�-X����<�=8=�2>=���Vj����w��������T�0��<�$=��\=�X=�^o�x����8�u<��<�B���w=�iP���=�.���=^�-�q2/��7=�U�<\-=��=nھ�?)��t%��|�<�,�� ��<��ݼ��*= V��@���,��.9�� ����n���YQ!��������L+~�M�B�&����B<��A=�׺p��O���Ļ �ͻ�xO�<�O�3s$��@�>Kb��qe���=v���1�<�SN���^<��</�C�Tx =���|Q?<~��3/=�����<-\L=F�G�ho�<�P<N"�<�ل�`�@�F��<E�<�W=�rv=�H<L�}�,_;���N�:�X=�M�<�[��7�ͻ|�"=�!��&�\��"K=��=�y=�瓼�r.8(��A=��Z<��<=��?=�4=@J1=��<PL3=f�$=01= �ź���˴�R<=�֋�t]��*a�E8
<eiZ=Hs�<�r�`o=����{��<��T+��B�;$lT����������s�R���E<X��^נ�'[ڼp��? )�&vR�Tp[;^"�UJ�*V�=Լ�֖<�ms=�8=�Lv=O�ϸ"="�i�u)'=�Y=b�{�
�=��=T	����	)T<�<�<��u�:y����n<ܻ�xG��L���d*=����t��\�����Ǽ�O�<TY�<k:=��=�u=��`��d<��F�%~N�h{=�07=0�'�E{P=��<W�p�t���Z�Y���<i��<��<�Fa=y$�<�!�����Yٻad=� ��n=�T��/0���*�_rl�F<�o����7�<�Ǒ<�}Z����	O=��5=�����;�(;*�`�'j���F=�<��<v�g�� �<��-��<�P;��I�G��<�2����^=�-�<�/=��+=��=[}�<��H<�E�e_���\=A��<��<���}��<w�=��;��>�v���$�)=��"�Z�=+Xo=�O�����<{�/�v�(=)�A�lR��A�;6?����;���<#�<T)�=|�i=l@�<����I�ܼ�k^�q{�<�94�>��;^�U���Ҽ���<��@�c�<���<}��<�>�;zv=�>�<�Lu��Y#=�Yp=�5�<����[����̼�Q��>	=�<$��8a<qxC��`ܼE=�V��輅W/=�'ջ�䲼X]��/~�;a2���h�vc2=��뼒��<���<g�߼⥣�WeY���<Z�9�q�O=]���7���zM���2 �M���@���"Y�4[���{<���<d�F��@B�#5=j1M=�#h<P��1��;�!�<����/�<90�;����ku�<��=&3�<��0�u�d�(�(=*8�p�<B�vJ =��)�	��� �h�D�3��7�<�o<���H��<B<ἡ�&=�+y=;��<��'=�Mj=����\=;�мA�<�)<������;�y	��`��%?�4��;�P�����<�Ζ�B�==��Ի=D�<}��<G�5=,&�ѽH=TJ�;ti��?�<�P����y���R�ӻ�h��=�=@�H=dT=�N=�=�����iP�a10�U(U=ɮջ�f;=��=H��<V7c���<|�T=K���~�;?�<	�<'��;�I<��D��Y�"A>���Y=�t�����`�*=�2$���4��/=�K�����v�����<i�<=X-�0����=���:[k�<��<;��<�H]�Uq����5=���9�T%=�8!=؛����<�cܼ���#���U95>=A���p�z<wɊ=�}Z=yY<�~=(�� ��ޙ�YiH�p�<�<�I�fu<� ?=]|�<f<��5��;�=@bd�cT'��=�����E��:<�5?��vU�K3��X�=�+�W��_k$=���=��u=Es�<*Qb��?�<���<jU��ƪ��:�<�<?�u�����W=}�=�b�����<ɌH�M]]<P�\��<�ǯ<�Yr=G�X=�	��x*�OQ_<��O=e<��xԭ���O���6=m}z����<.�I;��R=�̻� E;�t8=G⍻!_�r�׻?����=�1Rռ���<����^<�ܼ��?P�D���==����V,;�Հ���㼕�\�q��2I=kX+=��C=��9<+�;���G����&���,�<�~ =��<r�����q��	���2��j:�����#�m�|�bPn=���<�<L3�<4=Z.{;�E=R-=�$=�t<&9!=��?�"�;���<�����,���?��!=f T�ϡU��_�<R֖=�f5=��>=3l6���E;���C����>Q�7nB=|]�<�:�ual;�w�;
�P��nX����<X�<'ط��QJ���e�>J�ۇG�q[ ��U<t�m����緯�Z�Ƽ�C����>=սb<�1u=�IR=�ɶ<;KW���0�_>=�ړ���i���D=��{����X�íI��p�<�Uh����<���s
��Fh���=��&=g�B={7���<��4="�n=�A<]����p񼧗5�TJ���O�;�nY=O�q����-]=�K:Q��E,�;w��o&��v�Vw�z�[�{�;�:=��=֗����Z�}	��m�0=�c$<�q�D����=ĸ�<��m�\7�֒�<��9<�­<S틼�H�<�%�k�
�&��uz:=�V��3�=1;>�=tҐ<������м�8^�.)��UD��E`<(�=T@v�ZE"��=D�r<@��<�-v�>�F��4=P.=�
w��'��켓QF=��(<�f� g"� =���<��;=�Lڼ����d��TG=եݹ7�f;@��<��b�/��<���<��n�w�<�p��Q=���B�;!:N=K�:#r�<YO1��2.�VU��=P��<M9=��<ѩ></qͼ_Y���<��D�+9�U���`痼�"�%�=�(�<�<�(���c�����=�!h�I�>|��E =i��;� �<C�P={H�� �<3W��ύ����q����;�=-����=���1)������<ev�<(]=<��;Z�=�ջ��E=�&.9 R�䜀<J��]�<E�;9ac� :�<]���_b�� +��X��!6��Tn�j~�<Ee����N5��B�8�2�c��!E<ю	�܀�<�ͼ7!��S�4J�<.!R�~c<Z꼺�,=���9�<��"��B�4�=�p�<�6-���6c�<��L=�m=��+���<���W:K��U9<��5<�S�Sc3���ż�<6��<���;��,��,��D���3⹼��h=<N�ml'�O�-<$�:�μ�V@�+;LB��t�[=�x0��Ѽ�"<�=��P�]a-����A�%�_�q�&<t��Х�<��ݼ�Z<Ť8����<��C=�z�<g�Y<��<��5���%�iE]=K�l=���k=�+������4��<�?`=󘇼��:���=�?�<-4=R��"���.����CR=F��<G܆;�聼�e=�^��S=�ν���=��r�%;(=���<��=2�#�<YUмz}(=�L<���<��%=TP<�OP���#�C=��=W�u�4��<�A<:>RD=�뼇�*=�8�%L��|�L=���!X�;��<�t�ڍ��)<	c��Ay�����e�<4�O=��E=��<�?�rn<�G�<�0<xR2��U�<�}Ż�1��^�<ih�<A{�<^�<��i<�]���<u9=e�<j�Y��_�j��kR_��^=kJC<v��<�I��DJ=��A�0�̼���;\�ռ� ��vU��_=�P:��K�<���fZ<�Y=B}���;��:����I���=�)<�PS����;L��<�?�"�]����*���@��n���N��<�?�;�t;���<��к�L��i�������K<l��<�EL���<+�k=�nϼ�l���v�<C�8=�4�*�"���C�fh=gb
=�a=1=���<���<�pڻ������Y==wa�����̵�b��w���f�<>F=X��5�<�6�<�3���!O=ONh���=�m�=���<M�7��#�ڥ<g���m<C��<򈌺H��~�꼿F;X�$��sn=���;˜�<j�^��09<!S���3=D�=W��%�X;���<\���³/��W%���м��<�����E<�嬼��ϼr�z=E���sJ�<G��=��;k|�q�s�:Zü��=95�u(f=�����h���$�畴�5�!���a��LT�@��<��<�o=��@�O��;S��Z4]�z)=	���F�������\=|P��B�1?== 7����ǻ2M�;��� ��<�.�<�E;��~ܼVh'=~�=�H�,��|0�:o.;�7R;��ʼM2�w;4=��;�p�a*=����V��9�_^�&T���9�]��<,뼍9�*�c<�΁��M�%� �FК<����ձ�9F�3=�K=��
=Se=<3ż��ۼZ�.=}��=��L�/؝�B�:�;�;D���������d5=cL/��g3���6���p�D}h;�'�#�)=�N$= ����K=�'z=�n&�WF�<BTٺLa];#��<"=E�9=��=�W<=[�="�J�ݰ�<T����|=��#�T�b=p ��uNX<zQb�;+X��Un�l��=�ѭ<�P*��A=��Z�!;D�>8a<Jzj��v �vO��,2<8���y4�1�1��8^��=N)¼h�����V��X��v�~<�u"=3�%�w;'�U<�|�=�"����A���]=��=�*�1��x-�N��==($��	�;�*���Rz�<��t�V��<��"��9��^BG��W@<Z̅<p=u��<MPK<�Z��S=K%��O=��ż�}���<�X��a�<��<�w�A=���|+_��P�<�P��%�1�h�U;F=4�.�דl=$7�<!���s+=._O�	�X=S����2�;&�l�s�1���<DF�<��_=��Y=��M='�*�Zf+��&�Ku�<:hc����<�ͭ;�%e���Z=}(=�C8�܄a=���x�*����4��<��<Q����CH=a_T=��<S�9cx�jgS=ŶG=���y��<\�N��o�]�1�J�*<y��V�i<�=�<��#= �c�W�/=���<�N=�7=jƝ�<�,�`=Q�����D<N�_��� =��=Qv<=��=ڠ�<#􋽣}�2"=,-�<)�
��S��<�j,=��A��̪���j��<@�K���L=��V=^�=4)��ʻ��ټ�꿼9k��^��<Y>;) �����<�J=�=x�ڻ45G���غ��<�52=�@H=d�	=__��@��<`��<�$m=�%N����<u[c�a����v�;�ּUc�<��i���<�Q�������T��i����6=�����<k�K��{��Y7=}=����E��}8S�^��4�]�%h<�2F��Y<S2a<�~t<Ȥ�<_e��t��<G�ZHe<-�H=-��;W�Ǽ���ש#<l�/�l*'�T1<��3���=� 8=��k�TT?=�=5<H��uJ���=��=�I�;<0�p�ּ-[�8���8	�<*F�<X��g=0�H=��.��F�<��<�
�Fԏ<4^�^�
��A=���<eڝ<��OhE�3=yK�Ԇ=�^x;�xX=���<�$�<�I�#����;��K=�{���Q=���<�md�����\M�����<�����3��#f��=���e�=`%���`[=�?�G�< �e:RL��pK<H��<�5;B2�<�o<���x���n:��̺-qu<�2=�6<��ʻ􄽀���KQ=�vJ��0K=�x�:j�U�N�&�]G=��a�;��<"�U=���<&^� +%��%ۻN �<H�<�\��g)�az�<��=_� =�4��.Ѽ�c�<��ļ�=���i���=���<Sd<X�������0����٣�<�7���O=��1==\��(�:��պsR�<M"�<(:�G��<.��X	H�a��<�μ�f�<��';�&׼@P"=��M���<�H\��LY=	�Q�� �����4<DQ����J��;��H�w�<��]�<l�G=�*=��U'ټs|D=�[��Y��<��=�m��~\=⮇����ռ�46=S�	�����V,�6�!�E�L="�=TMڻ�e���<+rm=�ݼ��(=8�������v =� �<Ù<G�H��H*=��^<4S�;�S�^�<��=���<kt��V=�Ȼj�漕��@v�<�@A=�T����ʻ4@}�W.ʼ��;�/Պ��/V�4�<OCb=�(o�Ff_<�k�<�jl���ڼ��<�wY<ED��Z�=�;��V��Q������߼���?	<]�B=��o=�ֻl$=3�ؼ��<a�E=�W�ɤ;�3���n˼��!��rq=z��<�,6=c���y����<�lռf#�;3��m&=V�I=J�B� 
1=-C׼�5M=8�v��=K[w�2,��&���'Ҽ�;m=ѐ$��<�;#\�WN=q\�@��<w{ ����=�j���%q�q��<w�
=-M;���A��<�S�?Q=��|�x����q���O5�C�=����6	=�a<:)A�.x����;��I���	<��=�{ݺ��<���<g�<w���c�<�2$=�d(����;�hK�a���Y%e=�&��ܯ�����<��<\sL�TuV=�w�GU��ϭr;��r��햼�PT��=`"�i`�:̄���
�<�$E=���<-o�<fh�������KJ����/��<�C�<�<HZ�_0�<��D= >I���=��H<��ۻ�s5�keQ�!o=U{�yB�<�	�+�#�rTP=�-�<��<#A�<���<��k���л@��T�</�z=O�ۼ޳D���v;F�P=��^��w� ����ͻ���<�V;���S�R�v�N=C/X=��=J����ͼ�ֹ�/d�<x�D���/���C=8R��\�;o\<8�_<'у���<�4�F==�:���Q=yf
=�޼'�&��N��P;<��<�|CǼ���<����ß��0=��S��t<:1�&=�N��ϻ=:<�����l��;��<�Ѓ��͵<���<�즼�wa=Trd��(=�D=�U=~�A��)q={<)��ؑ�������(�-�S=.��E�.��}��.L=`G�aA
��`�:Vݼ�%���>���μ�)6����< k�(�
=��T�e�D=t�u=r5żW�%��]|�FQu����<���=�D��ZC.<!����`�;�w/�&=�����<������<�J=	&�����;�<��<�����n<��:�+d��!i=Ե;<ᙀ� [Z��=T���V��4�l=]ݼw��=��|�8�MC�ф����b�ߩ=0O3�K�-�4�5=���<�i<�5��'�
;��\�\��<8;y�f=��J�-=��3<݌�� *�3)s;TᢼjL�<�=�+�<����]e�6 a�D�+=��L=�ʾ��0=������=<,�"=��u���b��2=�9�<N�l�h�X���l;9M�&V�<�C�<�!�8�μ���i�^|�<�#=��<�I��$�<l�2=HL�<��^�ږ=��=�N��<�x<nQ-���к�\M�3J)�z*~<ެ��m����8v<�
���8���Z��==��D^��۹���H=���;w����+���<�G�
|q=x( ��^V<e��ltƼ:��K�t:�Ļ� ���J<7`;�;��O�?���0=iY��6�_3<
p6;R��aO_=��;�@ļ,�	����<(�*���$=/P&�	K��D�g�A=��I=��>=ǅ���;�s�J=��_��#߼��;*=0�7�ײ =eZf=ge=*�.=���;WS?�p�_=F=���<�yK�$�<:�g<0xx=ۻ��7��9X�_�>���9=� ��-b[=��G=��Լ^��	�n��"��, M=��$=.��P+=�X=���6+�<�=�F~�?=8������<��`������U�"(<9� =���<�,<<�خ:�OS=R�W=�:=�쯼W	5<9����i=o��cB=�?-����<�+w<'�S�u �9=9=�V<�x���<'��:�Y�;�^=��F=U
\��eD�r��:��R=�`���<�'���~�<Ie#�&v�6$�Վ�<���<s���I�<I�[=��S��1l�\=۽R�\E\�ɮ���i���!����9��=��,�__������$�Ѽ�D��I�#*=p�<R�)=@��������G=>�f<oй<�( <��?=�b���2=U�;�
��[3���<�R�;��j=��<��<��H�j��w'u���E="s�:_�!=�cj�[,=�;��N�<$�<���0K�<��PǺ���K]=bԻB�!�,��<�M"=�%9�"4����k�����0�=�6n=v��<�.���ʼ�<f��S��<ttǼ�|\=<�|�҃ �\�x=��F��n=Wy ���=j�1���v<-�1=������üN݈;��<^�<���<rj�<
k5=;�0���:=��=��m��?G����<��"<wqټ�mW��Q=3�޼���	G���Y�P�<'��<�B�<M�L=��=F���z�6�L<�ߤ^=�LO��II�֜=|!�-A=��<����=��]��}�<�*=R �<��<�]��"0һ݈�<�o<�0<R�(=zR�&xH=��<��;�<:=��h<N@@��"+�㛢��!B���*���<�F=r��<�N<i<Ta-=`�������n�=PՇ�̼��.;�Q����<s<��`�<��
����N�B���Q=f�%=e����E�  ��M��;�Bq=r=kK.<G�=��^=>����<ήg=o�J�y�)��b��9�MX���y�<:�%=�d<O���	@̼ �K�W-%���E=��a��[��������aռ.�i��)�<	�<BbN�l�<\�N=|�=��=�t�8ʃ��|q<�=���<G�<T�߼�����2���U=�e�ݭ��p���N���<`��<b�y<YC̼м&6{<u|}9��;76<#e�<��O=O��;9V��G~@=�7J��!��Է�Cɼ|����.<Z�/�|Kn��k%=��8=$���ꌽ�U/��1i�>�<u���<ûf�<��üݛ��"<=(���@�j�z51�g��;߃W�yC=�␻�9％�ʼj�I��j=�)=�H>�ֺ����I;���;�)=�E=�=�y��H��V,=}��/ob�5v=LX={�'���g��<G��<H�<	���6��5�@$�<�G��$Ļ��;4ꭻh}�C�|����<Q�����ü�]�;���ڞ=1�=�r��0M���l���=�"7=����0����K���#�w��<�����X�#=�RT�m���v�= "&�8H�QE==��$�q7v�DI4�E=}L�<{�<H-����<(�-r^=~���_(= ���f�U=y��<�&E���A������P,=*O]�!��<�4G=l�=�"E=�$��t����ԼQ�\��H=����2=�c�=��egJ���<��v<U�[=�H
<E��hj.=�(�ז��F�J=J�㺥;E=�G��ӓ�z�1=	׭<{�;y���Y??<�[<�xk=�?�<`Ch=�tz<�n���O�<��L;8K�<�7}�%;�:a�,�� n�R~A=�z�.�<x��9ք=���'�@��"��Q��=�V���.���Q=0��;L�3=I�<=|�c����<f��8]��GE=����!=�L>=�b�FP0����s�t��:�C���=܂i=�����?���<>g7=U��6����]==� =�<|�T<�Y�<�	b�p�o=A��;v؉�R#^���<ֱr�S�1�$��tB�p>�k�K��U=�����<"Y/<#��=��&=D^?=hؼsE,=0T=$��<��c=����+5<c��k8�<�Ǒ��T<=�Q=��i���_��^�6l�<S�|����;̬�;~��RM=�L�:�%j;�D�V�=\n0��n%���O��O��ކ��Y��TY��D�<e��<|�M=��\V@��`=  =Y�V��qy���*��)Q<��W=iNL�es�=�OO=��]�D�	=ئ:=�����@��S'�d9<!==:�����t%=����P=?���g�j��;�0�<��A=R��<(1+= �ۺ�،�?�I=�+<;�ʻ済�>u��\�
�Rc��C=YU=jKo;���,�<��--=��8c�<û
=c����H:�n��J��8I=$�W��������ͼ}ӎ=,;��vK���5�O����W=j��be=_h���R<�e�n�j�=�(X<r=1���	H=.m<��t<��q�<��<R(�!2�=Z�<�>�A��%�<G=���C��+=g:	�j�8�*xP�� B=����I\=>{&<I����)=�E�<[qG��u{������]��@4�J$�99=�7=��B�*8�;S�P=:�<�|I��06���0�Q�<0kM=�[�<+�~<��=�X�<���<�s*=�Ɔ=�Y�n�dS��:�*�<|��)�5:�v=��<�=1/�<l�1=ʭ=5=���&R<�i%<�`�:/�	��-�<usW�ebX��<=�n�^B=;)�2=�+�׿�<UN�<�xI=F=�;=aL=?�W=�X���<��n<@���q=��=0E=}��<�<=���<�E�=���<6Ӣ��4m=n�)=�>���!=��%=ڦ=��0��l$����<N:=u�Q����B�G;�B
= �#��<�r�^"=�{�<�=�S<l���#f�;�tb�7<����=�,�<s��;�G�9�/=��9����;Y�p<%���!���c<�s+<W�f�:�;�x?�ᳳ<i
��w�;��!�!��;������}=cL*=x\7�� \=��<��*<j��H��1(��-�@;3��z�Z=�[�=xY����W<��=K�[d"=o*-�,_��
:=��8=;�߼W�f8@�����`���=��S=�\Ҽ�2:;y'f��&A<�Q�<B1m<�{3�և<�:�����$�\�����Q7<5'���]=�O�:�I$=G�1=p��<!Q�,,4�����;���F����<�8(���C<�<��)���g����&Nc���F<�\�����:�=X�9��$\��<�<d*<��K<6�S<8y�<x͋;Ǌ;���)=���<�@=����8���4���E=Ϫ�@|\�'�8���=n��;u��<�q=^K��B{=�w�;$�=|�=�'�'��ִ��Q��&������P�3����Sj=�##�����b^<�(��<�a4=/0r<9��<�:=?F%��Fa��
B��f{��=q<D�'K�<K)�i���� R=��<�~�<�[�<�EE�W��=�	�	����3=���;��<�=��+��?V�����+'��0�{y;Ȕ<��D�4��/=�x����<�"7<<υ�\Ҽw!�<�";��%�Fc�<}�o�� �<�}�<������e�x= .=\�Ѽ\�=�[=��C��?�<=��
��"ٺu��f\��Lw˼M&0=���CV_=�<3�^;�wȼ}�A�ֻH=?H����q&=��X���<IǇ<�m�<����L��<18�<�8�=m� <t�W��>߸MP��1�<<�;�_Z��i?���޼�����3�J�Ի�<SAQ��	i=|Ų;��0=����}ؼ#}���V�=h�B;�PG�q�7�]�f;c2L=��8=�.��[<�
��:(��q=L�u�T}�<�䶽�=rV˼��w�Y)q=2["��^_=0���<�E�s/��%��#v���0=��c=�.��Zϼ>H����<B��=��*�<�ə<�$Z���
=�dۼD
򼾷i�Xw��!=�V=��Y���n�\��<�*�Ԭ\=c!��4�H��<Y�=�F���'=9>=Z]�;U>f=߮l<��;���o�y=m����D��j�<��M�mg��u�;p�d<��; y�<�o�<V�8==�'=l�(�;�����y<��:󹺼�U=�b5�eQi���P�!�Ⱥ�!Ǽc�=B�Z����<2:+�bu#�1�1=�e
=�<\=i[˺6�@=7>q�>nF=}�6�Gh<wgڼ�[�<bfM�Ρ��[A��؍��ck=�*������9����ź�+�:�f<	��<�?(������<ųл�ޚ���\=�]
�S���0�kGٸ)���=�b����<��<�O];`S�<�����=��<���X�"���0<� ���˼�,�[�=��C�x:���%8=Z���o} ��K��{�=�D;��:E<�y���=Ab���<��
�<p{
���'=!Q�<!3=队���<����@��Z�B8s*�<oTX�¶8=�_�YA��i=�g��0ԩ<��O�����7Q���<��*;K 	=��Q�)m�O	/�GeK�P�ټ�㛻��*=Ѻ� ]*�-��;k	�<
&=��6<����:�<"_�i�g<	��<�rm<LK�&䝼�+!=J*�<���3���u�tc��r�|<��=��$<j�<}�<��$�@����*]���7���<�|��z�%���xwϼ��+�.�#���=�ݼ��ռ�Z��̘L=� =��g���<�мw�,<������<�Pw:
���<rm�=|~= �_=��6��e=�9)=�>p<(�n<�Wg=4僼�(��S=R�Y��<��B�#;*Ԧ<Y���Q=T=r��d;nJ�<h�<��Қ�<������=�`�<O��<2�J�a�?<�; ��1=_�� ��ܟ<W�w��#=A���r���]H+=<>�<�����|���<�JB=�O����\����K���U���:��<<��
���l����9��:�so<�����A�<�hռ��R�SiQ�D��;߫2�ŏ�N���}1��z�<�?=Т=�$=W��<2q�<{ܹ<Mм޷���c���_<�&ʼbI�<H˻M!F=�"��g�8=g�_�t@V��f��Q��[�|�T=������������P;���9~w޼m�7�^�i��`%=�d`�F�={ק<��=|��4Gb��F�+�<M�<�|߼H+��� =HG�<�/B���t�d=nB���e9=�����Q<7�<��=0�y���n�=-r,�g�4�n��<��<s<�<:��B\=<cM=9���X��9z=I)�<�p�8=Q�;<̀��$
��T��<l�=t�����D����Q�"�����9e�k�GI���1��h�@�չ=S�=�[Y����؛񼝜=�xW��c���qƼVc}:�QX<S� =/(��3=�m�=!��S=��C�]M=�d<O?5=�A�8�\�<�M߼Ik���4=�ü�jż��:;V��<��};D
j���<�&��AQ<��r<��L����#��;(h)=��;��<���<I�<��)=<���e�V�*�=p�=Z�=΀D�Ob�;��Y��;AbT<I�A�E�9�/|<��\��rl�-�����g<x�c��<�*=��`=���9a�&�A=��<�ݜ<�l�;�N�;�=��'~d�C�ۼ�D�:���<ǁ0:7܅�"^<�;<0�*=�y5=#�>�U�$=��`=>�ȗ_���L<�e�@	�\���
N��cg=N�N��V��n���n==+:==�D� Si�6����2L�@=��<+	=�2��g=S�4��<�=�W���4޼�9==�:����<���<�[��z*�%W�:�'2��)�s�<w��s��<C��<#��&b�<uG�!�,=�;�\H�\�,=F���]=�yC�g.�;��9=R8$��'�}&�F�ޥ�<gC���=_�=��ʻ�=CX���Q���V�lF�8~�'˶<�K+�A��vb������J"�Tn��
Z�R��<�㻏@��}�<˚�;�6l���&�8)A=�*R=��%=��ʼk�0�ڦ�:��=�<�̼t�F=Y����E�<�ٳU�?D=x����5B=퇪��	�<�41=l�f�Ґ|=��V<��/��sS��渼����U�<$=��*<��$<��="�)=��n<@�<zy�=�׳<i�w�e+�<�˘<�
ͼs2˼�j|�7���@��k�?=��X�[%=�ھ�����~X=
(I���i=��;[���i��<T><�� <:�r=�9 �,��;GG=�i=�J6�)�&�<�C�HS6�,����:̴��	�_'=�G/<���(I�PL�Ŷs�n<^ʏ<d1*��p^=�� �Y�8�s�!=w�L
j<&2=�t����<9���ͺ�t�<�*=��=q���o�O���c�=�]<�y�<~�+=��$=��=��缘6�rm�� �=}.=R��<�b=��-<��!�g� �;�Z���Q=�n�<iL�%#�<#S=y��<Ԫ�G<C<n�V=3p��TŻx2@=}�
��< K�����<2&ͼ懄;{F��i�V=c�m=oLE=缔۱<�:�Y=��h;���;��=��ϼw17��(�<��j�Zߛ<G4:=��=_�<.�O�5��<}��<.;����<��V�1�p���y��Q��D�"�>�X;܋S�<�<�UN-<�C���N�p�B<7�-�]�;at^��RI��*�^:=�U�Կ�<c;��=�Gf:ة�=:B<$��<�=摻�K��	œ<��_�1Ń=6��<�����~<�Z'=�U��R%�H <�o�<"�9��z+��F=�����0�Z�A���1�ê�\��<<�c�Zf���;�D��+���+��H���༓��<���<�9="`�;�\U����<}&̺��e���<V9=�]��`�<�dҼ!��<Y���8_n��̼�\B�7�3�,T=Q=��1=c�3�k$�<�� ��������9r��{��� ��(��/=7rE;'$7=�I=��	�m�7=�JW�řm==O=��'�ڞ=�P�<�X�<ũ\<�I'�񿄻�SU�p��=�<��M�쌼��;=Q������?�;�ۼǇ=��z�Ķ|��9K��C��S,��%�<��s�ʔ>�� =	�_� ��;����n=kO�=!le=e�&=�-W<��ȼ�}!;u��<�Y�y�ټ���<�ej=���!A8�s��<��
�S��<hz���"��Ӧ<�Mļ��|�7��������/���(	�D�7=��O=��<��^=Q�0=pޡ90�
�R�@<��O��F����<=��	��P��j��E/	=p�$�՟G=�8�<*֫����;>v����R�<�`��e��:	|=֊W�+��<�!�:G���˄<ۓ�;�"=i�=a�l���=yc=��׼7v6��k�:������"o1=~���x�Q�����"�#���<�t�<c7�v{��W�����<�F<%R9;���KFi<���<��\�r�ɻ���<t	/���,=��=��;�	=�/v<嗶�����V�~1$<\�/=���;dT+��T�<��=�+��=�[�&	O�)B��C<w抽/c�����m��<�]<�%<TV�a�<����p�:wB�:�&F�]M�=1F="�C����Q�\�W5��J���r=W�{=E�&=M�#��]���)=���p�� Ҽ�^"��8E�a�<?��<U���@=��ؼ(��<?λ������)�'�;�Q�������v=p�&=�<=�p��#� ��e9�`�*�4�X<8�=e��<��=/�s=���<T7 =&��8<��A=�2��7�L�)����=��S=��	��e�뼘<��޼�� ��0E=�R{���=��4=?֞;��:PGV��<�=g��=51<0�*:Z��<[�8=�oƼ|b=�tH�(�ڼ���so:;�뻦�<rvj��ꐼ��^=kĢ�����5�U����;i��</$�<������|=�ދ<�J�;�I�<�=9=i�<��
=<l�)	A=�<�u����h�>1,�� ⼼w���S�艛<зe�Oŀ<�� ���=���|�i��M�:w���_r��r�U?~<���x����-�<��
���l<n�μ��<̲D�KG7�fR�k�l=�M=Ia���_<��-��� �1�~���ܼ��n�J���o�m��WW=�^���_�<��=5�"=�|�;7"����<=H?=f1=�}V=a�@���������O�!�~<T�z=\5G=�U��z<�25�$�[��b2��^���)4=�ť<��<��<P~R�񗻼�$�<��!�sP�ԩD=k�<�Ύ:���;���<K6e�*�ۧ�<��˼ ��};�77=��=��S���=Wڌ�i�0�|��-i��($=\��������<w�*=�mb<��"�7G���ˋ<J�_=l=^�=S-�<�]]=!�O<��N�����q������=�*:�^#=�H=���<���6S;��J㼷�=�+�<O	���;@� �=ɑ�<^AQ�>�A�=��(���t=��v�2�m�[��<�v-��#D=����*����;:��=�5���ߎ:�+ = ��yȼ\`ü��&�)ڻ,F�<}�T=@�&:{(��j��<x�<����K=<��`=��;�Zc=�m�!�V���d�lx	�����؛=��m�5��;����X�=�>I=�u���"��z�%=w}���&;��=���<�)1=c������<K�.Cl<k�	��.=�r)�0k�<!�a<wl)=�S����V�<�/�=�J�5�����<6�A�7�=��<�S���2]�q<-=16�<��p<Vi��7f-���[=�Nm��t=���<aߐ<G�һ�<м�["=��;����n�9|����7<S��<Gi6=*����]=�����==/�;�Ug�[K���L<��=Ӥ�-�@=[��<Mi��.:���l=�\���|���M=���J%<B��;��ʼ���<?g���/l~��%d��%=�����<�~��]q�<JJ<�J�<[e�<�qW���6��<�2�<�y��Z����<�&H=yo�=���x,'=� m=D��<����b�<��<���9<$\b=IY�������c�v���ż	��м�O �G����<�L�<���� 
�(�;=W�3=�����~1�{2ƺ�v��\�k�>V;<�����<����=�9�1'��%2�<BBW���+=(��;�8(�E�.���0=n��<��Լ.�=��Y=��>���=��	=�p�����<�s����N<u=RK; ��;Ձ��}�<�Zf�k��<�W̺9.W��)8;�4J=�u?����:x�����^� ��O�;\�˼i�0=[�A=出-&��%��;�o6�2RԼm�t���
��I=�m^=`?(=��<8�¼6s3;�`d=ީ��� ��N7�8�D<���:���;4���h[�<���=�H=����e�<Ի'=�l�<*���<�Gp������<�ZH��UN<۞��4=��D�k�W<M�Ӻc�<��\��=XΗ��e��n�<��E=�=��f�[�N9=61�;gs�|��<\Wl;��Q��W]<��<g�N=gc=��r��B��<o�;'�ͼp==[��jb��G�<H^k=��5�T=ςj�qB����<Q��2o�<�]�;� c=��l=�q =M��<�e�ߏ#�ዼ�Ɖ<D�[��`���G;�޶<�9L=R���#=�o�<�j���?���=��)����M�>=�!�<I�h���A�$Ja�$̖�C��B=��'=��\�}]�=QF���7<EF�<c_��=
=�H=�O=�8r=��<�_�O���yE��uo<�{F��E<�~E;��=I�%=hz2<�H+�R�=��ۻ��)���L�c��66I=���=�ؼcW��O�M�Z�M/V����c%!=��<�6�<S	=;�=U�<�9��ͺN�nW!=te����==�C���"��Q=1^�<4`��$�� �R�J�:0��|�g	)�}�"=�.�ι�<�8&<'Z��_�μ5J�=�q;��ϼ��Y���X=���7��<H�1=�����<7 ������A���	8�
t�<><���O�N=�p����<B�=��"<*5<|&-<J�=x'=@�:}O=2�l���y��;l���ޣ<!/=��c^o��=J�	<�=^ �;�T�:MBU�GK��K���E=��;R5?� J=W'n<�q�"�<5ֆ;�L�<��<cq�B�#X�<�z�w+3<��̼��<'��<���r6
��p�<���/
m=��D�k張��;�.�<5�E="���b��і<]�j=K�o=#cG��?�<�G{="E�}g�� v=��\�x��;�w�<?�8=�I;$��sT�<[%�;9W=8�w��m�<�#=Љ��9=v=Y��,==&����3�<�FO����*Uͼ�P��SO=�_���=��=<A���|=>)��3�3:A�Y=u�?=d�<�	����=��<}����<���H�<�F�x=�<��<'��;~�<#�?��~���n��tE�iS�:s�=��e�X�0;���:,��<l�+=l���޻]���>'9= �r���0:�j<��8<jYo�#U��� ��<<�?=�d(�3�j=���º�<�?0=V#=y ��Y^�SS�;��l��ju��=������j�X�{�<�܅=}ռ��8=%i<! �<�;,�b���<%hh��&=a���.���;�}=��>zk<�&=7/$='��x�<�-F�S����;U%�;߮�<�a0=��P��ݸ<�M���L=K/�;5��X�����<.r=�Ǿ<�8M=;u=\��;b��<"x�=eB���H=���E�*= "<E�=���<����mp;ŦT��r=:@=��A=G1���\w�J�<��b=�!�;��g���I��V���P@=��;=߯3��X�/�;���<>W3==�>n��v� �;�=�;�<�Z���q;՛<8\�<S��<�0^��#-�!��;���_q����ܷY=�%�_�;%�G;�y���6�
T�9��i�7r���̻d�!=2�=��z=6�e}=������=�0ӻ�=��W���Z\ =�$<>��v3%�*��;t4����C��<�;@8<+>�F�;.��=��A=ߺ���	�<�ȵ���}�?wO�����|���~�<d"W=� :=���X޼�� =t����B�j����=^'�<ȄK=S�r����<u5�<d�3,K� W����C=B���=���<�\�<��6�leP�M��a�;�~���6�5�[���>=C��_��_�����=<���=ɯ}��I�m�7��V����Feh=C��<A�Y=~��3D�@�9=�ּ�� =�u:��<�eH�:�<,#�<��ɻԍ�<=f3;�<���{�;�����+;>1�<�Xk=���<��;��6z�)!=p���Z=kt�w_=��=V�K<��5<*D#<���<��N�P�M�6�T=�3<�}n�BW<��;��19��g�Y݈<R!-=�J�C ��wܼ���sBW=��<.༛XQ=�)�<dM��H=���9ɼ7Ї<�X3<wXQ<��q�hC�<��F=~P,<��c=� ���܍=�bл o�� �H=�k��B =KV;=�
5��OE=�ۯ��0�#�.;_䍼��<�/����&��P��i+��nU<q;��u�<��A��c�=2�B=���='O�;��V��6=dX$����PM�<J?�<��<����t��A�S<�4�<��Z;��I=n5�(S<��:�<�j6=�X�P/����<k��<��%2g�È;��S6=v�t<�Qf�����i=�NY=���<�5=lȪ<��<&��<0ޱ���=>9
���<��3�|�<=�<�����O=�`<��=Kk,<�G=Fh�<���=�"��L_+=�
4<� !<�)�<,����J����<�dͼ�QC=Yλ�G2�?�<�^j=nc�<�P����%<�2���˩<�/�<�(2<�����r����<.?	=,�<�K9���<��.=��~=E��v`/����<};�*�m��<��<K��u6�<��P��Ur��z��恽������=��<��p=��ؼ��к��<�F�<1�=<�M �S�r=�I�<���<��$��ڮ<Z�ɼ�O����'=yO<�=T�r�:= ���Ã�q	"<E�7�+�;�i!����� ��J�H<�FR����<���<,-D��=�<(;=aF�����4|�;)d:<���w�k��%<X
>=ݼC�6��DR��t;|=�EZ=�<7=k����*;=���0��U��Z'<"�R=�s_���<��x=RY�g�t���"<��f�I�'�u�U<��.<�=��t�WC==�P=F<=ޞX�k*|=�m�W�ż<D�<�=���,�<���;wK=.�[=P�u�=��<�'�<�$/<�]@�����6��<Cv�Q��<��~=�?3;+#����
�!g�;V����{=��<̍9���\=ޫ}<��\���g��Vѯ;��J<�x�}]�<���;]���;='�Z�V��5'=k�D���4='	�188���һ�$3�9j��#�T�q��&�=ɦ���`�C� �y�q<^�����^=���<fB�\5Y���<�����J�
sN�tfC�L�=��.�J���"�#<��<خ,��mƼa:=	G��@!�5n-=~V!=s���`�뼨?=�S|=+.=�g��%�<݀K�Z+9<q�B�����f,8=��� m�M��<L�\�]�}fؼ���<⫃;��/��1�/�I���W=�ļu9'�<��<$,��}�P���<Q2�����<�?=����s&i�Dn=����<��O��e$=�<eӼ+�>���3=pǼ�.�`������*x���#;�,V=�tC�k�b�˦*�X��~�=�5=pyY=�t`=6��:.�����^d=#B���U���)-�<�&�;B��D�.�G6S=Z�A=M�<�	�;���S�����	o���=�_=�w0�h�L=��%�)2=~LC�;	�<�59<�仴�/<S��<�ԓ<%ǲ;�1��׆��L�����I;D�̼\v�Nu���v�z�_=Δ.=���<�x<��O�q�<1���m	=��A	b�j'=�^��L;�q</��<�@W=��;��p����<�%<=F����1=�һ��1���H<�H���pW��i@���$�����o�B��{f������<h�f<�י<1#�;_
=eE�< ��<���;m[�!���&��ۼ#=������︝;S�����`T�;9 �9��Cd�S�I��<6<�8�<HRZ=�`�y1���V�;��<��4��2���"-= �a<�T缁wa=��"�����<~���ڣU�ㇼ��<�Z,=O����;d��}�=�5=UW=`�=�$�<��G���`!<�Y?Ѽ�=>�o=_�=��[	=U���6���<�[�;�3˼h�=]��;G�<��	>&9�ˤ<��\<�c=P=s��<�8��ӷN��=�<m��H����_�z;:ܼ4'S=���k�j=Y�`<�g<��W<1n{=�@a���ּ0���mC!���<�j�W�q�T��;��ӼDc]<xT=��R=[U\=�F���<\�;�]��8.=
���f�;�̡;��<N<�Ag� (�<���<��A�#	����;�U��#�I��駽;�r���b���Q���%@<��4=�k��d\�N�<Ii�;!�c=v��/Uɼ-$�<|R�=�<�}ʼ;v޼��y��󻉴޼7鐼�C����@�^�<��߼�NQ�t��<�:���9����;�1K=�
��{�m��&��Τ����<3�j;%�+�,I�����M�{��<��q=��ۼ�#q<�ͼ�w=d(<˛�<�ȼY�ٻ��J�z��<.����u<ӡ=J��G�O<l�<�Y ����<���<�B=��	�j*S<	�^�I�n�.�u�;=#A�<_�2<��0��<e/��_/=b~�
IԼ �<�E=N8�����
-<� ��I�����;4(�Gt	�U���i=Ј��v�ڼ�/=G�;l�[���/=5�G=h�~���'=�EG�*H�������w-<3m���ZK<�q��풼@K"��zK=�9p;' =(F�;�e=��=ʊ?<�:V<��N=�2�<J�	<�M�ˀ��,Y=��=v�=&j(=ԞB<��߻e��<ă%=/#��$Z��&�O<<;�9��n+� Mݼ�͛��ZQ�i`<�+*��=q=�<õ�<y�$=����
<�**��h	=��:����a=W=�[�Kh�<������;�xZ=Ӓ׼s��MJ$='����[�\��N,��1<�$��A�������*��l�<r�e=.)Y=6"�=�F=N�:�UK<�<a�<%<E�=hqK=�Oֹ��<"&<�q��;Cw<�>�ڜ�<Z���jL�<�좼sȂ��Ӽ��
=ucb=7`=�tѼJ(i��V��)��$��v����C��m=�+o<�L���(c=�n��T�C¼�H<��<»+�G��"�<�|����m`�ܗɻn��9WL!=W�R���*�<�h4���K<�zI��%'� �<��>=����s=R=�gܼ@�>=���e(=m�L�&�K<41�I��:��^=�,���78���7;�E<��=�����û�K�I<b&U;��S���=6�D�c;<D�W�|���=@R~�ׅ=k��a�!�iS=�����<��C<LS+=�f��pT;gn=g�������T~Q<'�#���>���G=(M="=�z/�&g���U���V�8��֚;�TP��B�0�_=RA5�c�<���
� �+�����z��(�+3<#��<rۺ��u���=j���v���=�{�<�)@� 1^=n�==G�=��w=u:,��d=�ؼH*O�"`R�����#�<~��=B�+������V��O��^t=��\<���gbX�*AZ=!�E��|���Lu=�Oۻq��KE��:�<�=�.���=��<>��:�	d�N�7����'��<�E��+��D���m�A�� Ӽ=��<�k-��{�<>"�������V��=����=?3K;D�=fs}<z�<j�;�|���==n.���;=��<�x<=��:=(��;��<²!��<ȼ��ռ�̔��[��RG=-�/��j��G��;n�<�"�Q�g=w>l=�C=˺༉[�����R�<Զ�C�d�aa�<��I=��<}D<;i+�	U���><YA�vZ<�;-=q/,<_<�����ü� �;��P=8�y�����N=���<F��I�ʼ$�O�ׄ���1<���ѫ�<���<U�<t�H�u���������QH2�Şt=��<e.��,;�w=�u=5!"=�Ī;�5�}�ڼpq��fh=���<E�==[r�<8%	<��!�-q���h�ޜZ= ���>=p�@������	=�1D�_c=�c�=ɉ<��^=�==�9��%��Qr=�d��;!=�;�<��M<��A={��d�λ}����4�k'[=X�*�w�$��<�	�h�j�]bP=�*?=
?A=���� �<a�#=�B`<��<1kQ�̼̇���1x<�� =���<ڣ��_��
 =i�4�d�+���W��h���;�.h<���<�Լ�O� ��<�'�<��*;.%\=9�<38=���D<�՘<C[��?��O�<F(<*� �pY�#�0���<;9;5ck=|cܻ�8�;��D���<�P���`=2�t=�ڼ9�<CDD=uY�K��T�,=	4=Éa=k-μ�J"�uz=�
g��&�>�:;�<nZ�<(�n<�*��b==����Ķ�a�<�x����N<�)�cN��mK=��
�??X���ջ�"�<��<�!�<��R=���_<p�E<�=`�=�5=�I ��g=<�t:/��<T=�$�<l�b=�*I�#�T�9���W¼W�<��*���'�ӫ���
uw<Mɩ��a~��>�<���=��;:�Ĩ��!+=��N=ሼr��9�Y���z�|2#=�+��j�=c�1��4=qc��`X=����/�:��<ͩ=��(=��-<�HW=b���F��;L��=�� =�<�9��O%=M���!2�<Hڼ�H =�hż�T��BJ��n:�=��;�G����e2��<�;�c =��<�&�7�=�&4l<W	�|eC�	 )=��l=����?&�S9�<^���g<z'� kn<�e^���3=w`�<\�a=���.�8=�6���2��1+=��U<�u�׀=��c����;�_���SX�aY����\8��m�;�nU=�=q�Q=S��'y<%w��+]=C��<��;{[5�)�E=�ۼ�4�����_�=~eT���ż�d0=L�#=F^／v=U<�{!� $�h�;���<)���&=��=q�߻��<��l��M=&Z�`H��y�4r=�Xȼ1:8<���b�̗1��o���꼢��<�0��`=�s<
� ���R=�U�z-=֌H�s����QW<�a=��=am�<��F=%��!�d���B<��q<��=��BQ=�Oj=�5�"_Z���H����<�3���
�lF=�<��̕<�i�;Yqn=�0s=�3�Q5��q��~�<Aw*=
�W:(�R;�38=�#μ�������<S�[����<����=�F5�e��<��<��J=���;��޼q�N='�i�w0L=<f�$�;��Z=Z�C����<>�<C�$�a~!=�����:jJ<6ׯ<c���#�������|=�B�Qm�X4����'�׌�<u =��� =��;����=F�<\V��'A=k�U�3�d��=^�i="���3�swH=�m<ƅ;���;A�H=�O�<`�t�v�<=�:�JV��ݼ}�d<�`�*�\��ET�����H~��LT��p=��Ż��Լc�#=X�<��Z�LO���ͻ�^μ�W�<`�<l�Q<pk'�ki�<�>�<
q(�>b!���-�}��<G��<Ǩ<���Rd�<��%=�b�d$�;��>�8�֑x<T�1=�b��>�<��f��?/� *c;�S�4bq��6c��Q=O�s=-�/�-�=�`,=7�:�%��8*�:=���~f��0�;D' ���<��ּ�f�n,A<�s=.|/<"D=(f���$<��Y���<��1L��^�8?|=ٴD��pO��B=8�=�A<���Ǽvٿ�lk�<i�~=C���M=�M=�̼�2I���l���Q�Q�<�r(����A����:����mʻS�;�|�qb����ȼ��.�������7Ƽ�f[=�n�#���w��<�f@<D�I���= 6;$�<m�
�	�\=յ<�?<���<��$�&=:l�;j@z��6{=#�p����<��C��m�</m�;4=��滣�o��zV=�V�R�S�S�<=�����!�����O&=AfӼ���;K� �H*<H�=�Sؼ��/�Y߿��A���7��\����=��<���<Q�P=x�W=�%�=Vt��1=�c=tiX�,f<L�C��o=�j=��$�2<��I��N<��Ҽ��F<?0v<K�w�R�g�CyC=1s]=s����#f�R��e�m�	�>=�9<�\�;!�JB=sZ�<n�C��D=Q�����Ќ޼�%=1f��7��#=��:��n=��.=���96�<}I�<El�����QI_��)zG��r�<`g��1���ƻ�)��"�;zE����;	�%�_�RV)=<\�����n�9 �<t���h���L��<'��<��bk���i=���<ڶ=�"�<w=/
&��R>� ���ۆ=��R��ռ�k���V�"��j<��м���<�2��7t
=��=uQ��,*�w���<M�B��6A��3`����#-<َQ���ʼ��T��i=�����wμA,�z��<=�L�&�F��<tK=�=�z;�R*�cNw=�=�o=��<�%=�*&��+�<T=�2A���W=�t�%aӼ�S<0f6��&�<+&�k@=4�<u�<���q�ҼB�A<��<�����J���c<��ۼ�U�<0<O<�'�<xST�}寮.:���;��7x=0 h���>=��=��k��=<�D<�겼f�A�4`�c��;Eǧ� 6�PU��4����<��#�.k[=j��=Λ�<�_��������1(�b`=J]�<p6y<�n�e�j�h��A�Z��j
=�`<��8�R.,=�J���m=�R=)�=���3�p}<!��<�~� ��:?%�:���<�4�<�|��^3A=Y�g=�1z�Y��<�0�9�=ޥt=���~�=�q�;�v�:��;7qH��1Z=ޥ����<x�X�+���������%k/=�>��;g���Ӽ��P���4�/�v;ʛ�<���<Z�:3yI=+����_ٺp:�Yz<P�>��=_�+���ڼ{���d|=�=z�<Pї��c=-���;#=�)G<�U<W�<�y$���C�CN.�	�YP�<v��T�	�}�R��@E=g�<CQ<=f?<�Ģ:�M�Y��ءo=�ļ����p3�<5���%�lQ�=��p=�(</��<�t���%�ă�=Y�9;^+=�<^Hm=
&���>=���;-m�<������Q�5�2�!�<��=|}���V�M��<�z�Y+='�8=YE	�O&j=��L�?���l(���:���<=v�:�6��ʽx�3�'����[�;Ź<�Ļ�v���*=�/��,��;�$���u���G;��=dN�k�<x�k<��3�p0]�c�/��&9��y���!!<|\��F��Z�(<WF�D_@���<zʄ<��9=3�;���/@:T]l���պ�>=�y]=l���`IO;{��4R[<�յ�$ݒ:��C=IW=�H=&@q�ӄ���z�Qj�<�Q<s�o��yN���=�,�<i
���%�̲<��6=��<��#�3�~;���{�<�7�;k�^<�%�`�h<�h��F�=���SE<�.	�/ҏ;��ּ	��<E�J=��)=�a������7L�=�H�%^<�|�;�g=�r����y�DR�<;=�j����<X�=��&���K=�w<��+=�C�<8�ݼ�z=��
=a�8�$=�9=$�ۼG�F�!�8Z=�?��<�����|=��3�z=|��f8=�����f�6�;=��<B�=�a�ce=($���
��Mm=u9<IWb<�|Ҽܼ鼏,]=j���J�;oQ��λ�B=\`ݼ�����U=�P:FI"=�� =�|=%Eh=�=Q��ˣ��&�<�S=��<�<�n=���;0�_�O
R=�衼#�)�Ӳ�N��j/��x��#�c=)�Ǽ/>�<]j���[=)��_�����1���!�!%=魾;c��:��<c�=8���6����j�G���2�F�\� =M�<Qo<�4M<��Լi��0�<�AYE= ����g>=DμڤG�I�5=e�E=�+»v$��I��O�u>R�]	Լ��Ѽ�q���
M����+�s�֟�<,G=�X5��A�����/=���'�[=�rA=��V��=�Y�<N<u��������[�<�,3��W�5ם=/:$=B�ǻRf����� �:�<Y�1���=%�<�(9�K&A;
Xw��F=<n=��W��<�<=N#����k�u;l��Y��<���:8�Ǽ��_�4=�E�Q�c����/=��A=i��m���� �s&=�3��b!��ϼ�zC=��r�������G=��M=y�s<���;�O=I��;��g��Ֆ<�s!=�y�;�ͩ�!����<� �=Ȱg�n�D��[�=w�་��<��^<z�H�n.D��zh=_Q�Ef�<�	����[�(;$���S�0=�,=g�E=���<Ax=� ]�h�<8$��+'�P����/�Y�	�9=jȘ� =N��D�6�K�^=l��
J��k��FY�x^�<�v񻴮�� ñ��=1tN= J=��t��N�H©<3�=N��!I��꼝��:��<�=K�5=Sx=����0(=x�<�k���d=8u=R�����O=��,���g:Ԃ7�l�i=��H=P�:�{+���ɻ�R<�P�<֕�<W<�\-+��ђ��\뼞��6�<���a2-�x|�;��i=j.�[�;6[=
!��ȯ�B<_����P/��&�E� ��W��s�=	64<�&!=G���E><v<���;�pZ=�s==<ϊ<��I=�s����=l3��_t�3q�l��=��f��`Ѽ��K���=Cg��\��D����<�G������h���)6+��fU�z�ae`��J�_lB;�7=����$\�=�<;�����Y���<?=H�-��/��}��a�w=����������;T`,=@�K��h=�F�����k���L؄��'�Z��90A0�kr=��4=ơ����<P�;K����:u��;B����$=�����A�����K=6eO=a�3�J��Lؼ#��<.W�R��=�z;��(=��V=b��;��<N�<��==:�OH���=��=�g��c�<0bK=��1�{�<P�=#I����;�q��	��)�+=�`o<��\���r<�j1=�h�A=\f�<L=��}<�vn�$�<���;l�]=�R#=�C�<�H;fϿ:~�#=%�w��=|H�;�"i='�W?=�s�<Z�8=�N�<�)��I==�eN=�q{����0˥<�.���#���<�A��@_=�La��/���2��+2���.�Vd�<���<M4��v@P=�&2�`S�;	�=�|wE=%���y=n���x=I	�)P=��$<S�F���<���<�p,��X�e)V���<l~�;
�m�*�=���]=���<+����vɶ�z�<�'�.p �;^D5��:="i�<���<+�����n����	�I��6[<�><�{0��a���;=C>���l��;T�<1v�[�<��*�@��=�m6=��f<��ټ�f���Y<r̼�z=��<�#�<���F; �V���;sw.��X=�+�<�J�݀8;��6��"�;�)n�ݬ�<�Uf<�Ӽ���������=���<q屼��<Br1�*�r�f��?ؼ�.=T�1���U�=�*=^7�t�h���<[�
=hM���Zۻ�;X�J=�<���/~=�)J���=�RF��i�<�c=¾B��#I�>=�n5��uT����<��2��H�8�X�/=J/#�簜��L}�uo»,��<�A�3����=9j��w���G<^�����tZ��;�:+��;= ��Q�a=ȡ�`FH��,��P�;�2={�9<�$3=���K��L��<Tu=����Ց����ֻ͙<�9�<c���=�t�3u�<;`?<b}\=r7`���������:PXۼ��<d�f�k<켼w�<HJ���	=���Nd�6��d'�;,r��0�;n��&�<�����]�| E���=�9  ǼN�<��;�����<�V��*�w��G\<N���� �;)=�P;�b=���;�"�;Nك=k���81�Z��;܆��}�;'%���Ȼ��=��<p]�<k=j(���a<гǼ+�=����d]=a^N=|�0=�M<X;%������ۻ6+Q��aC=�F�D�==zb@=a�i<j�����:�$��`X=b�U�z�=rt=0H˼�ߥ<��h=�ż3I=D
�;��#��L�:Nm���3��K���<R�Y�y<�,=��;��H���ndǼ5:�<`D=c�h�ssF=���;̄=�R�<[g�<��7=�=q��<7�<:$;=�E	=�P��ϼ���;u���iy:�����H�^�_=<~)�e��<���;�؇<�!�x�	=я���n��K������u��0�aZ�<^n��|м:#=��"=
E
��=<gAf<��Z�~]x;c���b���z�<�/=�=����S=��A�>�<k`v=ː�����"|L��a<[W=��{�3�JZ=R�ʻ}ĺ�����%=V� i\��>�<֩*=[�<o�_��`���j�7����;�<�9X=��~<���W�<q~�����M����=�9&����<��Kb����LƋ<��/���$�G��<���<Uv=O=x�;=Cy��+��<.�������a&�W	 �f�A=Du��L�w<�8<��=#�L���^�T5=?=���<����
�&�<Ǩ�~�\�gw|�H��<�9�<����<�
=K�<��{^����I=�M=們<�F�;�M����TQ<=��<�����J=>{��vD ��R=Ɯ�;�#�O��>:=��I���<t�;.l5=%.\=:{�誻`$4=ػ!=�,=�a%�;K��X�ĻTƝ<�B�r�3��-b<#k�;�0i�mW�<��;�&=�銺Ë=U��<�0'��4�#�:4,H=���:-�M��/⼦n�<-���Hzp<�לּݜ#<�Nt���E;m%�#w?��]0���P;ZkA���<�%<�3.=�W����*��B==�ؗ</ú�껈�;���٧����!=f^X=cA���;����<��c=7c�<�TL��o�o�A�V8p=\�E�ͤV=�/�<�ns�U=�k�o��;�L�<�<��o�4�(<I�F�Y�G=��i��d\<�?H<ʏ�<����bog�%Q=������;t�=o&D�U]=jl�q��:�>缕Y$�0Q[�8c+�B��;�t<���>�K�ף���#�<Y���}�'= @=����.=YP����:|='o;=L܋<����Q�<e�G/=��4=@�Ҽ9�Y;��@�i]g����<ȶI��k=5��<��:�36\�	�ļz�=r+�T=�~s =*�v��fY���%=Q��"M<\�$���_��`��D�=�:��F�<�.2=\��<�����f��}��t�$<�xS��Z���<jb���\����:,�<43+=ּ;8q���I=���;%"�;w�c�1��eI=���:��f���{=v���ͬ��Q!����<��Y=.)�<���<�$v�t@���ܼ����t�a�Q��=�$���N����ә�<���<_�����;K��;��.�����=�=��x�p��<�q1������ ?=oj�y�k�4�=hR�<1�G<Ӳ��G�<�
;d�1�%�Z<>�<�=d��;�<:=��:�3D=e����A��	�<��<Iͤ<�lR=��.=���c�H<E�=<Z�Y=ב�<U$����R*=�].=��*�L�; �+=Ԃ
��-:<l�;Ch�������̼�[=]D<�3��������+h�u��PCҹO��5	=B{�<�)=}G<�rC�E0p�+�O��i��n�
/-�dX���>!�k����;���ͼ�) <�ꈼ?1�;t2�gD=�v�i;IBD��kѼ��v��C}��u�<�)�9g\<j8:<�/�O{�t�/��=�A=�>=��[<�??�@�={���He=R"=�EP=�t2��h���/=ZM=�(v<�b�<�D=�X���{AA=n�ռ0`���D���R<PC$<�����s9�;?�����=8=�<go�E��q�j�B:�}s=SY-��+A=�>�|v�<�$�<�y��"��(��b-8=i�*=!����e4+�ɗ&���y��a�[���1�;q �?Tq=/'�=$����=�4I��0=���<�K޼5�;�>(�q�>��l\=�YJ=�W+=��/=1-.�0r0=Y�=��-�h��:[�ػ�(�{`<|�����+=4f?��<�<�%��)���@�<���<E/��)�c�t�U���}��T8<iG���W=n�j���$�r���X�D�����D��<+�s=���ڈ�Kq_=�C��{/�:�r��G��p;���:��=�Ǥ<;������V�=�#�חQ=�d���H�]"�;��l=ǂ
=�;�s<P$��.Ud=곽;�3=b*��
�:_�1��h_=b==���W-�MѼ�/F=M��F%=8H,���<��9=�����;���;�=��<=�����<��B<�H�^	�;wc\=�ܒ<�PD���'=ϊa<:ͼ�q���=c+��dU�*�;�N�R��1�:�I�ϯ7�/�ܼ��#=G��<�d�<ê`�	�=�Q;�gW��P�<C�C�Kb<��09�.e�9W�0)!���<��R�=��<���.�t[�i3��*G���=�0F�e��<�;<U�A�r=��8�g3=�����;�x�:�� =T]J=��s=�Y*�H�K=%�Ӽ�\<��<�?��g�q߫<i�<Qfλ
�k<�?�� �M���/��U�;�(�ފ���ѭ��
d�w<�sN=�d���"=��*�脼@��<�ߠ;�&���v�l�T��Q=[=�`=-};-�r=2؎=ԥ��N�^�hK��[������Y,=ب�<�lR��@�<澲�0�3�x�����x��<�ٺ(�p<L�<=Fmȹ�.�<e[T��T�<�D��پ��==�O��I��Ս&=�.�<�R<�V=�찻��_�X�<�Y�<�%�2$=U�T=X�
T=��*=�^1�rS>��ZT�xr�;`�<��
=9X�<�%U�p2�����<��#��R=��m;6=��a���=;W����3�8,�:t�&���|�Ϫ�@<I1�Y�%�or��| ��8j��(T�█;9��<��a@��Ɓ1=�� =m���p0=�3U=mK��4�<=0�=�ѐ���<�1<D�M��fJ%=��@����'��]�
�e�E=�Q`��<�o9�������<OyF=V�WS`=QG�u�*��ᙼ��J�+�"=��:�2��!)�ȿ>=W��<z�=�h	=C�\��=�߉��J��=��<�[��J='˼�����nM�={�;�qM<�
��`?��#=Fi=T�Z�� K��<�se��.���[���=h����ŁO��==ӎ<��[<�Io����7=���Ɣ���W2���:���������U=�]����H�;"�	����<@<����;�b:�����.�"=�<��Iμ9��;�����2=T�<b7�٠�<��<��H��L������'=9�$�{z��/Z��+�T������j��9�I���g;��<k����2���<;�M�<��=Jca<P0=�U=��=R+�<�(<�һ�s�S<��׼"�N<��O��J�;���qC9�m1�V\=�%=|;׼dK�<��<\D��Y�@�1�@�Y�{�؊�����*��6=�g�<�� =�]�;ג��B%���:T"�<�y����	����<�c=�\=R(`�q6V��i�<��d=L�
=C�/�ļO�I�`r=�^5=��<�dܻ�d�;A2C9���'�|���E��c=l�!<���<�в�&�>�ר���ۼ��l�dTe=1�ռ^|)=�q+<8F=7���pf;��n�3�@���߼��=��~����:~�=��Ȼ/�Ҽ��<Å>��++<ϟ޼��m���̻�[);�i=HI=�P=��ڼ��4=:I����&<���<�G(�ij=E$<��U�<�ۼ����Zx��rn�Kݍ�����G<~]�<��@=���<���$�<C�F�"1��(���>��><��F=����8���<��I�ൻy2��^=�	N��ɯ<���7*��]_�5�<L�<,���gYL=�uZ�L7 �!�<w.=���Wn��X�=��/=g�<��<-��d��;�W<;`j=Ɗ�<X �=DM<�=�U4=M17��<�^�<��W=�>=_˻�I�;�n=��O= :�������	��u���W<�W�?�<�K<�ݾ<I8#�P�y;$�R���<x�J�3c>��V�<�e�<q���#�a<͞<=B�<�ؼ}{l==3e=�������JZ9=�[ܼ�6,<�q=Ȋ����<;�=U�޼�(5����<A�T�&��vl
�n�R�*�/��g�<rC+��j�<�<<*��U5=��b<��p=��<={]�=�n������f�;���ǧ�<#���9,��'��������N������=�޼1i�<G��;hÄ;����!꼜OC���O=�'�+�<�Ɛ��.=�:g=��=���;�nt�6�;=&를9]�<��_�<1��<�9�n�=�=%󰻑ס�d}��������^R�=�g�:���<� Y���<ɻ-��C����t=��D='�8=#ZA=�B <��V��G1=���<��B��uV=�5���b=�|U=cđ���/=�h=ӓ�<"��<��ļ1~=��=�<�����<O:=!�P��ڋ<Yzb�dTG�c��oY�<)Y�;kb�;��@���5=�aF��mJ���/����3B��D_<���<CVY�$Ѽ�.\�ɹ��F�?=�+^<zn�<d�=������u=[.�O�;Aݼ8�����&<��;��3���#�<��=� =#�H=y=�Zü�����y=�r��ۇ��|Ѽ�f=5 =SJ��!���= ���ǒ���<=���<Fw�����s�L�����l�9�(ɺ/{��6>��I�<�4D=W= �^=�t<a��<��2=��=VCh=��˻�-�<�<1�#�;&Լ)�2=qw��F��;d�f�L��?�5���b=V$�</Υ<�V:=�v!��t=��:M�-=f=A=*���g+=M��D�+��*G��Z=5�<@�A����<��*=JlL=,Ө<�:b<�cj=��:�'�K=��B��6<��H<G�="=d�<L =�5�=9�)�x�+<�Rb=h&=c2
<�{ɼ;�H��0���G<�*���^g�<{�#��&=�ͼc&��"!�֬��F=����е<΢<�0�ayʻp-�`D,��d�:���z�'<���;�'�:rZ�㸟��ϼ�"=G�=���<PZ=v�$=N�q=-�:���C��<�'7���j���;q =S+2<��;/�D� �A=��J<OA�; dD��<vp���C;z[j=S=F=��<��7=�Y���.�Uql=�@ؼ�
��?L��~-�k�c����<�G4=�?�9��=`�z�(/�<���;�iY<J��<m���n�<=U��ux=O =�0=���;����ħ��:Y�#��oa=�+B=�wt;�H<��X<�O��;�@�8�W�o<7}<��<�w�;V=Óu;��޼Q#=�Fr=o��h��=�A����<���<|�X=�Y=���_�i�sR��rh^�3�=��$=�68���<Su=3��<��9=�K�<�礼�e=]�<��C=cM��guH=�y=<�K���F��{7���X�DQ=�!\=K��z�@<�І�n��<�� �xw�<3��<h�%�3=�%�g��<�*�<�r��j�;�=����r��t<CoN=L�T���Q�_8#=���<'$w��ߤ<���6��<dP!=n�V�R�	�.7N=���<1
=�Q���?�~+�<�3=_X�jM�<���>���T�<X�	�����H޵<Ɲ��� �X�<&C�;��f�uB��9;�e�<b�-=�%=H;�<T�@�1qg<�,=<�&���FF�e����T�^f꼑�= �A=ş==)Gz=4L=8�����`�}�:=��L==�'e���1<�<=�,��h麧A=�Ж�po�<�YR<�QZ��Z��M�㚏�B��<_�r:�7�<48=�H=$e�<U.����wټ��<�����X�;� �<@�<Ea�;/
�<5��<�Hw<��h=��N��~�<�c;����R�<!�˻G��L�-SO=d��<yhK��j�<-@Ǽ���<�y�=��=�d���[!�O����U=>�y<�y@�*$D���O��1<R�G=^�;��˺hmº����Դ�:D$a<�;=��(�_z<���;��;/��;��[�u����>����:��
�m�=���<�����<��&��ݽ��ݟ<��R�@�><ᆳ<���5�~��R�c_S�3-���X�ЂU�a���ӕ�<����P^�Y=N�;1_�;K�0��/=ɩ � o|��2�4��ų�:�H=�l=%��;!E��?_��Ko�E�E�ּ���WѺ��<�叼��et���U=�e �lRL=N�e=7�+�������9�G8�Ṇ=`�j=�C<)�<�U$��r�^g��/n�W�O<�v�C0!=e�==�B�b=�JEM=9S�߈� ��|N|�l����A��l�`hi���#��~=���3�Ʀd�-y#������=Qt���%�d�;�5=xd��)�<���?Em=���5w4=�K�;Ib��������<E��<$��<0��<�]"��T]��k<Q=���G�=�=�=����n�mli�?�;^�;cB]�է-��P=�Z+�ɗ��*�Y<��缤 >=^��X��<��o��^o<�¼�K;)M�<�`<gs�<��~=o����� ?W����<	��+Z����<O�<b�=9�������V�)�<|O�:�]��<��Xv���;����}b=>��j뱼���δ7�ɱ���u�;U��<�=��^�kW��qȻ<c�<v��=��*�MG_=�3"=h��<���<ɆѼ	\;.������o�3�B��G��QL�����tG����<;������}HH�7mt=�.=_'��%+ټ�L�<7x�<{�;��B�<�6�<T��쯼��g<��:=�.��:Qk<�mt�q迼=�='Q����<=m�j@��I��?�=(�v�ؠE�M�u�=V�<
�=�
I<�~���~��6e=��'���o=X���� ��)�=�yK;�4=x����fs=l���Ñ�2���������Ӽ6=SЀ��oO=O��;��=��j�+�<0��xW=��D���\=T�<O=��?{�PE�<W9���p���꼎o=�U�<M*��vK�����K��=�<�������<�I�	���f%=�:�͛�P{=��z=�%=z}0�-`(<0d+= �;�sм-�;h�;�W�� U��h�<��r�ᤐ<��W=5'Y��
���<�	,={�=<5�f���=����c=�<�7Y��%��|<k��m�<:��<�*:=����ʸ<���<��x��ֲ��Ի��<���<�<��)���<�ɚ��*1�jta���)=҅�<Q9=\��=$�|=ΐV<6�1= ��V\q����������m<یȻ�<�eP=gp����ͼUa��P�E=U���~ =,4�<r~l=@õ;BL=V!0=ʢ���;h�F�<=*Y��g4����9�Ӡ=ā<?��S�k���?; �A=�#���=����? <���=�i|;�A;䞻�I�D�JJżyr��|��;9�$�@呼ב���<I��w�9��E���4�=��4���:�jܺ ��;�D]=&�;�Ǆ/<���<�n�<>�3=-�d<-u<%1=Ot�<�}����o��=�
V����<<����N����<k����8��s�<�P<B�C��i=>ۄ��#̼��r=�r��`��Լ�V =R�<[*��;<+n�<sPE��p���&=��=��t�ร<h;м|< �u��z=���+��<�Y������c`��<�4���Ɔ���<=]��qB߻�=��ǯ<r*�;e5�$<޶<�h5�
=j	�<N9�X��=��(�=�:<�V����ƀL=Ή>=�)� �=>r3�sf=���<��c=ǈ�=�g�<�4�����<u�_<J^<:�B=�A=b��5�;ޞ���'w=v�<��<��^=¯��5�c<���<5���ǟ<�l=�ap�o�1<O0+����<�_ܼ��<�`*�e�� i���U�Y.Y=���<�lƼ��~���a��9n��;DF���aX_��`��Wxe�%�"=%�X=m8?�q�;�=�=�T����<�	=���H�`��[��Gv����~�w���Ļ���<� s��]"��λ<0�%�b[@�3L�<c�����@uؼB|ռb*�=�ڇ�xW!�s7:�)}=�7O=�V<��<����K(<J7=,[<��B=�Vz=�1`<<.P=/�2���;bAK=��h<�OA�H�Ζu=� ����p��#�*<��;/�X�^����ސ=ꇛ�E+����=�$�<K�/=�tһ��K<j�<�=�j]=<D�6�(�ׇn=h�a���	�9I
���D�k��ѷ��\���!</짻½2<#�I<R0����;}�����v��;&�=�t~�<�s@�ؓ�<xJ=�J	=�=��V�%</v���k:�� <��;�<"�L<��T�(=	�>=���<�����a}�����?�<>�="''���X=��ɼVD�<��.��!��+��#D=wgv�U�J���>=�C�;hn=�=�t=���X�*�k�N��o3<{b<�9M=�E�����:�s�<��lW�;�3�el,��]9�_� =h�<���<�R=���P<�K�5�=�PF��<���;U�a�=�*=�$���T���D=c�_<o~=͓ۼ��Լh��<!���杼���<a�I=y��<	{�=ʂ=��a3>�6s���.,=��1=#?+=C��)޼�E<�{5;f��<�t�x=���>��<���;؄=��Y;�Q��[+�5�L��<
=��.����;�kn�]b����ѭ=��b<�k��o��M^�իN��=��K=T:</�&��tѼL�V����<�)O=V=w<�i ���=� ҷ</�;p�=�߲<��<"�	��)��lOL=�Pﺚ%�����=�bF��T9=�8�<��%������-Ҽ��=�����;�U�εH�?�ܼ��<4xZ���=|7���;5gj= 1ҹ���j�g<[��<���=#����4<��� �M= L��#��^��<��9=I�o=���(�[��y ��/z�@d��h�<�� Z/��;���:��.�<���)N=��F:��=�O��}�<�=��_�yQ�<�lj�3�_�<�<���;���,��:]5�;� �B��;�N=����
-5��P��V���L�b�=��<ıۼң�<�i�`:�uh~��k�m�7=�;Sxn=��z��r�<��o�;�A�rn<��K����<"=��'=���>��<�5t�F)�<��:<H =��<��1���<É�����!�+�pE@<ו�F�ż6h�<�<�<:�%���"=f�=,d��q��T�i2!;Z����!=�H��jG&<Ro2���ݼO�k�1j<q��=�_<�o�<�E�<��=���<5iD=�̼]�C��;6Z�<��)��]@�1kk��sM=:0>������9�K���0r�:���=+�<]��~;�Ѕ�!�7=�@= �<�u=+�O=����7=Z���)N0��m��3�Ҽ�i\�2�B<wY=he��xy<ϳ8�(�6�.Cf<���x� ;Ŝ��!:��չ#����^(�<����[=h�y<�%�<�e�<�2��d鼽e�<��R=5AƼ�*��{�;��=�b�<T"�
CY�m漠w���|A=��0=+Q��69��7߼{5=/pS�����<��<r=\;+�y�7-��ԎO="ױ;0����r<�X� ���I��5�a^=�aɺ�	�����<*&̻����M�	Z�N�e=VӉ<�c
��<�� ��<���<�8 =�ґ�,�c�qY� O=�7�<Yc�=W���~7�@� =�� =G�伛H���G�w���u��<�QK��Y�<�m0=nj0=���o�<3l�����='\Q=�)@=W	y�<��<�X��K����ý�=)տ<�CC<D��@�F=x!�=&� �P��; P���$=|��<n2���2�^W��϶�<���<j�c<�+��(1=���<v���_�	�l�R=�~R�<r|�=w���'H��y�;k�w=HƼ�C0����3�9����(���^�;�pd=ó=���x��<}?�<-�=����Y)�n�,=c��<<��<�t=T�'=аi<��9�[��<p�
�Fo?�A�ٰ\<����EF!�#~������<ެ2��ű�Z�
=�� ��ʻR<�<;pٻ�\<�sy�΂�<�&�<h+� �t�&�0�on�Ċ��1=k��bv���"=���;���<��Լ$�\�g�#=�v#=��,��K���V���!=J�I���h;Y�U��{�<;c=D��<��=������o���/�Tn�p>���<D00=��*�P�<-r�����<m�<=��=��(�1(J�v��<z9���f��-�&�#���W��=����B�Z=tG%<�q_�Kj����B�:.-;I5�<���<�f���q=q1*=�w
��rm� P�m��Q���	�;t�D=�of��}�<G��<啮��PF=]�\�0��<˿=��Y�����n|�<����ҿ)�	L<�^v;d��<���<s&/���<T�q<�!I�� Ӽ���9!s�=c��<+E&��k=�mW<�g<����7<K=����=0�;��T!���}�\�N=��Z�l<�G��.2ּ�S�ھA�-<��=��<� 1=�b�m�n�y�ƻ_��;ɇּ��C=r�<yka�'� �9_'�ߨ�<��e:�x
<jۃ=
�!=��<i�Ӽ
�N:濣<��p<�̼$�2=gd��vb�F^�;�(<�k<5{&<Y]	=N�W<�y];�,=#~���<{ݤ<w��;�C�<3X<�'�'�j͚;���<�_���[o�x/�<�dz���<� ���N<[��<��3�L�q�!��"=�H�������q��A=�=�j�<ߚ(�W]=D=���R�,�=�=KƄ���;�27�P�^����S�;ʫ=�9���y��*=��k��Y�;ww��7� =[��<�r�<��;��K"���X9n[Z��}�=X�-��< �=�6��B�M=���<���8��2�ͼ�G�;B�=�B=�B�<0�I=�=��[��5�<�M�<1�μ����n�W@��3Y��W�%<>ټ�;�<0*Q={9�:9B3���ļ��/�1pH�)��-��<H�O=N�s<<#�<�{�>����E^�c�==;w��ؠ�<�S�M�&���u=2V={���%펼�Ez�>�g��#�<v�;�KY���}�E�"ߕ�ޞ�1h3��#=�a�<���Z.T<��U=����h���<��<=H�<"Ϭ��`=�t=�t�<��1<$-�3�}l�<:'Ƽ�L��f���""���<�-����� Qx��~�ǯ�=3-T<��ӝy���=[G.�}���2"�8v��m!���Ҽ��<PO���=����T�<т�ĝB=�s��_��c��_~	��b={"�j�+�%{�z��|y=Y)��WM=�<����E�<j����;��U���.<;�k=�<f+-��H��6;=�d��O<a�k�H=�u���"=�g���+�0	l=�f�<;��<�Z|<K+"=;�=�����>=�A���=H<]w=��<o��ŧ���~#�T�&�����e��i`=�i=kw���Ƽ��<����zW�:��;�q(<͖)�Ȫ9<\�=�;>=.d1<>�»1I<I�Q��:�I$�c�6�� ���=�W̺	yD��:C<§E���ݼH~/����S�<��[=LE<<��<P�ٻL<A�)=4v����=# `�5Ԩ�?{X���;�N><Z�G���=2)��4�1=qq���=BG=��l=����nֻ)��q[����:=u59��Ҳ��w1�	+=�L��d���B�<!:%</�C=��4<�4����<	��:j�_<�@�<�+�<��<]A��Q>��.S�?BԻ����md=��u;(���e*�<|UJ�(%�< �ȼ��*;�V�<��#=#0Y<��k�P�=��x<�z�?Y����=���kw���D�=ʙ	=�Y�<�}w;Ga���LT<�Bw=�/=�?κw�P=D�P�W�S<��<H.X�N8�= \༜C<:�������%�<������8=�с�.G�<��=��*��	^�K+<��h���_Ph<c);;��;az���]<��<�|P�f���QOD<��$�m�}���7���\=�t��Q�C��h=>�=D$=r<
 ^�
�2=cz<�j=�D!=��|���1= y�<�W�=(�4< �񭔼mZ�=�;�; ޻1�ܼF���W��0U<E�b��=f�5���<�=D��<k�E=:�/���=�d�;�/x;��<B�l�������<�B[<zg!=Ȟ=8�A��=�O���ዑ:��^��.�<�;=�Y�� $��]i���ܼE>:���Y=�Sf�H8���~�<��D<o�p=��=�g�[�[u=&K�3����7����<�^<�2�� �< [=��M�C�<�yN�rx-�}�6���W=F�d=��;z^`=�s�=�;Z =>�0=+�q������%i<P�=;�`=QQ<r�=O_�<H�L<�ɼ�R�������4	�+t��H>� ��<G�<�Q�x���jT�r�};0Q�<V@/=�"����;34�<�<�<+}�<��l<��[�]����<` 1=�,��/��F<��޼|wĻ�ᅽ1�)�q-�ɚ =�:��X=y,:_�B;�W�<A`���Ӽ=��=U=�9B��8�<�n�<+�</�B�d<h��+m��FT�%=ׯ�<�vn��V���N�����T9<�$�<Ņ�<�L =�6=��h=P�=�%p��%��^�9��=�Q0=:<=ഈ<�g�Q#���]=k�X=�[9=�u<R�<-�=�fV����<b6=��L�&d9=��I�����#>=D;�<�������;�̀<b�,<�9��3�����l\<T�n=ʤu�S}üL4]<Ƽ��=����k<[i�W7��ؐ'�Fh�<�T�
2/;}s9<&�+=D��<O�<�w�;-=�Z׼�b�k�+��(3<އ2=4컻f��I-x�������L=���1^���	�Ցs<iV=��J�s&L=/V�;|kD<Nb����><��<0#��l鰼�Ip<�ľ<��< Ld=>4����ӼnS�;CO��y��K�O��A�;���<��ѹ:&�<-�=L��<A��,�T=��K����;-4+<����3��
���<��˼�n�<+����wƼS�м鼒�%=A��<�֭���>���ݼ�SZ�Y�$<�P(=���~����ͻ�g<��<Pq<,V<=̇����<x=>��A�=��Ӽ�o?��<��2���!<��;��=�X=ѭ�<��e�(�E�%�A�<���p=֦���'���=�f��o�;���	�[�m�R<�W���P�;�mv��t<�6F;_$�=Wp[<A�A���r=�׳���e=6RC���b=�d��nJ�Z=���p�==�.="��<�;��mE��o\<��(��T=�q��-�|<s���-EQ��==�E��iZ�L�����<e:��l���Y=�<���<b˼����`=�=��ż��1��)
�b(%��5���[��ڻт�<�e�[�= &c�%�����<8/�<B�2$=��3�N�ռo5"=��໹-$�C='K���W��ߞ<���+=u�	��o=�g<+s;�#<�c*<�s��M����<�6R=n��^�U<�7���T=�����{=$�L=��K��L=����O���<�Z.=�=T��k���2=����Zμ�,�K6=]��2�?=i1=G��p5A�b��<^T�n�;=��	�F6=]1�>.=y��<`M=���;��E���
�Q�9=	�8=W��� ^�i5�0�6�_'�<g����<(�4��J�;�ﻆ�:=��i�s���&�K�9�R�ټy=G��?=������<�w$�њ =/|L�C��<�HK�UbG=ěT<��<� !�N֍<�_�<��<�Ɗ<Hs�<7k~=���D�L=-cĻ�B=�b< Dӻ��5�
ix����W�r�Q6D���t=wK�<��7=H�=��<���<&K<��e=��>;6Eh��C�<�'��5��y\����;��<1��;��җ+�����˼���<ơK=�n���W���;i$(=D�=�$=��</ϼ��亖�>�X�;��&=��<؍�<�b�<���<��=�����f�L��<�.��v�����d<ixz=��zw���T����n�[=~���_��J^�<�=�=�Q�����:v�Y�$=��9=�q$�
Ab<ӝ�<��W�E�}�؎�:�u����<��ϼ�W�<���<���<���f�P��J><��C�.<��|� $�?ܟ�غԼ��ʻ�.��=�V���J,<�76�ʇv����e�]��S���I<����l�O`S����<�fb=(7X��=��<k=4<4�~���뼫���o�=vc$�f�f<f�<a�,=-�"=�ox<P��ߙ�<B��x��<� �.�!=��?��F����;�� =\bI�rU߼4��ڻ���;*��UT=X&=f1�H�[;;;݉y=aj=�����r*=c�r�d�N���L�1��<4m	���ӌ�<SFl��Mּm��_C�@X����h���'W&��ve�XBj����;Շ��§�Nl=�k-<��t<�W���{=��W��^�p$��v��=�p� �=��=ٍI��I��q'���==�:n��|���v;��-�~	�W�;=,��<�NX�&1=�!����h��H�6�=��={����N<ƙ{�ZI�9E�h<�麼�=�_3=pƚ<�C=��X=T}<9�:;	�:���;��<��v��Є˼?���i �? <rC=����b=�����-<4=�ш����<2�0��<�><�y=0�!=f"	���U��^׻g���f�=_F�&=CO�;��=�0�<h��<���ā%<Q����w���V=��;<��<�ѩ:򗋼�mf��%s<���<EJ�'���EL�e�c<�ό<r�X<�0�3S=�������<�����+<���F˼}��LϬ<D�<�m1��u==��<�m���=$=}�<��a�8?<�u@=r��<�U=�.=�H=�Ğ�m� ���t<�=��F<�|o=��<D�M:^���иa<K�=��<VZ��<.L=��V=�3�E����N<�={�"<���<�,��5��$��_&=7>==�M�<�Z=�?-� �'=y-=�ww�LT�< ʊ=o^_�ŔY�+�=�#z=�{��L+=�I�VI���c<�j)=��u�f���Ӵ�<x�)����;�!���z�d�V�B=��D=�2�l䙻y^y<�O��l��r1;�=9='4�<�RE<\q1=��;� =T='�=��<�}=�&��<za��.�����j��D��zd�c[�U�<Z|�O�K<�֫<�\n=���kS,�k����仟.�<2���k=��Ǽ^�ӻ��G=��<��ȼ<h=T��:�=D����9=L}���]O���=�o8==2�6=E	<���<)P���c�{Ţ<\�<���ɼ�ϔ�7�<bq�<�;X�N��<��<Jl<��=3�L�z��x�`=c��:l��<�T{<Q9�q�r<H`����RF8���q�?�g=�O��V��$�1R�<���C�r=[(
����h�=��4=
��<���<Iml<�zz��!M<ڦ@��[����d�p!=#�O���8�#�¼����71=#{ϼ��9��<W��`lz=ׯi=B��B����=`�r�C�*���8=ɬ5<o���|'��+>=��o=4#��)(�&ٴ<�j=%A�<���=�='1��Y=U��<��	�S���X��<N��^��<c���mRo=f��<�CP=����E�먻<���.׼P׎=�}��Řɼ�י��PR��?���'���)=��H��A7�V��<X���g���<*�)=�証Ǡ���~Z�$S=��%=X�<��)�����`���e%�S#=�޼~3�H�u��2�;�_���k1��A<<j}�;3��<�ٻ�:=w�1�B_f=�^����;��8=�/!��YW;��Ҽ%���y��;^X=Ǖ���-<`��s���Z�=��<q<�j�Z��;�g2=풑<^EL=.b�H�=S�:�+=x������rļ �1=e�b=��=uU��v"��5�<�U�!==�K=�y'���Ӽ�On�',I<��+=��;vo�D�G=�������������{���jK�����Z&�v����}S��.�<�.?�pٌ<��9�Y�85@Q=U>=�h=�R�<�&��8��<�-��t4<���滑�=<��4�*�?�Kn'�:�C��xE�u #���z<��i���g�}��m'6<���<��=��i:=�[����fPx<w�<.#���T������\�
�<�2\�9��<�~F���R=_�<�v^��)M��YY<g�^;3J��E�<d�M=T�=tr?�����{��h��8��<��ֺ�-��%��v��؆��&�;Qu��\�G�S!`=�Q�5Y*���<�U2P<�} �D��;ދK=؜]���$=��>=���=��D��l��b�n=ɂ������,C�<̎+�eA��8g�%
d=u5<=�!�Ƞ<�v<s\,��T�<l)=��:=x�G����<���<�J���%ּ��K=SŃ=�k�<Yݎ�7�#������;_y�<��5�ُ[=�;���=	�?�]��;���;Ϗ�䍽��<#�=ǽL�D(5�.@%=� ����<���<R���%��ə���<�k�;��9j=�j��������k�ռ�n0��5�<���;Id�=)�C�Vd�<=��<��H��ƈ�����=T�<���<qeB<�5���lG=�="<C��<���ӋQ����<&u��ی<xb�=������/���@�O3�͖J���=�e8�D�o��(��V5�<��M<�����榼Sl�<5�H;7�<�	P<������P��&d� B�;o/���x=���<;���=���f��<��߼Uv�	�<K��<����Xf=2o����,=�aC��W=�F���<0����-=
V�Ά�;��=#.U��>~���Z<t�7=�����=�+=��!=o��<����؈e�������E=�@=��͟A=q�<CW��s�Z��tk�G�a�=`�a=��<���xJ�ynV=/̇�[1���=q =�I9=��a������̻m�\���=iq��9�}�f�;^���t����h=DP<�T�xW����<��<��q=ݢ߼��V�)=m �<�"����+=R'<i�(��:<�8ż��=�0�� �;��6�}5J<�]<t�^=֩���1^=r�O	D��]�a]׼�L�𢡄;��:�F	=f�*�ضҺ������;��<��7�`d���`�X�I=��"�z����5=W�һa��I2���1����<s<=��B�vB�׼|�X�	=� 
<�S�<�\= ��:~���{�r���A�{�=�i=QL=k�= &*�g��;� �:�_�{<R������<�X^��[)=ՠD=o�=𹊽Fd=b�6Vu<5@c� &��b�Ջ�;K�v����<)�D<�T�﹬���}�sr�ՆB�Pf	�j����<ae8=��~�˚I=�Q�ۼ��M=��<Jz|<Cx�<�l����z҇=~����$<�m�<��;��:��<�v�
�m<�jz��_)��s>=�]�U�h<��=0��<�ͺ�=�t�=��\�<p�<�Ar=��=/a����;��=cʿ<)��<�7W=�~��u=N3��gc�;Q�����<h���Z���e��<�ܞ;�u�ĽA���=b,=>��[#I=�<��!��'=�9�Ph=�Uo��<� j�`��8���I=��;=?+��k3��~�<W�<�+X��8w=B�f=^�p=�'���"���<&��}�+�	�����=��%�_W�=��s�ռ/+5=�)=��5=}K�<�r����<�{*������:�<Q6k=isr=3�߼�@=��<9�z��ҼF��<4����; �G�D���zP�/a=\2E���)=�k.��� =��q=4� =wiM<�.�<N��<�=�B)=��<����	���Y=f�R=��(�7=��=˄C���<O=��=ʵP��欼��;�5<$�<< ��`;=2����μf<���<*v6�_�<پ0<C}ļ�I�<��=�0=�Ҽ�c���;\l�<�<<!�d��5�g�=�3��#�;�r.��8���<�V<^��<H*��
��I=��=������\=mz;|��<��F=a�M�Oм�<g	�</x�:�=�Ӽ�?>�G0�A(N��*d=ێ�����<J�E= ��93=���Nuм�1�t~ܼް�<��+=�(=~	����f;E:;u]=����h(��}���p�3�5s=�DD��N[<� =��S��K<{Q=��3=Ɠb=J�̱_=�;.=av<0�H=�⫼���O3��A<���;�P�H�ֻ�%�a'�h�=��/�~8���=:J��*�<BLa=1E��؆;��<��;V�|=�7�
ˀ���g=m�P=0���G���Ӑ�;�5_����)q=0�M=��
=�-��=m(c��[=���<� �;�����k��f�3�Ɩ =���</u���=5����{����<G�$��;�Zμ3���w��������� )=)r�<�;;�꫻�A<���<��8=��0=�#f=2�����Fm��D�<0��;uP�;�L�<B仵��<0;5�%<�K><��+=)�z��rK�1������q=u2M�ۆ6=�u�<G.ѻ�U�]�h�>��<GУ����,q�K)�h�=X��&�m�3~��@����<���;H=$�5<?����<���<�C�:%�,����=� �<X�p�{.�<74e���������&�K=]��<XC�;�]�<��9�[��:ͼ�:]�#�=h�5=A0�<�mO=��J��k�<W����<����K�i����҅;}3���=�Gl<gg���7�Uk���t�<* #��l5=|���)���=ϕb=\��eה;f%�<`���m����;����I�_<�- �%Y�<���,�=!k	�o﫼�ζ��
.��e1=L��<c#�<E�"<��,=]��<e0 =ЖH=/U=^j�:�n�;3����N4<Ț=(�d<��g�󻸈�<*^F�S�;�\Gy�9�o��Z����<@�=S7<��<��6�r�W�<o��<�Ҽ:�白1�=�/��h<t�	=���<�9�<|�żvX<`��;�
;F��<6mۼ��"�-�=?"</q<�?����-=�+1=n�#=�\=>�3�
��;/+i=DX�H�c�%��<b�6���`=x�C��F�<c�w��/I<ݕ�<#	�<~z1�;;B�=<���N=�<Xg|��w�<��<��K=/?��8=�9z=���νH��f=@���
�\�/�����<�"W<$��9IЃ=�}�<;o�M��Aʼٟ5�I�9��q<�w^=�P=�^绑�p�����ls#=.o1�t��!`|<�c��k���Z+=���9�'#���<f��A���3�)Fk<��t����X���R�<�s��cm1==KE���a=�n�;P�/=��G��=N�
�bq=��5�)�:�j�7<g�<<�t8<bZC�m�=������y=:&<ٺ2��s�<��,��<�E���Z�=�2�-��
L��%8�6^��bLE�g�L#���+=�[s<�A=(�>=����vXA�6��<���< a<Qw*�5�ʼ��J�{6�<��^�����/�;��;�=�
T=[m,��T��`���=\&=͌=�š<�x��>�����@�x��0��O�x<T��<�l<C�7���<U�:=��e��oe���'�h�<��1=��(��M@=��Z=z��<��k��@ɼ��O=�0�<
m��o<=
x�]�==:�(�{{c�%�|=�y=^�:��!��/Y�׵�mZ��5`�=�!��&_�Bۼ�jX��G=}܂=5`�<K�<~�X=�Fٹ�f�� *<�*���<�C=��:=����#��ʹ�<��?��2'���Q���2<Z�N=�c�؄0���T�*��=��C�Aw��-.=��=�]=񒻛��< ��<�/d=�(<=�	���;�˼��<�ES��乍�T=�S3�6".��M%=w��;;L�<�Q"=��=��<�H=�_=�8s�?�^=5Ƚ<�<}rt=�=��2�;�;V�55�<0鑽�F)=��%=UՁ;Q�<5T<C��<+4=����r��Dm����<��/�M��<]5=�@B��B��I�	�F�a=������R�j�8:�r;t�
��Y='�W=@�W���o�'灼�J���6=7-.��|c=-�J�MՁ�M��<��G=è�<��I
U���z=���'���~�%:r�)���QO=|m�<b캼�\4���m�aꜽ�$o;,�<q=�}|#���&�,�<}���f��䴼$mf=�N�}���j�<�M�D+�1�,�,R� ���j�����<1м<����=�gv�u��:LƬ��c:�(�\='P#��7C���<0>O�v�<�=+�(���.=U�ռc#L�Y�=��1����<���<�A��'�:'�<��n=��=S(#���y�i�+��=v2?�{<$~��񹼴j�<m�J��������<��z�ט���W�<�?���<�`�<R�
�w�=b��;Yq=GA�<��m�a��<�.@�	����!;���<@1<����<	�9��=Z�N<>c<�H�<��=@��Z=K=� t=-�<�I�<΀ջ[�s<\���ޮ\=X��;4h&=�Q�;)w@=��M�|%s;�����=(Da=��<s�f��f�U��<:	F�<�=�qļ��мŪ�Y�<�}��C>="Լ����U��C��3�9�*=�=��9�:K:�<��=!5=o����ʄ<��@�s������d�C;bǗ���=�<~�;񮦼�g<C�V�<��S�=�j���d=MZ=�¼MV�=�й�f����]d`=B��d�;.1漌zT��%d<7I�����9�<����h.M=[=����j��<h���|��<Y�:
�Ѽ�t������K�ܣ��^2�(;�<ͪ6���,<�����˻�2=�T���:��H�<����5�;dh�|��ϰ	<RDͼ�#�2��<,ij=���<�FE<��w<�)ļ.�'=�W��<^�f=g瞼X��;��R=�m�!�=�!�;2ļ!�)��<�ܹ���:��Ȼ�{c�o�F���{C=�<�3��<�,���d��T<]Y2=_7=���<�lB�m=F��<cA'=N6u��̼o��<l�(<�Fy=��=j�<2�<��/<bc����;��h�h&�<��D�A�.�
�<7�%<��<"���s8���|=DwN�^�U�#��<��b����<뢕<��^�p��:y��:#=�1�9/=
%l�-���c�<��-=��]=aS=�B��Z�'=�b��(;8=W$E��7=t,�H�=|S�=��:��E�L�m�% �<o�8=EX�<%�<��a<L�輧��: T=�o�%SK��k�7�����%�F�)<�5*��!��jm=P�n��o�oi��t�=�=h���Q����=���Rt�<�<��Y������=�4=3������z�<8';=��=F����iX=������<ެ�۾3=�P�{ŕ<ۖO�����*J=hػ��k=0z��(<�ւ={�'<�H=$=ӷ�<�}=⍗�LƼR�;S�}��K�<��U=��V=-y<�Q��̼m =��"7�<CAM�X L=����6=�
���)=m�<<��<\C'��9.��>[�j`�����;d�����<�;ck=�qZ����<7j�<x&���z�� ��O<f�,=_-Ƽ��F;���<�� D1=�CR�́"�gQ	=�ϼa�U<Q�4:K[5=�ʟ;��;��G���h(%�],Q�B����h=�'N��(a=/*m;�	����:?��x��G;��^5��,���vA=�7>��=S�u;��<��I�5ib�l�=)!�:i��<.=Ӫ ;_T=����,�@=ӌc=�4ʼ;S/=a��<�!1�
�=��U�r�c=w��^d|�7[Ҽ�<1(=7=1�e<�
��2Ӑ<aH<!U �	��;E�4�\�;�?-�=��|=�E��t>=Ҷ=��=�e��d�<�!���ݼv�¼<�9؈�<"S-�?�(=�sP�gԂ=��|<��<џ�<�[O�c+����B��<��==��2R=��<b��
={!=�_�<���<T�=�>�H���B׼�~8='��<��u=xj�F��<=�0���=�=`[+=i�l;&;��#�;P*<{D�v�i<����Z=�-/=7��<`v�����<��S�gwa=M�:��ͻ�d���s=qq�<��Լ�%�_n=<���QB�b�<�r�<]��n<�]=Г�<E�컎���.���4�7k��nO<�g0=<=l$,�+e)�� �9G=�E���}=��5����N-y�y�����A�L�p�����><u9����=��Ǽ�S<���:��=����OE��=@�\<.�=��b�����O�=ࠋ�`y~�y	�;f�1��y(=M2�|�n��׼(��<<��<M�Ӽ� ����<��;hD)=y�׼��� C=�3�ux���7�;YмMy*=Ξ�:Ō�t����c=̌�+ =A�-�$n�<硼��0=�5=]��<{����ܼ��ȼ$��<9��<O+�<P�"���w�y�����;<�<�
2=(�/=�U�<��<.��<d==8���Yl�S�s���&�O�)��<J��'S^��#=|��<��=ؑX�f�<{���[E�!�<�O�,mм;[T<��<"k����1�=�R.��֥�\�=����:f���}���J�2/=�Is���m<	�_=��#��𦼍
�=n��< =�GO�>]=t�G=<#ȼ�-z�/�*<��C=�!G��/�S=���ҏ�<�x<+15�n�<�%��;�3=��ӼI<ǈ<�̈́��
=����B���R��2�w<Q?��ª?�!G�E;f=ةl=����F�~�;R]�B�E=����5�=�=�9���U�"��<��s<cG�v�C=�7=8�)=�I=d�ռ�C=zm�NG��Yȼ]�.=: ��&'=��<�S��gP=[&���R���5=`u<v3�<S�&|(=�{�UO��'@H=��ϼ|1�<��=1(���&n�D<@����y[=nԡ�<t�;Ζ�:#Zj� ��r�?�'�����
;c謼��׼@٭<ޛT�{����NB=	�)=)�\��sd���H<�
��q��d<Ҽ�����;V-����2��@�=�%��9o�������;�
�<;�!�9��<�F�j`X��2�<�*x<���IC��:h�;����=��Ū=�+ռ��Y=�y&=}$��ބ<��-���@�.3Ǽ���[l=��@<B���n="xO;�����ٹ�:��<<��>��<S��gj<r��޼^�P���w~z<v;���J=~xg�؋�C-
��9���<r��=D�C��<���<8N0=0f(��=�ɞF<ƕ���*=�QF=��=��Ƽ�4*=��<�C��<�=��)���<�����.�<�&��<�Ѳ��K��M)=S���P�켕��<�3�#�B�ȸe=YS)�#��Vx�<di/���V=N�<Xa==N-�<�P�<%ch�����\JL=���"��<�B=�=��4�^�g_�h�=�c!�L�n���)=��;�zV=k��k�ʼ
�1��T�Ё��iE:=�敼�8ʼ<�o<-I=�� =�輼�����=���������1�<ȗ<��=�<:X-=F�|@���=���3�7�	l�;nP.=`�<>y�ơ
=���j�*��M��3��[Œ�Y؆<�Q˺�����%���C���wW���e=(����;�������<�k���vD=C���eq�LC�<�v��.<��;�#��|�V=�7;���~�X�=�O<��.=k����<=�]�<P1N��
<=�/�<�}�<<{S�þ�<y~=�t3�TW�<Ã��C��;�}ʼ�
5��;�1�$�M��<=(={!��KV���a=M#����͐=aIM=�.|=��f=a�j=��"��üj����@=�c$=��<$ѐ����<�
��|�<�C=���T��;�����;I
�#b<���jv<��,�CM���.漫����=q�<�]�<�v5�ݤ=�d<�w<�V<�`�:�hƼK`ռ�<�D�=�^w�֟!=<�a;���:�H��~ <MX���l=�S���o^� <��#��W@�Zu���l��=T�~���3<ព<^�ϼ�X=`ZX=ٱn=��a,�;no$=g�<�P�<l��<�7T9'ۇ�WQc=HkF��xd�j�`���<8�0�i<����{�<��	����<T�Z=E�<��C���,[�<7��<�n'�L%���6A�V�c<$43��'�<&�;tc�2/=�����e4;�A&�a���x;-���_Pe���H�0>��d��Q�<5��;p�����A��s�;��v=Mk=+�v�
L�˰";���9�_�<�	��hq=�L�<$��<�!b=b�0�+��&�Լx;���=7I<��z=LC�<�0=�8=r?��:|H=b����1q���I���.=�X�\kѺh�ļO���mH9=�ٍ<
��<�rټ�b=��Z�N�:<���O��7^n��.�=��<��i<�\�:a��K@E=�4<UO�<�<x�ּ*97�����tl�<=uN��=<�!:f�ߡ����T<���<ߩi��ռ�IA�0bϼ3wu�H��;�<�D����|�<�Z���<���<0"=ck;��������.��P'=�R�����7�<��p;�0=c|�<�X=;t�<5ɟ����<��j�������	�Cټ`(<�=H�H�F���a�<�:=˴<�=� ���,Y��w�۹��$���3��9~�┦<-����+=�b��V���}����5����|?�<�,=�5;)�H���?�����E��H/<���<��
=�_4����ެ<�3�CC#=�@�;���.8W��5�;�P2=m�t<�Yx=���K:-��&L�����=���Z��<t�<�jͼ��7=��8=FЙ=�]#=�?L��X��1�<��C=�HD=��;�b��h��=�m�=�~мm�"����9h��<}(켾h2���F=81ռ<���]��` =��l<B⊼7�w�v�C�-�8�
��u�j���oe=��w<#�(<�  ��q;=�}2<Y�D��N�;�����ho�%��:D?!�!	.����<�@9"(&��kx=u=����	=���:G����;5R����m�T<.���AP<�z�����<�@Ӽ���<��"<�͞���<�	@�{ ���(�%���g	�����]�=��=.���!,6��^R=��=�D�0�ӻ!������w�c�:C ����<��w=)�Y=�D=�^N<�.�W=hn=w+��EJ��8=S�{��DI�-�<T��<�4X=�10��q��^
�<C`�#?6�Ӳ�;�:�/%=�1d<��A<G 4��}H���6��SJ<��]���=[���	���<Q?����h�vm<J�ջ�Å��Lg�� ߼�t컟iR�-B�<4�<�q�<�t%�×=��O��3���=�Z=3�$%�á*=�r��1�<�.̼�&2;�,<%7ϼ�{]�;r=�Eܻ_�{<J]0�>�<I)������ =��2=��#=��^=�	K=�
����&�W�:�h�h�C���ۻ�v��N&���=���5���R�&=��*=��T�v�B��,�E�c�Cv<70=;�+=��?�B��<X?����z�?.U=�:F�Z@B��q"=�0<����3p3<�(��\p���7�?�N<��=G�d=���<d������>�G炽W,~:n�=��u=��v�a��<�ӡ������<���<�v��>^$<�J��6M=Ե��K:��"=_F=Q��:��<n����]��o�<�l==��Z=�S=@���;��μ��D=�^=�y=&�1:�����<��N��QK���]��Ǽ y�a�_��<E=>�e=�����+[�6;�<w���Ż;��^U=��=>�����<�dX��T=��e=E�4=��=	&��Qh��*�;`*��Os�K-z��=���:ޮ��Z�:=��>�=<6�<ω�<{œ��<&=�J������@�|�j��j^y�Xp�;�_(<��~��LK=�: �ڳ�k)��*v�:AQ��Q�:n���_�<�ݍ�i5=Ϲ�<��<��;zҍ<��<-=���;�{�<�]=�Q�o��<���<��?�2(=�2L�x[��d��A;̶M��G<�O����;u8�<�˟<�on=��T��C7�.�v���<~��zT��ju���R�1�<�z=|�<�<ܼ�?�;��]���<�ӻ��{=W�<�<����r<�;mvk='A(=����m�=-��<0j����=���<��t<_�H���j��ߴ���N<�\X<G���<ޗu���@=��V���pL���;�8�<��ʼ�Ծ<��'���:=绋,���9��4���V=�C<�a>�Q9�*���F�<�:����P:�e/=X�=^꛼h�;�%=da;=���<�Y'��{F��	���鼝�M�	+�=̖��H�3�[W�;rrH�<��<�0ǼI�c=@��;D5=��t�� X��l�<C�;>�9�%��<�o��~�:�U/=�v-:��%=J&=� 1�m�o='��<�g;�&>	�}!�S�
��^ʻ�S����%<QV��ʧ<�tO=����咼������A�L層�U=>.����6���{K�M�=�;���8=M={k=��<<�k��a3=+@=��I<)�:'�6�HL���ļ;_�(=���Ԡ
��z=�u#�!��M���+y���`<}��<VK3=Uz����%=?�<<K�`=��g��+w�C|�0�"������/�l�2�K5�<�ʼ��U='�����.�&=�j`�
�&=�F�8��pJ=����4X�;cb�<.7r<\�b�7��95��݋�@�?��L�<�C]=�2���;�v�<P�r<��D���\< <3_���ϻ��7��,�H���=坸<�̈́==�R=�c=�W\=���Q��\�~���X�3h?��5��Ҁ/���=��=傽����<����P<A%2�&"=6��<uv��JR=4�;=�ͬ�+�	=�4k=p�(<D��m�;���=�n#=��Z�Y��G�;f�T��m<^��b�<�-*=�ZE=�>R�(m�<�G=�W<��<��ѼU�|��.׼Q0A��&�ڋ<2�ѻ��+=���.�;�7����l=A�'��Yo=��L;�?=�ֻ
�_�5<�]!=�����;�i?��侼ų><�!ۼ�.=��o��=�k��dS�KƂ<-~���[���r<��<!k��}'=�S�����@';^�F��2��c8/�&��<2�2=�	W��3�<d�C=ko����;j�<e<ԇ��K�$=�:Y6%=+�P�P>j�'*==��<����������L��U=$b�F{]=�W�|=�%�v�=Ļ];)��<�-=�:R=A���G̼5���<-�=�5x��5�(�t��Ƽ0&�<�`�:�͸<?tJ��o9���5:&+0=
���ȼ�.<�^n�;�G=tǍ�{_�!.=��h����<�A���~;Ŵ"=�"K�ՄL���<=u�2��o���'E=z����Y�v5=�/��O���j���<��4=�Kf��B�<<N!�p����9=�� � v��P��\�<�d<	�C;�^c�ĩ��ڙ����̼����UD�V�����1=��;OE<�X�����]�=v�</ټ >��O����ݑ����;ݢa=6�<�M�Ʉ�<�C����y�0�e=�A�<����",=�Ӽ�_�<a��< ϼl}'=�6�<$���=-<3���E¼��/���:<��O#/=-�=���� =�u{���%<�GF���ڼK==�<߀=���S� @��"�w��<'b�<���p^n���*=j�E��z�;8�}��6\=��1�,,��v�E��|���KU1<(�G=P���q`=��f=*�-<=<.�<0=봳��dx=�A=���O%^<%=Y�=M`	���+<ʠl�R�-�o�P����A8=�1`<yt�:P��g1D=����:��sA=�����ļ!]�<�T<%#(�Yc�7D1�����ĝ;�zm���u���=�D=9~�<N�����ɧ:�];d����H�_�w=(E���Z���zL=+�=DQC=�b޻o�5=<�h�Ų����R�M<|zH<7�<����F�aJ&��<��<���_h(�)8~���!=�a3�m�F=+�4��=
�<4,<@�6���O��Qc�B��<U�K�|09�I�=�Y�� ]��J=��L=(D=
u�<NT�<kWg�v���g�*�üTC�ᛳ<N5 �d�����9��"l<�HZ�Pm���3!=��<�-l=ǼE=��]���[:�j�=Ku"� 1/=�X���F3=K·���1;f�N��3;��(�Ϲ�;��k<���j�<{�E�,o���F�W=v��K�s<� �<@�<1� �v;[�
����In��=hx'<�h�b���B�+���*=�%<s����=�A�RZ~<Y����yB��MC�9=FW�(Y ���R<�j��4#�Ĥ�;���I�ͼ2U��婱<�s]<���<k(=���<X[=6�=��J�eI-�X�	<�_7�`�<�8�=L��<��<
�~=��B=�>�:(O<�A����	���<�b�;�:��M?=o`<c�=KWa=�!޼V�=05���7�<��S��̼�rw�($�l7 �ܯ=��<5Q�ت˼̱�<�	&��¼ЄS��N>�ޝ*���O�U0i=�:��ķ]�r��}�9�r�-=U
_=�=��)=+Ĕ<�u*=�v#=�7="#���<@�=.E��"�	�KK�;x��<t��<^6�����<�9=�d���:�}����ûҷһ!Ǎ<�*��y�<��<%�ļ#�Ƽ?ާ��_)��
;��J7'��(Z=U�`<���<���|vt=LKt�0��<鼐��9�`:=�W�Q�p<�� =pP�~y�<�+=SH��_��<a�;9j�<A�������m��|L8;N�)e=����Ÿ���V���=�T��F��.���M=2l�<�@6<?<�;DR�'��<+oZ���:F���/=b��<svR�r�e�B!W��(=�<=T<%;=��4<�e��f�<(��<�\ܼ�%C=ݢ=��W���żM�H���mv=�&=����=�<�J��m+`�j���$�.�)2P=���<s)<6�<�-��=�w<���;�S�X<$�"���=���I���r��^"�;�%J��pv�|j�s:=�o�<8�d�����v��/�;�R�Kzm=�CF�N?�;]�;�#=tբ�[��<�� �$=
�r��2�<��eZ=��<%���uX�<�OU<�=��3=���0ƛ9�L��j�<��5��.��� �\�
��.�<��Ⱥ*>��]����<�,�o;�A����<bk��@"=�Kؼ��M=Y�=n�=y]޼�ԏ��Yr���=_?=٨<Z`� .;tw�:=��"�
�"=ޝ��&<��|=�#O=� �,뽼=�<�!U<E��<o��ߛ2�@��<�<=�]?��u1=���Q�c=h�=ް�<ib�&=��H?=�&����=���<_�<Ff�k`#�s�<�Χ��Q=���ЀW=g�c;$# <��%=Z&B=���D�u��y8�%��<	�=�8�<?9�=��D���<��:P�I�KO�|x=yD���'=���	�;�{�<|L^:ha<�u�<��/��r<=#F��0�Q���N�<.�<�x%<�~=����e��Z$��Y69������<1�F=ʮ�<z�j��Q�7�E�D�W=��W�v�K�,�?����h�Y=6�i=��V=�;z����;�=q\�����:�[��>[=�L�<����b���c�<��H�vZJ�
���VL�Aa�<�c �^�\�]�R�A=�2�<�Z���;ټYԼ}�<G��{?��ܼL�Z=*��H<��Da=�*:�u�=x����4w�e.3=��U1����l:���<�9*��
�<t#i=D��bO󼄫�VrQ=P����
�?"�<Tr="��V�1���K�V��<��^<v�H��LS��]0=`�r��؅������:��ݼ�N3�n���|������˒�r��<8 ��bJ�J����_��&GH=M�h;��=�� ���Z=�7=�R�;`�=5�<]�f���<Qcg�E`�<
��;W4���O�ޓ1����<�\�tЬ����� ;+b�QA3���[= #<��ؼ�E�9�4v��9@�eI���S��_��}��1O�;�����<��Y<,Xo�0�<���<�02�w=ӄo<<=D=Qr����=ӖU=ȟ�<�F��=u�&��Ӵ���=M�=����1�<)����bʼ"=�%�<�gf���?��<'�q��.=�V�<xzH=.o�*��<Y�v=��;�bk�gQ$����<sW�����J	=��<>�H4=�KM������=�a<��)�l�N<�t2=8�N=8�1=��<� D��1U��=<�cj:1=af����\꼑~3�ı5��lY��;~�=�|�&�=@]����<@�2<�_�<GrӼ�Zu=�\>=R�z=�Ca=<��<5=����<�.��>����d=��e���u�g)#=	+)=$ =H�<�:<�m�<a��<�F<#��$�;������=�.[=yG�<Ѻ>=_ *<��<)�ĻK�Y��D(���<<9��ˆ<  ;���<��<E�<z悼�bP��w<{[<	٣�^�w=��<�K�ΥѼ<ܠ��,�;��i=�϶��d�<I�,���M=�b`9���<��I�~<�Һ<�+���3��l'���y�k漬tQ=_c���V���;נ�;�+c�(.o�_����J��n���L=�.�<�]^��&]<��H=c�Ӽ
��B�=�	I�<�֚������6=�=��缙���o���'�:=�w�uʒ����<��V�Җh�<�H���bJ[=���<�	ʼ��;�w����=F�L=C�<������y�>�żj0= F<}������7�k��6i=k4F=����-N���='��V@��gD+=��&�Rd+=F7�;�;��C����z�q#ϻ1�)�V�ռ��l����c=�M�+��L =nW�yZ=c�ټ�|���y�=���v��;");�i�<���<�h������󺜑�5�=A�?<�4��"0�;���<T�;���7=#O[=��6=;kڼ>�m�'y�m4=Q�X<�,���ռZU�$�	_0=ڈ4=�GM�O>�J(=z��< �X=Uɯ�w�
<+@�<�l�e�<D�=1n��T=~(ǻl>���'��*�6�%'{=����ڷV��W���@��O�,=.��<�w�<D	�� d��|D��m)=:Vƻ�E����<jv=��;)�H=�c���l=>��ּ��h�	�������:�w��<��;vR��a6�Y�=��c=v�;��ڼK�4�s�==��=�L=��U<Q@�<�t�;iD=�.=n���P�<�y=���<�
<�WFY�0P�������<���;︝<j����Ǽ�&u�R����<�� =��)=�+l=��o���"�ϫ =�ڡ<$�#����H�����<��SӼ�T&��N�<�*������=�=.�=`�g=��+=|��<�a�<c�z<Hw�2C.����<�R�<ոH���R=�%U�ّ�;b�==�J@�=GûYTs=[p;=US!<X�?��D��t��; f=TԼ���4�=<�0|�q2�{��:�c��-�;r,�<��T��&f<��=�\@�3�A�@��Q�=�^+	��ҙ<0�=�� J��D��<��:=�g�Pw��ʰG<*�󺪪��TF=�x)�Be�=ι�<{[=v.�=E_��	=9kRļ��R<\g�I��<^+Ȼ�� ��C�;���<v�8��2<��,�(� ==g�����3Ė<�O<=��=�NV��X���/=�ho���<��;��;�����~����<���8\�<=W��:�!d��E=����Frɼ�p=єi<��=2=pKB�2�$<�м<��O=_i��R=H���q���E{��'�<A�Ҽ���v	�<��$=���K��;U㼼I�����
�+�<n�x�W���&�L�9�%L=僚���h�n���*:��V=cF|=�F=(nܻ����ڤ���;�l�<�b�<�[��N*�x��Q&�<�{���S�X� r�(E�:���<[��<��]�a2=A�]�Үh<��<�l)��<����g��'8=���<-��<5�R�:�ϼ�ތ��/=�<�	[��菽�\���B���;��=�w<)==_S��<�I�<��(=.�M�8|<@��=v�y<t�<$W`<��<Gɻ<G�B=+9���컱`�<�c�H�<�5s<8e=r���To=M/�<_�3=��h������<��}�Y�8�h��;�n*��C�<���\v�~QM<ۺ)��7��\������:\?=-^L��TV<�0r<�-O=uvM��cͻ��=�u���=n9;��T<�0�<�7��SK���e%=qv�<g�o�4=>�!=��"=A��F�z=����u�>=��e=��]�Ӷ���k�>c���(={5=Q�����r�!5��]0=����!N<� �:��=�6�;�&�]�:;�/<����!�@=Ւ%���:������S�λ9�9����%;%/�&�<ŏ�9���J�Z��"��H<�B�"�{"M=B@�<�O1���X�x�A8�ڱ�@��<í����=�?g�,��~ޘ;��B���$={0�<{:L=ǶY=�=�m+<t�4;�^�<�;"<C�1�"��I��q>N���޼�q�<��d=��)�@ז<�i=�BF����<�����`=�!�;y�c�F$3��S�;K�3=�ז<85=�"[���=ӓT����:����2$���v=Y��� ���=zdV�m,���r;5��<�/�ؿd� �I�~w��ȩ˼% =�=��;�
.߼n�}�-����|e=;C�c|�<�h=��n�k��<b�'<��<S�<��t<�*.�;�=��=��u��K��z�<��@�r{3��A?=c��;�Ȓ<1�:id=� =;�<����Ƽ~�a=����z;=ts��uk=l�~�0=Ɖ�;N�b<�mQ���<�d�jX�,�<�ѧ<v�f��Y=��=JD)=��=�^��ja=(�<d��K�U=ke=�僽�@5=�l@�e�4=+pB�h:�s�J�!r ��:�<G9?�U3Ǻa�σ�;������k=�W�� =�xX���
=�7=�
0�E];e�/��Լ�j#=�JO�j���7I=��:
"�;?65�r�[�!%=L�]=�8$��[1�Ct�<�5<j=�X8���;~��;��=�3;Y=�E}=a <��<�3=�$=��;���1<n��JX:;z�=�l����\�}�l=�Α��u*<c��:��,��Qϼ��q=�� <Jge=�}��2T����<f}�Y1Y=�i�����&���%;�"U=��L�ۣ�<��3�C�����=< �a=��ۼ't���<��9���q=H���X@=C��_?=`�J�ݭ��@=�A�A[��P�L�h�V:u�jG =h�=�c�<I�z�א�<�E��s��:=��<q8���.޻�R�;%`=L*<�s>�}~z�_Xȼ[,L�&=�U�&�6}W=%R�:� Լ1X���;H��;[�$=�~�<*�O=���0�!=t#�2D�=�j�<U��<���%�=ﬨ�6�
�f��<㛏�w>=N�� u
�;�A=�8C=Aq=�)���;��	�L�����V��>O=���<
�<:��N�3��⺋��2��7�(=ڝ�<2�<�:<��OH���<�TP<ce�<1�(=�v���*�<�Q=_��<�\� �p�j��WS=�R?����<M7���<��wp�<%�2"�;�a�<�nG=��-�=����O;��x�D�ͼ�Rּbn���:�K��A�[$=���i�<=L�<�q"==1;t��;�jf<�*���d�U�m0<� �<�*��;���Z�;ف�<;�`;2�=D���ݍ���_=���<~;=v%X�qw=O���I����<	�&��|����E�	�b�xD»��F<��;j­�t�X��Vk������<27C=Ϗ�<*���W�uu���C=V�Y<�ⷤ'=li.�Qr#=�J=�Y =�V�= h,��� <���rw�<�L.<��O=S�=h3;<m'���)=��/��7:�2��m��hA�F��7_<>��<���<D Z=^��yT<*#6��A�<�=�<H�-�.=Ym�����ΐ�=��</�h��="����<�CY<�7-��6<��=��.��,ܺ��d�-�ټ<�,=@��<k��=���!���g���S�: ?{=Z;���$?�:囼vQ���;x�ɼMS��[4<�n��2�����aw��3]=�
N=f~�:*��;<xռ�Us;�+��3i����<<5d�TrA���!��1��d<��f=��`���<�@�<��/��Q�۞���<��F��n���<��ݼe<�, =#/;�q=�:�nz���"<�a,=��:����\1<�Ỽx�8�_~N=ʤ�=�g=��ռ�	Q���g�/<���<!�ռ�1.=�(���<g|ļкw�A2�<�<��
��x���A%=&g�<Ζ�<G�g��̭���<�o？����<��<��#�ļ6�������=Y&=�;��W͟<l�<9V=pxd��ȉ<ֵ�М�<B�z<��P���;$�I=�6�;Qd=HU<�=�a|��=�;��|���=M&�<�>����;ɚE�e�<�p=pD:�)�b���^���j<L5&=��=9��=��;��=V"����;|�"=�J=�[�<Q�%=��=̮�<H��{��<��</)�'`C<�*#��^���=��y�<�L=Qf:�br�t��<!��;��M=p�(=󮝼�Z��t:=HƟ<G�a�ֻ�<W�B=Z��<�M׼Mw�7=Z�B�,@I=���L�(=8F�բC�GW���u@:N�\���+�B��U�>Is=X�J�t$�<C�<S�R�e�V�<<t����(<�`&��!�<���T����:f���<��8=K�<Ł�<���<�#꼭g =v*=EM�����d���ռN�Ҽy��<���n�^����@	E��`p�@�=��U;��9=[��<�&=DtH�a�h;cW�<�ٶ��V��[h ;�\v;+�A���U=
=�;=�j;n\�j����<�d=�h�ھ����q�A������L<[���@*=k�V=��$=�|v�w��2t�<t7=M�B=q�@��[��ȤA���:=��k�;�ټ�u<'jp=eLh;jf=�3���Y���A�u�>=9�Q�r�]-=]�<�)=�����R=8��<�"=��YD=E�O0=���<������991h=+�=#{<O��<p�#�.=9�W����`\��V���3��-�<C��(�������~n�
����p���@=��j<u$4=��5=�T�Q�=�6=��*=�U/=|=U��Vm�;�h<�2<��6<̼L:=��Q<��;�����P�9�?<29W����<�fk<���<o��@��9.q����<�F<��@����<p�'=���<ÊQ=
y ���<��]�<e�<A=F�L=�B�<)<�z�<��0<��Y<7�%�v�;Ƞ�_GǼ.��SZ���9��1.=��*�0�n;r�==fI=LH���2=���<
���S=�=9ɻt{k��=$���N
��f=�w��z0M�I�����Z=�T��L��S�=���<�T=�=��K{ƻӃ:L�;�h���Uؼ�Ta��\;='i���K���=*n�eg<��<$B=a��(=S$_��H<h�켂�'<�����=4�9=cm[9����dJ�N<m'�;��ȞA����<�df��<<�T=`�<"�%=?�a=
=.V�&8=�۸��*5=��<#��<���R4�C�o=��s=��5��%5=S��A=2�<��T=o@��j<�@=(*�;�<�=Ȟ=�v�;J��B\��:�qt�<`�{���Z��p��m�1=Ut�<�^=1\_=Ȥ$=�NA<:��[=h7�<̋4=�h=�m����<��9�=R�9ȣB=��O<9�b=Mڥ�Gx/������?G<�L=ԓ�Ƨ;��B=�#��:��Y���%���k=Гż�`s<�����v=v��S�*=>5s<�o =XO`��A�>�$<��!=�S��We �5�������9�ƻ�=�-ؼ�&a=f�r�����Au�`��<Tv�<_x�V��;H�W=�N�<��p=[�&��� =��&="�<��=#�1=1�Y=��=��9=��=���zW=tq���1`�j�=l�z�L�����c����<��6<��|�����LC�<W顼d��<E�j��]5=�q��68��oS=mH���<Z*����x<�{L=��E�N俼�u�=U�=׻-=�K*<�!l<)6:���커9����-={�%=�>����[��]3=N���h=s��<�{�6�
=Qb<sI(=�<)㶼��k�X��to<:�O����E;*����ʚԼ��<l.��F)��{M=d�,���/�N�=X`����<����s5�� ���]�������N��/,�5�<��	=��Y<_(����L������
=��=+�D=O<�N�<ht�<�C�<)=�Լ^��AJ�8�O<%s#�L�R��g=�e��u�<���zE<x-�ˤ��^��
Q'=������<V<���v!=Z@=l��� O=W�9�M�<�{�<��%=R�/=���}w<B��(vV=2��<�k�<Q��%
ּ��W=�<޼GZ=�'I�B�;lc=��
��DY�UkJ<����3ﻪcH<m��<�~�|)�<`/O�
�;�hs�;���~M�G%��^`���f�<��,=�1�%=r��<Ȣ�<(�h�)T(�4P �{PH=��.<3�<�R<�Xm�*��P�|]�:��)�&���4<�*=b���<��?=`�$����Ʊ��ݥ�<��<��1�%v�;;x/���-=v/<y�,=�0�<Y�6=�o�w��;���<�����<���<���1v�<*X��[����=�J�</�������<C�T�^�ut��<E�;U@���K��M6��B�<�~M=9�C=�:!��[8��P)���O=�1�<�LP�J����׼_�b=0M�<�+�=�b�<޿�<�t�+ּ<?I�lI����=�`��{C<�v���:=W�ؕ��&<�w��l�<�=%��6&=��8�L�$=S5<�=~,L����n�<�t���I���=��V��@Q��b=Md��sb�<@>=��C=��I��y�<j�=�;C=�PQ�5��<b�4<�DZ<W09�O�ɼ>rn=G�w=�����Z���G�%��<�8�<KK�^4�;<=<;O=�*��^=�"�]����<u<=��=�Z�)=�8<��|�}V=��ֻ��X�%/��g�<\���a�<�횻�������_��;�ļ�ƻ�ټ���F a=CeT=�o�� =s&��|�Z\J��8q�C�45�=:������<[�_�+�8=f =j�n�<a-�[��<�r=������<i�$=�Hj<�ۘ<��0=��ƻ�;E6f=ޜ9���)=6���?\X��ͻ�_$��=�L=��Q���<���<��Z=��
���q���#=~
+�Ff����(=�[5=�@�<&��@��������<���=$oϼ,��<��F��R�<D%��0V=�yt�X�s���,�F=	)�<��C=��㼼�<���<e�<$�7=�<�<��g�\9>�c;�<�R��4��;���������<��ٞ�4�+=��%=����Sz���#=�7���gM�W�c<t8��.O=�5W�{F<V� =>a�<	h����>����w��<�
`=a�;�Ba<���<�<	=���<�vJ�!�D=��M=d��+@�4��w5�<+j��O�<UO�<�L=_�w��><z��Y��7��Hނ�ذ�<��=�e�<�dC=t�=Ȕ�<��;	�@=�A�;������μL���/=ld=�>6�k�=C��t�<�rf<ɱP=	ی���־f=�v�<�er<�N!=WSE�*T�<a�=�uL����;�D=�":=k�K�k@~��>�<w~9=O�c�S⇻�L�
�2=��<r
$�5�:�c��=g�T��WW;!��<'[���0b�eN%�x�<8�78�L�b0�<<~=n�ټK`��
P=�D�IC=V�׼A����<��=�A���?�<��p�w���Pȼ�����ܼ�T����<_�J�u�V;�jx�\B�S:=�҄<?�9�_�k���<�#.��Q�<�Ϗ;цp=�O�;��#=�";�??=���v�;�K�+u=���9�6��<[���;k@��m<"<-�+�R�\=Y'���C��f=t��<7��A:=A`�0�=Mq���g����a<�CZ�+���,����;3���� =�񩼹�� ]=�!2���!��5=�'^���9pμ!��mN
=o�I�@�����V=�|8=��&�.-<$���ը%��Z0=G�G���;;����)�u���(
'�o�m�~Q=��\��8a�d�b���߼B-=���<B=��{������x���7<c�(��O���`�����fH=/��:�%=,h���L�QI"���B��<�;
��<y�����N0�T����=�w:[��ce�=l
=��<�	<�Z�f�����3; ��?F����+=�9<����|���.=�Gּ�K8���
=�|�<�|򼅧����w=r�v=�)M<9
��o;=�Z=<x<�#���h��u=�Cs��.=�D�<X�=g��r�<�"�<i���=�:�B=+���-�<=c=�8�<��R=�U<�4]<��ڼ��<�x�<C�.=��缔pO�� =��<`���h��)�<h����B==.���=�J�<����YR<!9=l`���v����ܼ�����h=�8=ޫ�;�41=0�a���"=^�;�����?=�Y�B��4�
=G�h��=Z�=Hh�N�)��<M�g=~T\�%�N�6�<�)���@9���C=��G;7�ѻ�
��Jic�VB�;g�<Y�<����0�<��<4Eμ,=[���a�k�ϼ��;�*O=tA3�#䇼ǱZ�!I�<h����t�����B=�^�>�P�ʭ.=b��<�w������.��آ'=���h�:�C�7��`�;f�8<�]F<(�y~.�w=�����I=<(3��_=�X��u���ϒ;�w1�(=ߵ��;���$;�����<~-=Q�=�@f=;�W��?�<���;qU!=�GͼX�Q:��=����p�4�=:3l��
=�?<>�6=�N�<�EV<'�LQ<�@�>����;�(��{÷��=�| =�R5���;�
)���<'{-�I���d'0=�{R;�=<<e=ܼ�֞��d�<qH���a�Q[Һ��6=��9=0�:� ��L��0o�<pM\<����I	���g���<��[=�f.����v�<��R�/};{'f��(���2=���*��;	M�:m��9��j��eQ<b>���=IF<�]!���;�/=��U�������C<��T=�9,=����T���=��~�_����i����<�̑��k�<읭=n-��c�;|�B�]��<��/�^<D7�;�����=�R�E=�S��\ =�m�^t�<��K=�Pݼ9�<������_��J;=5�<�P=�>5�Đs����c����U��/(=s0����<��亣*��~=-��<���fj����<��K=HL+<��:y:<�\=&`���<R&P=$�μ5�K�va�;y�.;�U���Ը<���<p�m�)}=#��<e5��ӷ<_Y�;ph>�/�<�a��=��ϼ =�w��+�<�	#��<�eB�d6=	V�Y�\�s��<�۞���ۼc�36�;:N=�Tༀ�޼�3�<*vm=E�:<q�޼=�=�<=�<;(�&�� =��L=�tǼ��6���%)=��4=�C>=�H=l�=��y=g�+��N#:Q��>�<�:�<Pws='GD�m� �<�_���-��4=�w~=:Ya�_�<��6�Va=zx|<w+8=�-B�}.���.=���<��E=�\�=���<��=��U:"?=>+�<g�_=�r�<� 9��˻<:����������<��M�����
�K=�T�<g*T�a�Z<8;@=��\��O<ݲ���<`L����"<�K5=ng��V�<=�r�S* =�5�ɠ�<Ç�C=��=m�.�Z�>����.=��;ߗ�<�Z8�����|I�V�:��<���<oyc��Y2�ԅ���-P��7=@%�<@�c=�$	�Tp����<E �'S��yA=aJ=��4�j�<��Z���=z�H< ��)�ݻ�-���ʕ<8W[��c�����V�E�K�s��<7o�;�J�'H�<\�<F0��󻪓�;a�r=��'��4'�/	�<1*μD��9�,=��s�k=���q��<9?=�8�d�;�٧�*;�6=�%'=ή�;��/�
dR=%�����@�~_<��#�p���-�F<�~�<��<"��<4n\�q�=Y:I<���<�}$��a�4o��L�-�����<J*=�Ћ�}�߼��U�����;�,=�.=.�K<2/D�����qE<��K��0�8�<�����:����
��C�;�=<w{�B�g;���N� =,�Ӽ��k���f=ɡ�;͹r�9u%=�B;�럼�� =�� �4�H�dI�+=�Yм�0D� x��sN�E��aX���+�Z�>��-f=�P�;�=#[�<�b0=��z��-/����:�]R<�o�
޼���n=�U<���<	&ܼ�_=�9:�ܘ;$�<���<|e\=*�<=%9!�@�Ҽ-w�|�%����<��<�=�S�;�A,<o��nӼ��7=��b:1<M�<S�߻-@
�v�=�Tu=�Jq=�N2=��*���==A2�VN�<�ƚ=^�����I�p\�lJ���E׼ы�<w] ����D#�ϫ�<���3})��(�93�d��o=G����a����gݙ��=�0;(a��%H=x<F�CD�����om =��u=L=�	v=#˻�D�j�^��<�+8=�`�?P�<F⼙C�4�m�=��<��<�;�Ѳ�<ڿ����B=у0=)�：��;��W�w�h:[����=�e?=�� =Z��<~�;��6�r��<�>�
9 ���=���;h�,<R}=���<�d�<�}i=d��=��?����:o=
�<񛮼�fD=�{ʼY+��P���[�;�"p�1-<�T�@����˙;�6$=s:��Nƶ<8��Ĝ��O��:�x��2Z�� I�d�޼�C�=�P�g��T@�;�ż��j=���<�x�&q�;�4���z=����;�d=b/;���<�+%�)'�<���6����<
�i���O<�@=m/w<�O=@�C��צ<J*���Y�$�)J��8�=�z��]�b�H��6��j�OY=Ф���-=F�r�I�NS=�~a=�n�װ�<�4�xq�<�dҼ����#�<���1<6�ÿ1=�K<%�v= $�5�Ҽ4�G<��:��|�c�X=��ּ������[�(��8Z=�1_:�%5�<i�<v)R�m���E<��C=��I;��x�D�S=��4=�t	;�2�YP�<�H9���<�V=�<�\?Y<n��<�֫��n�<�ܼ3nC��Y1=z]=�\���(!��&�<9�A���)��lλ�s���G=������<R��<	�+=\���G����<�tY;rG)��l	�D��o�S�	O=_�G=:��#۹��m�P�̻����%=�$S�g�=N�'�Hm=��:==�r�R�Z=�e��L��OT����<�-�N��<��<��X�R�U&�cj+=bi'=�%<�e�<B��G=uH�:�����";��@=��{��4"=��}��/S��vܼ�}%=���<4�p=�k-=���Ba�I&�;�u��rR��2G=C� =s&�p+a=�5����;��ż�Z�<+)��LF���<Ȑ�<�ﴼ�4ͼG�ڼ�м�L:4�p��ll�2
�<i/=Oh=�p�� 8=�0ȼ������`=j!�4�A�W�n�<��::}���/�.;%�&=�W8=�`���<��1�0H0��)7=̋�<[ĸ����<M7������ۼ7?j=��N� n7=݂�<�^�<���<�|=}�<f	 �*~=P�<�S�т^��D�'A�P�6<��d�;�9=u6=π�<Jt�<�J=�=�|J=�̘�@���~ f=`���Saf�nZ�M�<%�v�[�ż­�<3�,��.c��bؼ�/���i<��,�f�5;|�]�5q�����/���%��t���=��=���\�;6=j<k2�o�+�D�$��� �=���"����qxٻ�S=G\=<�������@��[��A*<u�;Tϣ�t��|F���=�����S=i�"=`=�<�Y[�� �=��ؼ7 ü��e�� �;�����<�x;�S=��P<S::<�jżZ���U�k��v��"��:CcF�C��<�څ=�J�<-��I�=�M�/�L������r���d��;+�9C?=0C9=}T9=��Q=GGR=ѽK�����*�>z�=ѓ�;���Z�5=x)=��$��b(<��
�������<��]��vF��4X���.-=����6+��A���y�<Ꜽ����ˤG=by�;��ޓ<\r8��\�<EŴ<�Y=��:�Cn��<F�q ��@=�<2Kj=th=FlY=k�=��y<7j=$�)=ẑ�6/=+7>=o5k���K=s�=g	����<1�	��Ig=�/=#�L<bM�9X�<-9ѱ:�[�:Nep<p�=Wq���{<:G�3xl��=��-�4J=����=�}�lh�?�<�%�<�O�<H�p�Ac�<c�?=ܼ��
~^��}���0n�=��<e�H�J~Z��S���<��<�
�� �ީ1=��<�؃��YV�" �<��F��x|��� ���5=��Ż1\i���3���Իt,*=���<�&�<'A=�+��hȀ���(<�u �/��<���<c�X<|ͼ�7=�<tJ��q�p��i}=zE�<	�<�J�<<=���c	<�l�<�_6<��D=|��=�'��:!�.Ѓ<�2�1�+:=�8~�)�Z�YN�;~칼�z;��T<�$^�� ��H�;���V�伩	��
��<;��<�w=.���ڰ��Qw�<E�(< �ǼAї�Yx<A{A��3�;�������$���vR=�]V<@�<<v=˩�<�Lm����<��<Uy[� � �ܜ�>��<��O��b=��&�ICY=�i����,==l#��D0<�p����*<Ļȼ�yV�AK3��$\=�6�<i�;�M:={��<}f�;�q�<�ռ$=�������0��]�Y=�(�3�=���<ݬ¼�SJ�DXE��=�K�<��(�m�D��K�=!��<�]�<��:="�x;�@><}K%�J�n<�e=:%�X�λ(������<"`ܼ�5=��,<�?��FF�࣒=^���p�<��0��_d<�$���É���IwM��N*�$�=爻�9=�<W��=�KW=��Z=r���ސ;�Ի��~����;u��W�=��-<{E�@���8�C=�'�#�:���A@@=|Nܻ�����F<�ټ�3�o�<�ޫ�/���<���<F?;�ʼ��)=,�y���;I9�@���b=�[=l�ɼ�j;l�ּ�Dϼ|�ټF8�;s�S� ۼ9n�=|�<*G��������3=S=d={�<4n1=�`�<_�e���r=;\=���=V#`��y�b-�X}�<��o)';�4���U.<�E=���<`�D������1=/�߻5ia=���o0���N;+Vۼٮ"��E�<j:S=5W]��W�(-�7�
<���<<�ۼNp7�H���<��;>dG��PZ=0=¦R�5�Z��0E<�6�<���g*�bt1;��ȼ�/ٻ������H<��/=4!�F-P=:/޻ A���
=e;�g�i;DO�:S��<�z��f��S(=G���=�G=`�D=��_=���<7�,=��A�N;�<NK=�u=��m�=|�<��=9�3��	<72n��jy�=���<�<���<�L�;�}<�ȅ<�|��`ǻWڼ�hz=��;m��{�F�J=v�b<)~�Q;��:=]�?������<o� =ؓR=I�g��u<j�;�ȍ�g�c=ZC=�U.��%�u�g�&��b7�9�)���;O�-�HP �	��<���<]F�<��w�׷���_J=�q^�k#|�&�Y�n����5ƕ��j��� =?=��
=��>�y���=c�<9ɻށ�<�<=b��<��T��S�Z�䦐<�2z�Ve3��zX�ٌ<a����Ee:;��SŶ���<�ʁ<��d�lpb;Q��FQ$<�
=�b,=+�<�����L=&��=nqE�h�0���d&=������<��2=-G.=�%o�r�a��J��J �&�:�==J�1�p�ﻌ�<x�����d<9yt=�=V=OỐ�E=�sn��eM��ˑ�ú[���=���)�=LbX��A���D<������<��b�&=��~��<���;^CQ<DS_=y"!�UQ�<(27=��<HU�Ѐ=�FL�p{ͼ�J
�"s<��\M<�""�5AJ;E�=W�<a,�;�H�皱<��F�X.c�=�'=ΤL���<6_>�hEC�+=f�8<0�e=���<���:! ɼ�:=��<hG=0L���=/R�<�Q=�^�<�c�<��h�q��<Ѫ�=B�T=��ػ�,1=c�&=��=�$=�	�;p��<_m�;��|��?=��;e��<E��=<0)������
��ߪ�lRX<%�Ǽ�|�<4=��h��w�T=�1=͗T=K[=��<l�z<[�z=���L*˼���<�<��*�X�:��\=ʖ=L���n =�.�<6G;YP��'�O9��T<�ź�c�<���;=U�ɼY��ʺ#= X=Qlg=���<� �ȴL=��=P��;L=f�L"�<S��<�K1=��2<�yx;��<�E�T�S�M���<"9N��N�<��ϼb<S=ˣ�1`=�r��;Y�c�	<`k������(_=Ra
�{d=�cb<��/��f�<���C��7|���<�1�� 6�4��=�Z�j,ϼ�~[<{E��f������i��L�L<��>=Lǵ���<6��	3�Mr�<�<r=�;780��{�<]�ټ�
�E�~�	Z���NT=�h��֚<�P<�-����=r =�IC����5#�b:�8Z���k��2�?-���}x=<=H�"ρ���=��=�u1=�)���+�R�=�1<rt����(=0��<��<��<#[G=�Ӽ�5�
�e<�̻��<-�/��,0���U��n���kO=�3���2=�?�<<rd=v��<��<LA'��3n��}W�p�*��̼�o�J�< �k�\�=l�*�1@�;�Cb���3��C<��<����l=��$�G��D0=|�4�(��;΀�;+�ڼW��<X ����e���E=�����P1=��=��k�z_7�Qc<����f���<>ڼ��6˼v�t�#��� MJ�'|�B��<}�4=�/��a\�<ρv�"�0=������!�=0D<�Y=�
==kļ(*�;�	<��Y=����Er; �za+=�=-n�<0�=��ܼ!:;�D���,�`���[��t�t?��Oq�6��g=~r伃gY9���<,����X:���`="��n��t=/�>=R=�<��hoY���;F�<�f<��<�=t��<�s��'==�l=�4��|�<E'��7P6��*���<d������rG�|��<�~�84�}E��s7<�D6=�+,��Q�<jش<�̽��YE=V�
=/���x�9�=M�<��;<:��X�E>���ռ�fS�n�<��<;Ub�<�-��yO�:�9=_/��8y�H����0(=�T�����;T����s¼�B���;�ږ<����[���Q�_ݺ>Ie�Pġ:&>�xB*�E=��A��eD��=��<&�k��޹<��F���ZQs=��=�@=�ϻ}ƼM�=`JI=L"=��N�W�O�]M	="޻��<K��ڊc�v�=��0<��X(X�����I\Q;q�m=��T0j<���I]H��j�<��I<��<�=��=
E?=B#�;sV=� >���	<���
IɼJe�5�=��E���;H7��߼�(l<CM�<�*��
=��*�=�� �;�Bo��F
�+c�<�_V�,� =�qG=e45=>��;��=&r:�
r��^��<�T�<��;���E8t�+���M�=b�8=LN3=ގ0=ǯ����h�;=d_�=�+�<~A;=Xc���M;]�ܻ+t.���~<?K='��n��b;�%��@~���l�<[�!�A,=�8g�Z����(y:��=d�k=�<\$=R�;��;�!�<��Kh�<P�C=n�d��U���<�x=aKR=	)#�����H�=}�@�2�=? "��7��xԼ|�=�1w<��<�,W���+���=�t��(=��h���B=K�N��~*=�0g=�W����<Də=y���4p���+4=7�*�D�f���	�8�׼�h<�8�=~�E=>V���+���e��#�;�� ���@=�UF�~7O��$�˷��®;ӡ�� �=Qy=�+�<�6��֠<��=��=�o��@5�<�vK��mJ������߻����V�{���Qy�<0�I=�g\<H7Y���}�6r";v�j�ɍD=SF;m+;�W<V�<v���h���\=�V�<��0���7=ާ�;lq��*s\���5��\=ri\�ğ�4#;�,&<�� ��u�<Z����N���=���<�� ���%=�VK<��*=�h=v�ӼĹ8�Fa���<Y-��<��=�V���i��N����+/L�	�+��
��Q,=�ל�E��<L#a��Ni=D���n=�[�<��ü�7]=%�(��V����.��;�����<y�<`8{����Ik<���\<~�8���輧��<��</T<����܊=A=��<���Y��<�	��T�<��лɋ �/�=� =�?��gd<��M=� V��N8���r=:6x��-ڼ���T�$=�c<W�@���[=�|�~�׼W��<|�|��Ӑ��#�4	�<��B=�Ѽ�/?<E!N<�k;��
=~���׼w��;�ۚ���<�9����:�<�9��= =�r,=��<~2<;���<�@¼0td=k�Y��l=��<X�$�}�!����q2=�IܻjRB��
�u�M=&H�V=���<a=b�qn�=��&���~��o������;�z,�ǫ���G<є���Cݼ<�ع܊м�bF=�{v�t�J���׺W�Z=�>��Q���M _=[�=B���2S<�T�=�SL=�6'=Ѻӻ%g7=$s=��D�n�����$�d^�<`�<�L���<KF�t�&�{+�<e�\=;^<�I����<C<&=~8=��?=�T��=fǧ�x�<7��<(s};Ԩ=ҲѼ�������@��IPڼ�<B=d�j=,T=��r��O/������=���;��ܼ��;ǯ亻ZT�B�<�� =+�;@�Y��{��NR���a=
,��&/��=�~}���q�|�#<��1<J�L=Z�[߃�`�Y���z�����ټ������q<>6(�ќ���+=Q��<�K��ҏc�iB=%H+�l����B��� =ۿ
=|�=&��<�A=�V�;��Ӽ�e�<^B�`�׼!��;Bd=�8���E;|�<K�P}8=�<�<�k<�U=Vٻ�l��lk<7d��,�G<�ɒ���k��μeM�`a}=�D��=�3�<E��*
��'R;i���<=�@�<V=i<���ރk=m.�����b5�<�	=?e�ٚJ= �<=Oo�<$?Y���<Pf=*o,���g<�H������R�<F*Ƽ����2N���6����<��4�|���%�`�<#t�<�=�W�<���<��e��� ��D�<���;xA���(�� E< /��J$��=�=6���:�A�v%m<�E �uD=�SмPt�3n<L<o&s=OG6�m]�<�4�;�i=�O��"d;�S�<��N���,�.�����M=y��<�!��Ɂ<��;�$ӼO�=�QF=� ��c0=$b<'�n=[�$��z'�#ȼ/��`Ay��s%����^�����U��Q��<gH�
U��r�<h��<O)��-=�Z�C`���<���2;_];>Gn=�d+��ŀ�/t����s=h���7&ּ(�9�����8�r����<%[�I�%����<|޼�DE<
�|�i˻�ŎH=-�v<�� �)*��~�>��d=���Qq��ܒw��ͼ'�J=�c=/2r�
��<�+��&�U<�ە��UT�}	6=��Fg�<�b�:�F< ��IC����_��D����:|��f��BD�����1ZC=v�<BIX�.��#��y���rg<��U=��S=�DU=��&=;O���<�X[���
=޲��$4��*=Ã��$�B=ڐ=L}c�����x�=1�=�u ��ew<�t<?Y<{��O=�x(=Q+�<�_m<�$S�Mё<r�Լ��˼��=�B`==Ug��	=��=�=�r����@����<*,��B�=1���c�I;p�=��Q��s=���7��8��Iƻ�N��p�мNj;�y�+�;�
<��W"����rY�~B=Q{<�B�<Q~ɹ��<�}�;=�<?�`��劼'�<���{�;-w.��S�<�l=�D�<�pɼ7I�;����*�����>=����.���=;��Z��T��<3~�<�;4nM�M;��������,<�q����ɼC74<��=�y)�aH� W=����""���<���-=8�d`������l�����;q�=��׼y�x;횐;x�,�vUt=ϳ��=��<@��<�W[=���ae�<�M�C���� !=�B���eg���CF=U���M�<5�;sy����
=N�@=!I���<�5=�F0=#�_=b)Z��l=�YҼ�|{(<S�x=��?�4m$����<����1桻���<= 	��Ʊ<\%�<��=k�I=9�ż���n��B]=	�"=����<��#=�(S���=d=.�w�<H�:�i�<�0�Z���#W�:0=;�Y=���#&�M7���ߕ<��.=楜����<�J���c=�A �'��<`
7�k';��㼡&-���A��b9=b�����:&�����~7=�ɉ;:u�<�wO�o�1��Zi=�L������tN��!G=Q�];�ê��͊<�=�4O���	ɼ�1Y�A����<SZG�|}�:��<vJ<6�T=T�<�/��=�-7�~�<8��'�4;�j�o��<��<92�;�7+=�?S�f������|�X=�� �#DJ��r&<��^���~�P-=�]J<i�=�>�<��&�l&���Ӧ;V>1�s�/�,gH=��"���j.��r=��H�8u�Qv�	u�:�M:�{	ٻ��H�f�f���_�� �XZW=X8�l]/��sO�d���i=hE��~˞<�F=!���r =��"�U?=z�=�(=��{�R��<D3�w��;r�<�?�<3'[=-��=`�=���Φ=�hx:e�V�_�:��#=z_�|#=X�=�L =j���ǵ��}<qS3=��<�><�sX<-#����<D��:W�<h�}=)�ռO2b=�W$<<j�l_b<�3�+sT��y�c��A͗<�2�=]K=t	��-"��&�ĸ��e=#���(����^���<�=j��)��<ȁ<��:;�Z�<>�ؼyҠ��/=e�����4=�</��2�vl�ؾ�<ו8=s2';�4=��1=%==Q��
'+���'�LNG�T���Lm=��|�:�S�!�t�LSN��-I=��,=1�2=>�C���z<�$(�����ERT=�)<
�_�g�-����;/S%�̐;�=�^�;g�̼0�H�#�>�֬�
���x�Y�׼<Rɧ�^�'�~�ֻP�-��a�� #�u�?=д;��n��!i�KT�l�^<2
V���#=T�=��J�
z]���`��9�ʯ<�w�c*�ĹH<�8����<�b=�I��`��D�c=̤<�x�	=�V���J=z? =�ܝ;�GI=3D�6ž<�rۼ�=����w+��Jm��d!=M�<��U:-���~=
�<C�B�>=���<W%Ż:&�<c�=�о<b=���<y�<>�<@rK=_M;�(<ϊ<SW��:#"���K=
�=`���?�<�����e=}:K=z�\=�*=Cn�<�R.�F3=�1j��Y���Bȼ�K�<R٦��X0�k��O˒<�T"�_�!�
�=(�T��B#��� (���~�2���A�<�Z����H�=
A�г�9>���غ��b=������=vC!���Z�����f�8�=_ȫ<G��������T(<5�/=��輭��L�<&k��j=��z�F�vs�E�C��d���V���	���<r�Z���껒 =k]=B|�;W�k=ұv�!b	=r =�G���<������P=�Ӌ<�
���`�{#=\�'<�7�lZ�;w�;ގϼ��Q�^�<�h��H�G=��j=�<
�2;=����\���|<�"R���P�ԓ=��C=Y���<���v<z���TE=\SE�ά�(��<���=�&�<���"4��:�1�7���_<��K���w=���<�o���c.=�9=�Y�<�!��<==���;U��<ק$�)Ʌ����<��Z�V5ȼ�7���i��e=�Ś��$U��EI==�"��d�[w=�u༎���,�<��H�v�:"�7=��Of�;"��=/{o������=�Ș���<�l���.���"�&c*=�=#=�J�uO=�|O��6��? �7�<b�<0�<�@��E��=�6�m��<t�t�m���j|I=��6a(=bڼb;Z=�w��)O�.��x��|��<�;��3�[��<8iѻ�1�<�6=�:%<^Tl:�X=�C=AS=�x���q.<l�V<�����;�J=�d&<e(M=?���a�)=I�"��!���<�Zл�＞yӻ��̻[�!=B ���}k�9�bM�������~�߼�1��.W==\x��T༩�.=
�<��:�X<�v�<�<�O�a;l���m�2������<k�~��8Mg=I��y�	�ۜt����<]
�<���</�Ӽ����'�ɻ$��;a߅<����q
�_�Y<��G����D��O�<�Y�X��<'��a��<.>F=�t���<=E�����zԻ�[	���<�<�9��Q�i�r���!��Q<lHc����<m��<��P�<J���=:�[=�W��)��ʼ�P^=���Q'9<"gѼU�E=�[�#Kt�J�V��>���"����	x=?�3�Y��<��<S���FI,��	�����;~F�<��N�Jq�k��hU <��k�<�����0��Ū�����u�<����ͼ��<е-=}(�<�-f�.���Ԋ:%�?=��C=0ؒ<fC�<1&<�=u5�<)��<��X�F0=�/��Ȉ� eK=�<=�;�o@=�{ּ"�g�$4*=x;�=$s�ڭ9�w�M��6q<Z8�;�m��
М<�ǃ�s��;3+<�p�<�lf=�v׼��ļ��=BF=GO�<�H=xü��<F�ܼs���%�p�t��0��<^G߼e�����/yP=�4�=�`s�Q@�g���r<��G=6�<M@�<7�h=��@�
���J=���<"W�;T��:|��;�����W�G��lC���B=�D>���I=���m�~��;���xO�w@w=P"m���=�Ah<Ӡv�@t:���J�vI6=��</S��(��jV�����e��q�|q=�ׂ<��!���V9a�<���I'<�8l=�0��\T=��<��s�݂b����5�@<��}�E��<����OH< ���-��;;'���0t�ġ:x,�&<�<�yA�*���R=I0�;֋6=��#��<�>�<{N���Z�;K��<������M=�3ۼ�±������<|�e�����_]�/�=���<F@8=COv��	���&=�<8B�IJo�(��T�[<L�J=3��<�DP�oߏ=�O6����=�<��d;ґ�⚍=��;J�=�.6�4� = �b�O<��a�A!"=�P�r���\��<�ӿ�K,E�S����Y�.sX�tf:1�ǻ��:OW4<zA���T<�h(=�;><�z7=n����z�?��=]J�;����gP=�a=�㣻`�����<��a=u�Q<��)�����ּ�<���^=���k��z�<en���;��;=	E���{���mL=�U��};/�zs��A�<:B����=w"�:R_�<3��IS���=h��|9x=6�˫��=����T�4=��a<=��F<�� ��~�<��=/*�<�J�j��s�6�я�<�%<4G�<WQ���2��|�7�V�� �V\J=M�<=̻Ƽ�ڦ���O���	ȼ�!���O=�H��Ҁ�ϛ�<�Dj���P=\��<H�h=�=3�$������<��a<�$�S���F=��)��়��&�s[K�ª�.�� b�=
(;@����U=8:ػ���y�;m�S=�F��݊��l�������kL�3����N�<>�<1N
=��,=R��=�)]�}�4��x��g<�3�;Ft�<�)�ͺ�j�=!�ټ�'=$���6輸��<��<͐ �Xtf<\
=iy��H��<�e����;I��
��b
��!��%7�S��<�O:�hI=�*���=�M� �ĸ��*=��p=����1Y5=h�O�,��:����3�;Y�9�4�<|;=cRK���<HoZ<W���=�Ƌ<*�<Z�D<T�:���=�:�=�;2).�$�7�][=+]��d=�!��\ѵ<���S�;�FHW�c#�<?aH��&H=n�#���=ܕ�<a���ڛ<&�=<4 �k�=A�5�.f=kz�;�R�<�e���=?t0��X(����<������<ԣ���,�#��<���<\y<��l=�1ٻ@�=�֪�9U�=�-=���N�J�"�I;��b��廹�B�k�=Mv��O�F�f=�\��Ӽ�
}:ō_=�"�=�M����Z=E��qv����$�
=���;Tp<H�7�E�0=��	=^��´�<܎5�'�=����M����<��9=�`�a�/�U�O;P�?=n�<,3��:='м�#=�9��CWD=�m=?�y=�s�)��<[��UĻY�ؼ&�Q<�0���N==��
=/�:#��<�ͪ��;����<�J;*4��l��P���':Nq�?o[�����y�<��1<��<�O =����b=��$=�ѼQ��;}�2=a��ѻF�K��:]�<�u�&֎=M��<�_6=ե0<~$n��Z�R�2=�?�;��=���N����<p�	=����}N�A���^��g,{��(+�O�D�:���Ż�_�<>�m�H�
<{==���; �2���:֑<�B�<�cd=��=Z�C=o�̼��T��]<V�鼜<A��A7��c��R�<�<샠<}�F�{`���=�9=�R���s=���
U=�)<��M=����Hg�(�ļ��=�4�<�v�y�M=�T�Um<�
����O��Su=�<<w�=�
�����%=uzx=8���лμt�<�S���C=��=p�Ҽ=Tn�5�R�_H����<-��;����2�=��~�<��=K�<����Z��<$v�;��a���1�+�¼��M��b=N�'�����0��<
�=k&��8ػ�[V�h?=��S</
=t켈7Ż�:<�Z�<�y�=�iS��DJ��N�9�ZE=���������H�;��{=�E<�<�b9����������a=@H:=�����W��g_;2/=��V��)k=˻��E=�*6��]^=�s���#;��_<ݏ/��{�	M�<+=�-���/�%A��bL;]�/�jd��RK��'�<B
����軝;ü�=��*��]<^�<��̃=�_�=;#x��J=	�Y=3�Q<#��$+ԼS	S=Da����<�d5�H���邼�}?=[F�;��;L�M� �U=ك�<�2���a=,8�;����<�!�(J=r�=$c<�@=R�!=�޼���h���u=�VX�6�H=m�+=���<Z5�<���<���;��<�� <�i0�~�$�ǉ<{KW�ƶܼDlO��0��V.=�����,������<�z�<�k,��jh=��)=T-׼O���kI<k��3������<���J�����;ʬ���dI��A=��x<�5�.T�<q2<\����]==/��f�w�ӹ�;}-=���<�
k=GS�<Y���c�<����vS<%Q!=��q;i��R!��0W<V����*�'6��kZ��'�C=�6=�=�u�<�G0��� ��m:�������;!&ɼ3�=�䀼�Y]��o����b=�G<��|<*��u�S=B�]=Cwo�l㕻LbS�<�<���;�B=u�[�X��j0��C9;J��<l-F<Ջ<�L���+��"=�-�;Ds�aaX��W(�W��� <"�A�W�e���"�G��<H=� {=d,�~%ü7����#=}л�����ax=��;=��(X��Zɼ:Y�<��@=���<�0��� �-3h;b�߻-/Z�$#��S�o�`<�|���a<��=b��j� ��i4�q��<0h!�go�s�#���^�p
8<���;,@=���F�w=K1�#�ۻI�ǻ.�K=�7#��)=/U;b|I=�é�~*"=
��� x�<�Tc�`*�<ѭO=TB��w�;In�<�Ԝ<RỺYM=RA=�l���Z�G��<S<�;��9<�};Gʻ�RAy���=.���%�c=������<^�f�x�O=�xY�"��3xo������(6=�|=�D�a�3��m�<��s=�	�Ƿ���=�ME�5��{�=1�0=ô)��Ɲ;�G�<�l�;I�C�zl���2��'��=%0׼�ː<��<(=8ꔼ���k�N���O=&縼��f=���;��p��`��5=�>߻݁<=������k���!=;��z�"���y<�'-=MH�qD�=��oS;�(��;�}�;q�<�4��8��Z8o<x�<,�Q=������B�7)�<� �\1=���B�<z���=6ep=���<���0e5<�b�<i��F�;�Ql�~�B<Sx����<Q�<y�M=����˼�V�i*I���?�px=�C���7���t<�3��GW<?�=��<���"�̹<.�>=f�4�ꝅ9��[=���� {���Q�Yص�^$�<�QA����<��2<�-��i<�w��'��<7�e��c�<���<�~��b�<�����Xn�(�=0��q�O�
4&=|輗�/�\c��ۜ����i��Z�5�phW�1�#�u�r�G"��7�(��
�=MA�;�<��=m�<�ц�9Qg<B�<���߉C�46���=?���=>�O��$<s����0��?�>�k�E;W"=���;0��<\Ϙ<�h=|��n�< K;�u��ꥼ?A<8T=�J�<@�=o���<�ʀ;��y=��S<Ph�՗�<�V#=־���t<d|�<+�=�/=��;@ �ۗ;=i~�<[DY<�-n�t��<6)�t㼙\=u��<8?��1�=�V&=S�*=�.��@��;v�<�Lܼ�3+=I/f<gے�x	�<�	5=��d<�=��|<�L< �X��.��7'�H�]<��<�	��$U<�nF=`�=]���ƻ�$ϼ���<1x�<3��{��Wռ2����Ψ<J���?4=�T@<F�:����q�T
�<�Y<��I�<�<���<<�<�y��(ٽ<�>=��=?O={�x<@H�������$�h�μ�H�<c��%�<��������g=���;�~�;yf��P=f 6==����6<ݙ<����,�;�J=��]���C��������;�Z=(=�Ym=�D<�T���	���=�gx�E�4�k���>�#���:���o<�v�s6�<�r�����Qk=�1>�4=��;�i�<8	��i1�+9J��0=��Q=e�=���:�F��+����ڹ.y�9L�h;C�2�n;��s=��-=�(��7=���<$�n=��9��el�>q�;�$��E�:�ﵻ���<d��<j��s�
=ŷ<ۯR�^�9=" �<-������M�p�^\=f ��K/���=�LX���˼���fL��;=�E@��ֻ��r����<HH'�Gһ�ݦ<�6:L5���=��=F�M��8�}��<�(.=eG����~e�q�e��%V��{����u��Es<�� =��9��\�K.x=��ɼZ�y��]u�=eN��s=b}�������Ἐ�_���N�w&���>���=�ʁ=�x���9;/�J��5�������%ڼ�f�KV�+�<TM�����;ޱ=;��ث�<�Wp�@���$7���/<}�(���S<���<M�=n�n��%�<y�����O�<�3=��;^L�<� &=�a�;�＿��.@#<M}F=z85�@���ټ����V�9�I��<F�M=�W�<kT=���l59�Z~G��-��!��XGJ=IT4� #���,=��%=��T�[m�:o�<��żlf���><������B=d��<��ּY�����;v肼�PI= S����ӻ.�=;�����μ+h<��<�W���;.H<v�-��&�oD\���/=��Z�<�Pv;j#6=Vh<�um�dϱ:xH;=�J"=����/���A�=��<��f�uv¼;<��<�V��CѼ��j���|���O����<�3+=������S��E���Nt:���WƠ���;`u�<0�i=�Y=��\�E�q�O�B=�`�[�M���=� K�<������<�"Y�T�Z���4���1=TP޼E���"[�=k"=������׃<j����
������d��/8�EI=,_:�A�=�'ݼ�t=z�w��+�=K������pa�/a�<6�B�lvM<���<_��;9A����?=_QQ���C<TQJ=m-���M=K|:�z>=�^ =�WD:��%<ξ)����<�5�<�ӕ�GT�t���?06��~��܍�?���*�G>#<�6:��h5���0=cL����oR��"���R=�M<ʗ�;ޛ�<UǑ<&�Ǽ�j��J5���=E����d=~�c=C�<ܿ�<2�<���izv��a��qmF=��g=��p���=��?=4k��(P=N�V�nxg�׋�< ��|fm���=��K��f=���<|䖻�D��zO<��<B�<6��1*<������!���<Y]�BA�<Q-����;z��������.���s<���K��<e�0=�%�=�<��<l�L��#=	� <�I�=>,�è=� K<i�M=[~=�Y��\+�j�z=2�!��dY=�GK�V7=�ҟ<l��kB� �ϼ��-��	L=��8=!d=�ݼ1���%�\	=�	��,��Q:��;d0=��m��H=�P�<�Ml�]��<�I=S�m�=�:�KH���~`
<��R='S����5����==�S�� ���H=*_ܼ�#I:Mg&����<�ż�G��:D<��t:�m	�b�9=��N=݉�<W8n<X�;=�{�;fX=~9�Ŧ
=��I��un=�6r�n�<"'��
}<m�	�ǐB���>X���P����,<CX��O�=$/2=m��<ws�<& j;hI����=F=e��v�;<6�6��e�p�<��;�FL;��ź�HE=j�����<郩�j�-���=�@�(:ּ�ys=/��<별�+<\��;^��<dT =LØ���(�zkl���8<J5y��`�<����DCԼ��<x��5$N���=8j��T�=�P-���Ѽܽ�;1��q���)p���)[==�>=	��</��<u�<l�A���50f=-=�Z=��߼��
���=J咼)�]<F�<�	�Ĥ�<��c=�7(=?>�<�4>��x<DN;��<=$*M==0�<suL�~�V=�w^�G���_?�M�r���_�-�<����_tἶ?L�2N8���c=��_=h\<e��	��<�	-= ����<�>�<�O<pr�����Eqʼ3=���u=��>;v���X=������<������c��*ɼ=�r�?����;�q�+̻�˾��H�q�k���W�;��<�%*<��!��ּ��m<Q_�`��n���`ܼ�3� ���?=�Il<^Ԭ�c�ǻ�IE=�EH�<���V��9��<�!k=`�-=[���,��$�d�>=�<zj��)/=L�&�K�]=B��<�Uo<�A�'�<1�<^u�uw2=���9@-<��</_�<<$�<���;M��<]�׺��m)��?��60�6��=��/<��B���P�����Q%���"��F�<���<p�=�If=Y�;��g=VM��v7=Y�0<�e_=� ��`5=T�˼qH����=W1�<��h=g0��D9=�˘;�g�<&=�����<��4�_;9=ďG<Z�<��O��[���J}���<7�n<0_^=� �K�x��'&��=I�=���;��#�s�=JC8�x⤼ق��Wʼ�f==yH�<OL�=�!:�샯��P?=H?����x=&'�1)˺��A���V����<H�<@�;$�������������Ƽg��`�=F�����x�\=9,�<�2z=�Һo�W���W<=Lf�<%;ɱ��T|�
5Z=�_�<��a�)1�p+<��=���<���<i���?U;�X��?�<9�@�Jv:�bG�(M��==5۟��[=�(�b'�)<�G#=���<f�U<_�=�ِ�*��9!�1��H�u�u�<�4=��0����b��8�)=7���9û�Ye��ݚ<��=��:@��m����]���F�i<�?���h:���<L���IN��U'=嵺;���<f�U<[zH=$Ұ���%=�ͦ;$�i:\�=Z��0/E��S<wܠ�G�=���<�;���=w���;�#=� �N�O�b*p=��=�%�����ʋ�-	=\q�.����<q�0��Q�:W���i�;8�v= �=�ƻ�T�`�$�	;M=Ph�;J�+�o�<���vۧ���r�%�6��b��U�;D[.��Y��a={(ؼ�8ļ	Q���>�

=��<L��<e�<G�=�g������m6=U�=-�$��S;�(=�.=�ų��`#��غ�~<J�/��O:���<rY<]��=An�=�ߺ<h䡼_��=u��<L Ҽ��＆xy��B��2���U�K�Jׂ<�ߤ�b� <2Y<!�6=0�g���?�O�<ԋ�<��s:J���;���^�����r��0���B��x#=I�<�`G��Ֆ���i�;0�*=�7=:'󼔔�����-���#0;�&=ꗽcf=Y�u�ay�<�'5=��=gAH�XF�<�.Q97���Bk�;�]�=��[<�Ṽȏ <D��<T�Qp@�4k��Z
���wwټq9=���<׾4;~�9zQ�>��/�R=X\�=��S`��ڼ�"<�wE�<�UA=��p�k�<�|�<�UI=<u#��!���ZW�Ϲ'�����i=Jh@� �:�ޖj��8<��l ����<�<=k:`��g<�O�@�&=e&�#*��;�8O=�v(�;�+=gT=�^o���,=��S==���%=\-=/ƻ�J =%��<c�Z=𞅽��e=b�'=0����<=$<<�"�����<��n���_�;�Fe<�|��!˼P�Z�����1���FO�<=��<�Ђ;��ܼ3��:�J�ּ�Լ �<�:H�m=ZPB�µB=hm=�u��W�;�X=�=�Q;=���<I�̼�g�����Os2�dD<I�B=��Q��K4=E�=��<?�m�����:=$���{1=������?=�J(=�<Y�����<���=ӷ�=��:]FL�y��;��=�Y=��=Q�;��T���;���6�_m���);��6Y9<Y��<�C��?�U�@<^�<�����<5_>=�`�<_�a=�p���Y��AD=LE�<M@<���<���=UPp���򼅰#���3�[R5�e� =dM���<{3'=T޹<S�r=@����c�<y"�<��o��9=<�E=�J�<��<��L�������<\+e�I�ӻ����D�?=��;<)Q�����&P�~�׼׃㼹�=���zD<!�A=jq�)�=��W�m���Լd~�<D���O��;ף��K=U�J=W��+'m<��s�po���Ƽ��^=�L�;t�<}<=ɥ)��a+��cB�$ټ����T�<�p�;��B�0j<=�3<b�� ��*�є��s��<��=h*l�W�<�u)=�[�;�#�<�O�<�nּ�I;`eԼ?��:��t0=\�����̼�Pq���x�aJ4���=S�?�U9�(�.=�\%�=�E!���=?Z�:�(�^�����<�>�m��k���u�<`�M=K�=�<;#�=�)׼�ԣ��`#=39=>�̼t��m>�<��`�sC�<@Nݼy�=����g�<�]!�<��J�'=�m==��*=�?=�4h��K4<F���[<%��v#�T(�<�:3=��&<�=>-�<�?�=���9�b3<)W�;�P�<8�]���<�
Ẑ7���=Pێ��ƼH� ���n��C׼�8�<�� ����A= M=��P=tH&�l9c�|?=�B=y�=�(�:�$�<c�<=�㣺Y� =c ɼ��v=��r��Yl=XV����=��WH
=�ݻ<�Ou�T[\��Z����<Wh=�6�X�N=�d�=R�4�������iP[=�1<mr?�\Q(�
T��ds=�"����9=W�<�c<p�U��|��'�OR2<�z;�
[���=�b��_>����5=��m���!��ѿ<��^=�=<��b�k�d�F�(���༄�;_�<�ļ��E��-���?�i)u���Q=�O2;��B��l��d�<;=_�=�������	C�>��<�&��9k=��<��( �.[�M�
=�e|����;��+��M;�!�E=�`=�rB=0�L=�c=����P��~q��=�&����e=,�3=]��; �,��(�;��"=��<�J=S-�i##=��;=�bR����;ݦ�<?m=mw,�ԙ���м�C�;��ӻn����Nn=���<~� �'�\=�rݹ��Q�%��<J�0=���;ݟ �$T<B��T�@<%~z��:�=&Y=^�=����
;��<P�H<���_"ٻV��<.a��N�<��T���W<����<9 $������?<�;�<̦�h����w<�iR���A�+m	���Z=OT���~=�W�<a»��8=��-=�q�G34=𘎻�]�;��3<uʻ滑����<1_��` = 
-�?�X���3=c�&=��E���������<�-=�k�<D0�?C��i|k�۩_���<�I�;���<c��e����K�<;Ʌ�� =�n\��t���2=�߶��`�:U=����&�<�R�Ծ>�P��zH/�eu߼)�A=��l=5M=5�.����<'K
�i�o=/�x��SG<��<V�_<鲿<ϭ�;�+���%e��*��u<6SI<8`�:��%���< O=���<&<�w�+n={}�Fo<�==�K<�_�����<�W=�J����<.�*M�<�����O��:=�Q�<pZ8��c�;��I�7�Yq����m<�g%=��=8F��ѹ2=�G=����˼��9[�c�G=�Mt=�P�<�k�=�ur��CU<���;��i��e��t��"7~�]H =�O�{����|���2<��<��(=�Df��z<h�<�<|52=���;>�8:��<�]�����Yw�<;fq�jJ�p�(���L�7̻��<�ؤ�VI��=.���p���D=4Z<&i����T=T=����I�2��;3I=�,�����G=4��<�W4=7d�<ؒ>�Y�R���Fk��1y>=��3="l<Q��<ts��H�u��Z*�;jx=��<��2<Y�G�=��Ђ�L��;� ����i�5uE=�\�<�W�<"9��;8=ZI/=�<��t!���=��c�d�#<V(=m�����=�t����=v�<��)=.�=E��<�[R=e����<��� H=(�g�.c=Ŧ'=F=��;�P0\�-u�<�%�;��=mQ���s�%�L�p���:�"��ɜ���h=��A=�f=��j���A��I�p�;��k;��=��0��U=+�?���B<�	|=J��<��=<�M:�����N�A?<�#M=���;}!�<��V�v�X=�9=��M��_{�p�$=�

<mu*�}�����=j_��d�$�%�=N45<�=5��E��\��";8���A)�<�1h=�9=��
=���8�A�~u`=��֞
����G4;=��=n�I=�>c=�V�<�:�|����p!�<�W=���;$�n��c뼾su=&6=���������ߝ����<U�'�Cx�;�z=ءc����]*=F��<��x鎽�%���\=�;=���:���<�4I=d}}<X{�B]*�d�d=��:�5=n�=��R<@ =��;]7-��c<��E=	�< ~�;�V�<D�:
r�� �"��R#=6�=	���+�	�[����!'n=Wﺾ�'<J�5��żOy=��K<v��<0=TB�;.�2=9�Y���A�<!�<!/4==�r+�*��uS=Z8M�i!=Z9;����u=��;���*��%Fe���=tGͼV�c<��\�,e<^�;�e"�ِ=ɂ=@�qW�<�O�;|=��=���;B
����M=�m�<�]� v<���Z�<Q��_�=2�a�yk=r�Z=C.���)�<�'#=�V�<Ϟ���͊��?�/B�%�E=[���¶<��<o�t��i=��9%�����;�B�����l�� C<bI�[�%�,`��؆
=N��<\�<[,��W��_=��;��h=�=#�Z:��ռ �Ǽ�J���0�<��/=n�k<�2Ƽv�V�$�`<��2j��;��K�a<�T<��ۼO�ټ���!�ʺ2�<އ,�`8B=$�=�����Ϥ��It=�ݖ��l�<b��;�=!_�<ه;y2�Aq!����<��P���$<��'=ͭ}��ɼb�c�@�b���D�5/<A̅=pZ-<T��<�\d=f����~:����l�D<�)�����I�q�.��<!i���i�R��=]\<2�=7�<���;��C����<.uc=I�=^9�<D;p���(�7=e�.<�<Zݹ�#=���<��=�lм�7=�n=�Q�<2OU����[��<jH�:����+�<�?^=�*,=]Uw:�8=��FQ�<��;=�6v=�� ���8=��<��&=Z�,%�<��[�w;O��3E<��]����p=��(=��=��7=[}=ٰd<>HS��(3=4����<�3;��<���<]Y���2���9<��i���Ѽc��<�@n=��<h�2��I �C��#=$yE�|vu<�k����<L�9<��K=�4;�ܷۼ���<�?�����^��������#��w=��"<��缁��;�&����~�x=��;��%�a=�O;��߼g�1=���֒�k �<��"=f�=�aż�_�<�QX�O�0�2j�+;'�)��d,=��I��$.����;�g�F�~<05�<xQҼ��=�l�;��<
L@<���<|�Ƽh9D�͈i;#^z=�W��L#=H�*�[��~?��j$=�s<��������ѻ�<Y�<r�<��j�P�n=�}&=с�<��������;\��~=�侺񕵼�`�=�n��=�˼�I�;��<�G(<���;0���9㡼b�<6�O=��<ʟɼG�=��;�k<yE�<��%�!��WU�D\u<Z�q<�8�.��;7g�<Ħ/<Ո<=�m=1�^��R�< ��<П3;�ƈ���-��r���N=���;V<�9m=AjW���V�
�ռ;�<H�a�x7�c��<mtZ���F���<�%;�@�_�}<3j=5�!=X�꼢D<y\�<��\�&W<��㼳\=\����r�/bv:��O=��=;�=�$-;a{켟�<a��<P�;=8[%��r1���O��֗�,=��,<�~��\MԼ�� ;1Ф<K
�%�]��<ҷ<S� �Uss��)��{%=;)�<��G�}��;���<-ˣ�b�T���3=7ڊ��I_���>=�W˻��1=����f�<%n����= �<nՖ�$+<�r�<^a(<�9$=K�;=�yp��TI�0�����5�
�n��<�4?;��&=�e��j�һ����==���9���1N����<���F��t�v=��$���K<{<��$����t��;�����1=̍����B�\�]<�ϗ�E����<N�m����<{�O=u����@<�k��<&� �� �W00�e�\=�t��$�@U=��#�B��;bt���5E��z<��=R7l=��L���������ʊ<e�Z=����̀=��J<��O<L����r(=<� ���v=jsE=��d=q;¼�����A�}����\�l�@��⻽>�<�����H="Tn�|�v�]Yg=o���c�����]�Z��gT�;��n=��<�%�n�'=�.���=�8�hH�<  ��A;&m[�]Y����>=H�=j\����U���e=÷����1��#��5�8�)��<;�=���</�g��s<���;��=�Ҏ;Z�4�7�<C*�o7�<�@{<f=������<�(1�]W�<+)!=~�
���<���;���<�	�;Ge<�v��1)���;=�a=�%K=��(��LE<�;�dG�\��7 �y⁽�ü`�w�n<�q��P=��M<����6@�9�5�>��<���<P�/�1:t=���#��7�+=v[\=s�v��Ϟ<��=�SN��qD��)=a�M�V��ܰJ�߂`��k=��<�ؼnƴ<�{�<�ـ<!���Q�s��<�g=��9�u���
���</R� �<n�D������|;f-8��I=��;���<bXؼ:1+�(Y��C��=��!=w��DӼ�>o=!'�;������n<�;�<b�����uT�<�rb=��=ԁ;W�I������9B<mc=F!�<�h漍zs���;��<L5<��E�]���y'���?��3=�W�<�����V��U�=>��z��<�_=_�=fe�<�yt;�J���Ƽ2G#=�'��o�^�u<C5ƼK�i:wt(���\=0=�����j=𴳼�������<�����<�t�����¼�і��b�m��<X�%�@1��	��Y�=�A��W���ް<TE=ΰ=Fzl��u
��A-=2B�:�Ӽ��<�b2<f2黙�<��(=*_r�2ȑ<�@=c�������g=���j��<L�μ��Y=GO6�5"�<��<���<���7����?�BS��;,��c�a=Cvݻ����F����w<��G;�~��u�Ӽ&#Ƽ�2=ǃ7��'=��j� ,L�M.=�
����L�@�=qD�<�g?=%F=��߻l�׼S	�<�D<�Xg;�!;�A�
<_����Q�;
��<��������z���y�i�X�\��<'��:`=������<Q�����I��}�<[�.�<I�� ���q[� B̻<�*=���<K����<&H=G_�<��5<�*]�S��	%������2���j=��a���v=!��<�����=���<h�����<ο�<d9	���Ѽ;�vV=x�ͼ��D=ܩ2=C˙�~"I��M��xtƻ��=�h=�U	�����0׼-==�&<��=}P)=�ļ����O���_=9m=§���=�y��ݲ˼g��<1P =?_����ٻ��j�2����:2=~�P�^r���׼��;�;<?H`=]��=�ս;�w�(4�<=��<2<�T=�=Y=xkV��8*=[R=��z<�,�<B�1���<�Z!�+��uH�^S��kO=ص=!�NT��N����;H~�<����O���H��:6=4�X<�H#=<W�<�d=�&J�����3����zR�D%f=4ם<��=�͆�h��;�+���W��]==�ꤻ�����=�L4�sg�^QG8t�n��a�<�N=i2�{^�hᴼD�<�X�<%>��40��=*E��4X-=}ˍ�e!:��%���<l1B={4P<����G=�D�Xҳ���i���I�Y;5����<!Q��qY=A}�<��<F��<;��<'�<w�>=��1�F<xw߼!�<�30;�A���=3�<P��r�k�%��<�:�m�#���^��$�<d�<y��<��估5`��=�(8�5H3��@==m�3=� ��֫�7/�;wO<]B]<�z��e�*=	�h<�<�4(=�!;��I��<C<�̼�S<$S)�+(h<���(H&=�.��	Y�/R��d�!g�<	(�4�\�e�%��3<c�<��=��6=�9=G����`;f����;L�*��d�W&��� =�9=;�a=�����]=T_�^����޼<�H���=�Z@=Կ�JY�<˼�,r��0"=���;p�ϼe	=���<�������A�Jq�i�=��<�}n=l�=巄=�PN=�'�<k�=� ����R����V<��<%8�/B��U���=4�]=�Oi<�؅=�]���<��E=�[�w�K�~�i=!���_=!C���;��ؼ�_��>�==�g|=���<�b�<j��<ϯx<js�<�C<��'=��9U�6����DQ<1==��;�ˢ<�(=��(=�oz�2���F5r<kKG=мO=<t=�kQ=���;&5�D�<��;� �<�o���=�	-=]a@<�S<��<�d[���
�8=��hv=؎�<�/]=p�K=z�=�����߼���<��<?�&=��@���[�ū+<�����X=�T;9=�J�����/?=�l�<��M<<��<[x<�sx<r�;c=��x=D�R=D<5���=������;�|E��S=$���<���<��=�1=bU��n���་6F���<�gU�KK<%�=^|H�.r��/��f���� �VtE�T��rF��F=<��1=��磊��'Q=�8(=��;7S��?==��H<`%=� ��F=ݺi��#��:<v�g=l��=4�<o{��ݒ�e� ==	���8=WE�<�!Q�ZJL�Gw���5�G�;勐<ϡ	�OY��\�<�E��q$�����h� � �<m�K���r��{������O=�?K=К(�T	�C)R=}<���C�¼P�=��<oU�,'=5�L=Iɝ��E��CJ<S�-B�<��#<��=<�!#=h�:=k;���w<$=A=~i<��<$���K����
=������p������{��C�<��e�R=o`�<Qϻ����΄3�̌�<ق<=<*Y��=,��<�h;�g�j=7 <=E�E�$�;�P�;�B;=�v�dz�D�O=�q<���<�`V����L�<��H�Y<t-�=f��<�09=W��e=�<��5T=�h�t�O<}M�<��G���6;u�=�PO��׋��޶;�7�²'���G�+�U�0L@�G�;<�
\�or='�� /[��iJ<�6ϼ���<cL"�EN�<W��<�o�Z~:=kS�=*[=�}̼c�<���=�L���m���<(Ld=�%�]-�n�c��)e��"���P<[�м:~/=9�G���P��|�<1�����%=/��ݎ:􍧼[&
<�L<%p����@�,�	uC=��<��>*�b��;��=�9�<�T��'���7�hW=+d=��g=M��d�=�SN=��4=|6�<ɶO�+�=�H=�J��W�u�8�<��,=�y>=��J=���;M��\��<�+żGN*=3Q=ƥ#�²>��f��g�<.<��Z�١f���;�W�=t6м�μ�8���<�
=I���&Q�=$��*3��3<�<E��5�=8��r;���������V=�0¼��<��(<.����s�<k�=�w��ME���V;;ji=U�R=���0n�=���<��<-4���μ>V��eC=D呼?;&�=C�<�3R=�S��qS����4強�)��5�<�G=�y�;�AI��Y��W�z�h<�綼��;��_ =�v��=��b�����j�໵S=�(#=�_=z�O=|&<�z��#��]���m�<>ܑ<��$<T�=Y���'<�ټ�M=�uG�Kf����;y��(μ[�<�#�;�3<�]q�U*���~P���~<i���B;3�#C���;�S�<V}=z*S�eR=N�+=�oW�'<��<�<�/7����<�ji=i������G߇� �u<�v�-j�<�}�<S��<��	==giT�6�D�]�A��f��D^���{'�\W�<y��<��;���<W�,=�?�=<��;A�!���H=&�;ƙ�p��N��=�[W�x�˼7z�;��=�)��Q�6<�E=SH<��ӻ�L<AXF<2��Tː;^u�r'˼3�%=�ǈ;;�$=�d����r����:�8s��]�)�F��Z/9	��<b}�rt �ލ<薈�TE鼡�A<�+o��=	;���=��c�@�C��2f=�v\=?L����=��q��`�<���|Ԯ��&�:��D=�����M=��^=YG=U
=l��<{a�<���<�W�"u� �1=�w�֪N<�K~��os<��J;3��<�h漴��:�T�<8��<F@꼕$=79><�"|<�i�<*�2<�V���ü�����o;˹L�3f�<�����1��L��9��<��=Wcx�cz�K�/;ZZ>�9.����<�z���g=��f=�c\���/=�ﻧ^b�am�py0<Y�߼S��<�rI=�Je�r�(;�jM<��������;!�m�T\�<��[=�]=�����3���m=1�h�(W�:6)=*�.���׼�9�<�;�O�<oG=�J=ԏϼ��<�@b�o<�Jn��\=�x��V��;�4K��0��s�<\�\�c�!������B��w�;�����ּ��q=0<]=f\���H=�c=��<rV���Ѽ�fg<sK��?^e�����8@����pY��3$:=()���V��?<=�4�<��V�;R#<1��<��m<§�<���x�=p�M=���� =��<�����8%���8=�b>=<b^�w>k=�=>�~C+< �<�f�<�ϼ�<���R�<��5��[=��μ5�$���<�.�;o'�<Kgc<�r�;��5�B�=�C=�G��bP�U�\��
��O��<Yc<��=��v�aʀ���R���<� @����<�+=T��[g`=�P0=C�e={L�2�W���:jx⼌X�����|S����;���[=�#=EԻ�VHo=�&5<zg�<X�/<8b6;�����U^� �(���D=�ե<���#q=o����ؼ�����;G���W�<S=����W��"H��N;<��^=F���9����޼!2C=ыs�	/���)3=�����/��N��<�*R=�="[=�1*<��<�q==�(��+
���ib�aІ<�������i�3=���<~�=�
�:�8w�
:,=�*E=8N,����<%��<JU2=E��<|2ּ:��P�#�AJ�;�n=Ҹ�;��<J��<1�u<wmw���B�=jE༠�C<�ӌ<es}�����.'�(T=3=�L�9o-�<���1/=����L=#1Y����<�/=���$W=�J=)L�SD˼����tǿ;�_`=��<"K��^��c�Ѽ�#�<��<��=#�<��<a?��ȷ�<'=��`=�wE����:,��ת�{�d�䈏<����o;E=��������}�<z�.��T�<����'=3��sD�z��m^�;�L���+�<������<������<��q�6е<m�A=@�\��v�0F�;�����/=K�=#Ⱦ�=zy=S�E=Is]=�=�<���O��3�Ἅ;����<q�*�5=(h���<ѝ)<$��<'�=#��<����@�_<u�Z���R�ݫ<��;#]�`=��z =�<$���j�:�V�u��F�ѼJ6��wE<t�>����+<��t4=$�"��M<��2�{1ֺ��<	����F�'97�|� 2�<yD＞Ap�KZ�<�,B=\>���Ǽ�5ѼG =3����<�̼	��;mq�<��=���Q��Y�י�;,�[<9=)��7��T�8����<��=�+�,5X<�Rw=s4=�8T�nK[��|-��Z�<�\4=,�L=��=�Ƣ�}B��7��$KC�כ�v[��Du=0��<ȁ.<$n��Y��tO;�Q�?Ƴ<+(�<���<w�F<�=l�4^X��=v�)=���<�4���#�;�)��u�.P�L+�<��|=��u=�yf=�s�<�tV=�O,=��<k'�=Oy�<��=��J;�1p=��s;ҝ�<�]�;M�=�_��J8=Z�ȼm��tC?=��W=]]b��Nμ�������,��S�+�*���Q��"�<�p��$�I<���<�y�0�+=uF)��=?&)��'H�7�=�ӼrpN=3�ɼ�Y_����qOh�
F8�o
˻���:�ƼgM:=�މ<��E��=ļCvI;h=�)�;�dF���<�0H�zZ
�����=B<�=vPa=2Z<�۪J=W^�;��E�]+2=�=���Y�<���;ڨ:��1��sI��U$<k=�n�,�0�QJ=U�:�6+���6{=	,G<~g1=��P�6���=�<��<���Uh=e���|񮼘#�<e����U�9�U��<M,����G��6Ռ<�.=^9<��:��<)_5=ʇE=|&/=�W��C��<����\�μ��<vC-=�IѼ_z��2=��=�nb<5����.�<a�&�(�<���i��;��x<��T=L���"��N=��=G�-=����<��"=nG@��<����#�Ü=�Z���=����#=[=3$Y=�=��"����<�� ���<�(����u#�:��==[-><�+�v2��.=�$C�I�=(<�I���<�,���=zy����A�eވ��3��kƜ<0�[�9�<�4<�(��~���\W�;<+=��_< �����d����<�ݜ<@e�p�;	f�h�<�`��� =�(=�WB���=!i-≠z���0�m.v=��&�������;�16���}�/+=��=
p��~�M=��C=Վ2�뼕M�������С�_|-��#���M���C����~�<��c=,��IGf=LHX<yUD=�R������d;(��c���<��3�����<�>�C�I<�V)=�~��;=�O�t=y�=;X=Zq��l��2=*�1��pʼ��V����<J�;Ds�<j�<d1=��7RW<��<3/E=?���Tȼ}�+��D�;%z��)���^Ӽޟ+=*6</|�<<&8���X=|滼�=Y�9;����c��E¶<DJ=�`�<;�I�;g�<��6=3s|=�� =bW�<K��� �<�6��d�<�05<R k<D�=6%\=��R��TE=7�p�)�?A��r����kP=os�<��^=I1<N�=�^<���<_7�b�:m+�+(=�]k���\=��g=�=^�<3=戡<�b�<͉���=�8R�	�[��X�<�c¼N����;0�W��l�;�ȸ�#��f���́���C��\�Q�˼�	ܻ���4^�=�7���=��Y��~��j��/<�=dH;��1�ޛ=N=�ȑ��'T=��(=.�K��=m����;�3��� =w�
=�_�"I�<cyN�),�:f�<l�9=���EPq�vT<Ԃ�;ǿG����=�5=ya�<�y�����<�y�<I�\<8j�<���}�%�NS���1���=ɘ���n=�ȍ;@��<]򼤾e��A�+�T�'e=�B=YS�0=BpT�UR��������Һ��9�i4�<�����.G<����]{=�5�n*P=`��<@;���/=cZ!=�->�=;����<k��R�A=L�ɼ���{�
=x�=z�=*�,�Bh���d=����Eo�(X�<�==Wm��1��#$=��<��u�(d鼡�=o�����K=��7�?�=�)=���G�Ք=�(�<�*&�ZR8���������I��<&=)����<��<��]=�dݼ^�O��4;?8�)�y=�c�;��=PV=��Y<dL���P7�М�<T���!=1#�8�t�`���y�T��(�<GnI�We	=�С<��<V�P;@S|<��;T��<��<�/�<:I2=�7�<N�� =�=��q<�{:�a���.����G<]*/=��0��;�`=�;:=5���=���\������b<V^�<��9��S�����m$�;�;e<��1=�tT=);H����9�!�݅��!��<H�0=�)9=]b�;�*={w�:nq[��~�<��N<ൾ�_�ռ96<<6Q��¥D=�T=�⇼GS�<![����
Oü�� =�]��Y<����,= �{,==�-<�s=�ݻ<��L���3=��'<�=�A㼙Y,��e=+\=�F�<���by<_v��C"-=�����C3���<Z��<q�<�q��N�"���=T��Y�<������<H+j9G�=��?<\�y���<@3�B5]��<ʠ�5�==��<�

<��l��|����},��[=&��<��a�V=������=�A��ƹ�<"�<�n�;JƔ<�|O�{d�;0���"��+$�<fP=�
���ļ^=i1f�gY�<3�b<H�G;;*v�9:�<;���*=}��9Y{<��R��	�<�?=q��:�G�:8Xk���=��Q��O:B�A�LPü�l�7�~=#��hҺ��r��6�:�O<Ī˼L�
<U?�<��~<i]<���i�8�>?\<�w�D=4��;�f(�q�<�1&=�Fһ�q��ZH�<��'�E��<b0�<Rm�0	;
�-<� ���<�h��SC��c~���;6
���(<��]�W��<e���(x<�<��]=$�Ȼ8՝<�&B=�B8=L}m��x=܅���=&���j��d�u=���<ͦt��F�<�:�q�<>:X<���<V|v<1�L�F�9=�X�<T����S���R���I=���a =��ڻ�<�]�;p�S=m��<o��"��< B=�ɼ%|��
(=3��F5;, �<fEH�+��;��<?*M��4��'�"��<j;	=@n.�]KB�<:�<��l��<i� =42H��v<�?=i��&��9���=^���+<����G$=x-�<�th��J=�f<�7=����=�>(����<��^��|���O�iYټ�)=
c7<�=�T�;���<�Nj=�?�V5�osV<�cȼ�ܞ�B�Q���C=�� �<�<dĴ<�4;<�n�ʻY=����7=J�:��<A�<=B�߹����
َ�<'`�����^�f�U�;wT=����_ꦼ|1�<Zr=��B=��=%��<Q�|�b ��ܚ<5����(<L�D���<��<��RpT=h��;N�=h��I�,;�b��'5=l��;����3T���I<���*����cy=[����&������`_=�0�;�����F=4S�&A��  �<X4��qL�����ir�:���.CT=�p\��=���q�<NT�;�.ݼ����G���v]=C��o�<g���K����=z�9�dA��r�ڻ��*��4=o�d<(ּ��<��E= �.�?��<!1?�c�Y=>=u>Ǽ�8v<��	�o*߼�8=�*=G���#>���%=خ9�� =eN�p=� M<-�'=E�<*ؼj�P=24�����(�$��Dd��8^��޼�.<�����;gmB=˶`�������=s�K�1s=��<�)�yj1=n�Z���7���<s(:�_*O��F��.#��{�<Jx���x������1�<����������<m*=s��:�;5X9�?U�'p=�x��S�	�M5�=<=wow=ˣ[�qe=�rSG���/; �=�$`<r��"���sv=HTI���,=�]w��}�<�b�<c�<z��?f�<ۦ\��_6<jA�M5�~;�<54�<i��<
��;(��;� 
�#�<OY�m}=��Ǽe2-=hh�<X �<�<�}Y=EXL=�L
�PO>�!͢<Į6=�� ���8=f�1�(=�uq��{�<���<at%<ٛb<쫇<�ق=uJg=WKZ=��=�[�\:-M�Ӗ:��;��ZF�f0<z�j<�耼Ԋ�<
�=(S���r��
=4�b<��)���%�p�s<������/��5Z�0�=�Jg<��@�BG׼4ʛ���]=��:Y]:Y���/�@��\1=^��<y$7�O��y|�V{�Wf%=q!⼬���S�J����<kd=ځw��:X=�X��6�=ռ<��;�#=1�i<O�I�%��<�=�ݠ<��}='�X=��Z=w鵼�1=ݳ�<(��<W)����=1�'<�	�<���<�y5=)=3G=�����S=�;����e=Ѿ<l�<)�S�/ �� ����[���K�Yl��.���+Q<H=/��:t�Y�̏4=��<;�ɼ�D<��:�z<��a���#=���>�x������<�)P<�pg�<�`=�\s=�s&=f��<S���@��#=�Н�Rw;y���d���߻���7�%�<7��<��N4�Peм!�=�u���K1=��<�3 =�U
���u��&B�&4<��M����~=����Ӥ��W�Ѽ��ż��v=F(=b�'&�<�<���'=��8���_<+�.�\m<�|;$�?<�ۢ��4�<�����S�<�)��M�����i����<.r�<�T��|�v��;*�<��<�뜼�<�l<ݦU�7��;_���3�G/��><O����<��U=k�n=���[f<�e�<���;?{��7�A=�΀���G=�h̼������<1�5=��T�.=�=�}r=
�H��s�<
���Ǵ;$������8�<�I�<g������<��ػ^ǧ<b=�ϗ<�{S<(x�;��{;����'l:��׀<�@���Z���~�8Y��?A���C�ua����1=)=�~[��5��1���	�=�s��<눗�z���AE<<�6�wTC�43=\XT�b�ɻ��7���W��A�<��9=&�,=q�W�k%A�:�'<�j���� �<I�ݼ"������=��F=��Y���<���R�%�/!�"`(;��G��o�:��N=j���o<ҁ�<��=��=ǫ=�ʻ���,Ѽ��;�p�%=_zS<h&=):L=�ɒ�t�=/�a=r�z��g"���7;�<	�޻2��v��<$;�=���<1�N=��f��<0̢:N�A=�s�Lȼ�5����q�>W(��S���5=�	źS.q=��W=�-��#�<�*�<&"'�\���D= �(=���<i��H�m<�_b���/<�0y��Qj<'�N��M�A;�������=�X��[�<)�a<��<=��;�����=q����A;0�\�@��<,~<�g��h�<_׼�.���a=�Y=�)A<��e;��7=�$=�Dq=6��F�<o'=�K� �4���?�&$�x�C<����d�<�@=w�;�)=��Bm=�0=��7<w�$=�q�<��̼��<η���kU=�7=j���lQ=���=�K��<����lfd��yX<ͥv��6�ȇ��b<|��u�<��#�x�V;��<��"=!�%��X�^�P���b� �'�'�� �<d�������%�P;�<*��:�B��l�<Xż�[U<�<�Q!�_q9=��r���ռ@�<m�<�d���	;�����e�v�=�����ǼV&�����;#� ���;���,�3����t���_��Iڼ6�<��s=Vh�<}�7=�!<��m=�Ç=6弨}F=[F�����4v���>d:�8'�$D��Ү:�p����H=���<�`8=}��:��ټ�f���T�<T��;*��<���<FX7���U���-=d�3=%�=�)/��a�;G�<I�<��	��k�:X%�<u=M�׼J�,�I��;��s�vZ=C"�Gwt<���<3���F�<{�<"<����m=8D�<6O��W�0���`<ͻ~ke=�����5�|�*�������;���=�;��l���kN�^=_M׼�����1������e4�oeH�O$�;��ۼ�f*<�&E�=�Fo���=<L =X���`���Y:��P�<�޿<��<Q�=>?=Ko=-��<.�<͑%�����Hμm�P�0=.,0�N���<!wj��g�В<���<1�+<};<��]���k=.�<��0�Gؔ<ӭQ�o7���k�PUл��<R�S=��`=��=��;*����<�DO�W����Gļ�h����=�`�<����O�8<�!���{=�B=��=�w�;m�=D��g-=Sg��~=�o���F�%`,��ȯ<�7��y�:!��;#�E<���ü��=�e<N�<��	=!hj��b�<l{�<���s�`�</�`�^qg�m{y���;��<π<�J��<��P;�g<�U�^�e�L�hW���򻼣&v=b�$��Ȧ��8+���=:�E�;����|f=bų�L�<k�=Θ�<(����#�4=g��p5=�/<�N���D&=+� ��U=�B8=qb���*T=��k������< �;�V=��9<�2=��<Z6b��>Q;����y���;м�o�<�홼}�y�����*��v����Tu��0�<P�=&/�r']=�=��������G�8-=��ȼ8�]<��-A�0=��;��_��(=\q�=�'�<��<��b=n]U�#�I�DZR��!�@]M=��˼��=:���:}(=�-��^�=�⺻����]�ϵ�<)��]:`=��R=�~Z�W뽼VMR�R_��	9=$�:�O��9�a=Ӓ;ݝO<<Z�<2$M���C=���'� �L9��X_��м��ڻ� 6�(��+o�;�#��4��1��*b�H}���:�юd<���<)�/=�?D=��@=#�J�!���ކ���`�؟4=�ٻ�c��[<����Ԍ��`}��������Vr��	�����<b|=K�q��ix��61<�_=z�&��h�Jj=�B5=�~�<�n���ͼ[ <��&�=�.��0��l <�"�=m�:���;� ����G=��u<1M����<A3=1�_;,<��*<Sp�:�Z2���;�+x=�-���aF<5�=%B]���~<��;�����b�R�6�O=����8̼��'�Pw?=!# �m�T�R)={P�<�fb���Z=���<
�W=�Z;yIH���¼c�����#� �.�������d�앯<]]Q�T=�㎼ߙ�<��#��v:<s9'<�BO=��<<櫻x�1����FN=+��<�D��������=́<�[ =-U/�b�6=��<�3�;�@<,8���9�Nc=^�C;+IQ=�q��"�;�i�n�_�v;%&B�;�<��<}�{<�[=�9V��i`<b@3���H=ز⼠�N=�l,�h%]< AB�:u.�����o<�S�<#�߼>&�;���;�"��=�<3E�����YX=�؄=]=�=�z�<�.:�����mR=\X�`w�9(8����<3D��L
\<��;W�����N=	�t��=q=�^���Ļ�W�<8t�|XU=b�����$=��hZ�Z�2=X�k8�<�e=z&�;u�<~�<�MO��Ĕ��<���Y�g�<5Ǔ�p�6����:(́<�E>��ʬ� *��Z���:�P��u!=��4=�z;ȣk=�xӻ�e:=�h���)=��;d�V�'9�s}���p< �ļ��<V�[����<'�ӺN�����/[=�!$=���&Ȼ7"&�(:�g�L�5]V��S�]�H���G�Rĉ;]5�<4��<�Z(��K`<0Լ��H;��C��{!�3�a�u]�D�H�<�����Ƽ�S^=3/���-=ޮ�KC�;^�һ
zV����� �r�#��3F=��v��~%=)Y�<E��߇ =�L��O;?\���ּJ���f\μ=��[�	s�=�?=���C=��<�K¼.d=�b<�1E=���<[�9����<��<1&=��J=c�<�{�����]�N�A=�QM�����=-X��uع��<n[!<u�;  =k|�<�f6���<��<C*<��~�i�ļפ)=b��<�d���%=�O<=��v<�n �;2�=���<a�AAU<藃�e%��r�==��Q=!�ؼ�;J��36k<�R���b<_�;��<005=Gi<�wV���M���;� L�<!���I}<[��AҪ<<�1�<]jǶn<�����K���Ѽ�k=�f_��P��+�<�� ���=^I���Ϻ3�<�G��h�<�e\�N�Ҽ+��Zp˼��3��s�<�Mo�tr�<�2M��aw�^�<�3j��t<�}�7�v%=VX`��G�8I���(=9�B��B��1U���K<��<��<�g=��O���S=�6��x<��|u���2=K�y�ּ��_=�~=�s�<t�4=�<L�o�=	P&��V/�TW=�
0�;��P=R�+�������6�Vq+=�i�<�#=��b��ռ7�;���W�B!����7D=��|;���<�����&=�Z����� �<�\D����=�=�<�a��}=���<jO�<=cS�*��<j�O� ;޼�=�>�<�>=˥8<�g/����<,A��D= y�<i-S;:��<�q���a���N�<���;�<!;��;T+d����<�u���ࡼ3��<cFW���<���x�S=;����;DZ�;_����P��lJ=.	�<�:��9=����@=I�A=o�2���
�:)7&=b�˼V� =g�"��&=�/�<$�μC ;)���B�0���R�a��;��<Kא=b<MT��y�<$Vk=�L���Q�;�Ȳ<� ���
����+<=�&=��1��=�we���L�qBT=�=��+�7Z'��P�ё�<�wB��L��G#��N���+K���h�QN;��D�<�n=HԢ��|;��h�߷�b3�������C=�M�K�5=@�<=�I!<f�"�K�g����A�˼��
�A�<�{Y���+�|2	=�<ټ�� ���`�f���W-���f=b�����܇w��[7����u��z��l�<��d=`�ܼ�-���?� �V�: �<(P$=�lX=�}<��=z*=�;,�	=��|b����<m=I�r�2�AO��� �(=�X;=^�=�E�"4=H	����;Ʋ�<WP	=��n=(��T���h=��6�����=�x��;Cw���;Z�`��3N=�h�F�)�{��<�<>=��zT��^�<h'�����:x:�=j]9{{��]���5�GW�;�Oμ���_�`::;Q�<�Uf������X<*�=��X��bϼ���<)O1<�ƻ�v��l{Z=ġ(�!��8��qͻ�E�0<��x=�w�<Gd=������;s<i+��<��H=~�2�����w�b����H=��K�!���?��2�����.+�x�=���=z�Ӽ%�/�Ue�=?���c�<n'*�9�	��<E�D=�v=��5��Uǻpc�2�#�#
N=tIh<���<��	=��<��ݼ�ي��=���i��<8*�<f��C=e�=���\< �<-~=�l3h=��n�f�(�|��<�&=��<We��M<�m�<X$���<Y/������=m��<'0�qm]�}]=��;�G<��Y=+z-��Ƭ�Ⱦ���3=(�<T�:�N�a<ʖG����;�ǚ9QTS�ď@=�a��`=���;S\3�5����H;\�e�>� <��N�vL��n���K>������<�K=��<���<�^a���:���;��8"K;=K��;��������s�m��)�<"�n=�z�偲;�)M=��3<c�[=�*����*��	=�g,������"�<x��<v����&�� nt<Or=bqo�w~]�:E,�T��V	�<�[_���T=��� ���I#O����ρ�=�AD���e=�;�i;�F��ʦ�%�n=,�/=�D=��}��e�<4�<��(����<��C���z<�*l7=Ʊ�;_� =~��c�<��
=~��<����#��^ۼ�=@x�}C=4�;����;���<l��<���X=%�]=�=v����n��rm��A���j��A��c��g�;Kbӹ��&<x0?=smѼ��4<�!p<���<�w�o�=�
"�d�,=`_�<0�k=��G=]5�<a�<f�?<\{a=D�=B���Y,�H�A�%�@�C�ټ�b<��T�;����1��n�.�W;=�F�ʍ[���I�A�;<�I=���<�a�</	=��~��&���г;��&<�᳼r����O�%�.<��<��F�DjӼǦ��-�<�ҁ=��{=�C�<�m0��i�<��ǼiH+=6|�e��;j�����A���f<)��;V��ѣ�*��<��ż��b�u�<=WZ��<<��g��+#<�څ;p�X=9�R=.�z<��|=��j=`��<^�@�{����<��<u繫D =Э"��y�<�S�=�@����<+'
�peE���@=��;�w�)���U<��4=56=㙼�2=�9�1=-x(=?�p����<D]T�h�;A`0����<��D�)��i.=��<�+�<#��<�|G<���:��<S�>=O�<�;���b�<)���i'f��~�<�ۍ�|�o��='�j"=ʱ����T<2Y�c�Z��ѵ�C�=թ�:��=ĵ�<�D���<!�=���@�k���"=�2�y��u�Z�G&=F��q��92X=X�\�x�B=�6=���8��<ռꨚ;Ͳ��B%�<�$>=���<,4��)˼j1��E0
��3=$��<f�m<�2=�%M=}�9<O3;��<`���WV8��R3=
�x�j�Q<��:�<@�Wυ��P9;KД<F��f����r@�<Z_.=9�G=���;�vt=��)<Rs:=лe=�>�����(��P�9��e��W<��=���<�������������sE=;j�<΁�<�/��H
=�����Y�S��8p�%���%���BL�<��=�{�<��;<�XM�Y.���Y=RU=��<��<�KG=۾B��?t=�C�[Ɂ<A`ݼ�2=�b�����:=g8��Ӈ���X�i�F=�O+=���<9DF���h=hT�<�h$�	p�<H�Y��K<�+��v�9��<�y�2���G�r(<�,�<���Ei*=�X�9V�=���<�u-={+<-�ͼ�*
���R��%<=h�Z<�B���M��N�<�տ����$���h6=/�=�h=w��<c-4��I=d�<�x�<�ݼ9���[{l��/=�v��&:�/o����<k�<;Ho�N&=Y~�JW�o��?��;2��<yPN�8.�<�w�ֆ�;˵.=z�:mDg<�s@<�I�<}�=o�(=��=`b���K�<y@�<#�<��`=�h�����s�D�'=8�j<�g�;e�G��0�#�7P�l<.��&C��;���a=��<�*���������=�NZ��ü��T=��C��9�<�qf;1󿺥,������;����`<����l.��M+<�s&=4��<efU��Bo�{��	���05=zt��yC�:��<���<¨=�ڎ;��$=x��<Y��=&�(���_<��X}����;R�<��= �����<\�$<��=m�>=�==��=���;H���^<�pj=���� ��;7=0���<2D��k�V������żT�?<��`^=�C�nW<x�<�a=U�Ἕ��	���/���=����^�żF;�0�<װf��j=.��;�A��/�Y�X��L�<2�k,M�,=p5:�����JP<�O"=�DX��0����3���û�U	����<��I���,=Ts�̭<�Z6=��;���(@o<c|���m[=��ż�=Y�ݼC�=s7�<n���t�v=�vc�:o�H@�<;�� �2=g��<7�<z*��:.�<bH]�ytM=�⦼��w;ɲ̼o�;��=�μ�PԻ/T�<h��<���#O0��F���5=�r>=H9p<�<{�i=Xn9�ƍ9=�u?��O��y0�)�b�Y�'�^y�<�����<JB�9���:=>�|�q�n�>͠<�;��h�ҼU\����:�y=��1�6���w�<�:�>o=��<��"��ı9]�8<o�u���;��>5���<B��<"�=�[C='H�<��z<�]<Jr�<����<)���O=�F�<��/=fcz=��9�K'�� f��w`��������< �.�9A�<8�i=A�;��eѼ�*`�4*=�#�W��<�~��輰GU�� C=����g�<��=��z;&��]&e=�p�<����4< ��F`<���5�ܼ�
�Y��R����=�/�<}o�z��<���<j��<�<���c��'i�)-����<m� =��6=��e�T��:��Ѽ6( =�=��,��A<9��0�e��d=W�<�qC=�+=�x;�R�<�#�:AT=��jq:9.<���=A�r�%żǘ=V�̼4�;�;P����<+`�<����5R<ɳ/��Q�<�jJ���N���l��<?W�;�M=t��庀=H ���<�û�]��>2=4ﯼJ� =�Ki�Yb�<���S�;���5�I�=�O)<���C�?��@�<���<�Ξ�^���(TM�̬;]��;V�b
ļ=.�`=�F�!	Z=���<�\�<�{=��8��cI;����9:<��?���\�@l =���[�<��@=�l=Axh=x��;�
=��뼣{���,�<�#�</�G;�Os=;8x���}��F��m���1E���l=�_=����_�S�μzX9��v�</�s�,��<�Z=1�A�ቼ<�Ha����<{=:=lK
����<4��n�=\N�{[�<��h=X�ۻ�8׼(�2�^=��o=�Ȼ'!K���=�O<6�ݼZ�P��>(��SZ=F���@'=�F@���<�٨���?=�3�׺�;�GԼe<n��ae�<�xn<�چ�,�/��u=�(h=<��z=��y�=#2���1=�>(='�z��I��)=�� �����,���6�{����.��!3��_F�7�,��#<�JU�k�L����<&����q���˼�Q��*<J��a"=-R!<'�1<;i^�(�����j�I=ֻ=&��U��<������X	��F!�{��<_��<xr��� =��,=G����Ѽ�¼;�M#=m�7=99�Z�z�];i?Z=��t����XEE�;�<m+b=<�<�f�����k`+<����Q���Y=�jL<��O�š`=?=��<҈7=�*=z<�<�f�<2A��	=�<��K=������;�}���L=��ȼ�b(�KV������<�]�<���<��<��?=F#=��6=K��<UI����������o�<����hߺI,"�1}t=�Hy<��;�@<�K'�1�=�JO=�o"=�&=xnt=u�;p���M���qS=��=X�;� ��~~Ѽn�<e��;�@�[Ҹ�>��� Z�<�P�MvQ��H/�ClS=p��i�<���/a)=�B�<F1�<®��~;��p@<��;o��<B�
��q���i�e<��k�Ȼ#���8���<���
�F�3���d�<���<�5=��+�j/���,=��U��&N=�6��ℼ=U!���<5�=jٻ�a���6�mc1=�=�*J��1-=E��<ˮ|��k�F5
�uT�[H =�)J=*�e<�u;=|~�<5=�̼"n:�HZ=N|-�.rZ��O=�ܑ��@¼+c��@=�,h=E^ �r�'=-��:m�]<*��0�N�<>޼V�{�8��.��(=8Ya�����z�L<f��<}y=����?��<�^�=��g�#F�<6=�
=�ꉼ9�f=%=�H<m��;][���>�
�-��QW����<���<�b<�RU=�8z=��?��e���;h�^�����-л���<a�K=�������;'����Yl�{���7û�G�|��<�V�=:1��=��B=sޣ;��6<K,w=��s:!t[����<>f���z���F,޼��<���m��)<��%��­<�1S�ԥ����<���=�dV+��ҽ�G_2��J�<Beλ�
���-=<_?�<�i�ƠG�6D5�4�N�&�=#"�ޭ�<��<�7Q�e��Zڼ[*S=�R��T��;M�r�$�{Z|�"�>�7�B��r"��C�<#]D=H�=�CD=,ٲ��x_���;I8 :�2#=�4���*=QA=�e�;�0!�?)<�+��0=�6����̼����G7�<%�^�������F���8<X�r;?>����4=M���g�<O�k=m�)�cj<�ɋ=x#��X�<�=@?�<�X�<�H��d�4��==)��<5�;��{�R�=?�a=ӫ�<��ü3��9�J��h�<Э8=��=&/6=԰<
N�=�"*=H�\=c�"���˼Ӽ��ѻ���<��t<���<o�~=��м�v�b�弯0=�`��D&�<��<i��<=;_����t>=����\}<9��<�˼�m�<Y�k�:�2�>4�<���=O߂=��e� ����K�ΰ1�H=�/vZ=��`?=�S����B<�)�=&ݼ�Ś<��_<�u�==�/�iki=Jû�.���N��:����=Yi�<e6?��U=�E��(�=
�<1�&:��9�OF���.Y=�s=]��nڐ<�T��Q[:�h�=]=�
=�EQ=�����=��<�Z
<8�d����g��<�v=��<'�j���6��	/�u׌��F6=��g�'I�x��;e��[~h���f�tge�� =|��<Q@H��"U=�W�<BJ�=<M=�=7���R�H<���^gϺ�/M��l;��Y;.8`<�2Z=Z��<�ā���м��{�$=v'�<V=�٭��[��ȕ�<ē����L=�?�� _<�0,<�?�)�<�n=�v=�^�<�Hr=W�b��C�:��������<W#=k=KS=6}���oڻ w�q1���V���ٻr�һI�/=t/=<4�<�ZF�_z�Ak<�y˺v�0=��N=����2<�'�O>>�@n�1>~=a��<=Z=�����<��[�m�<�ܪ���>��k<v�<9�<Pm�,U�|�t=����9�q�+��D�R��Xd���0�rx2=6��;=��<���V����!<.x6�2H�%�=�%7<��=��?��N���X=�˗�k��
�=�U�;EJf����<d�ļ�1���������<ik;�'��}^�;=���<�Y*=5=e�}�?�3<R�=k+��c�B���)<`M=;�S<#[����<�ʺ�t��3ר<��=�jH=�Q<��T�JY��4�<��ֻ}�<��Ѽ��.����;�@;Q^�<��^�bT��u�=�w=D�<ξf<���;kg1���M��=?����JҼ�I'�XO�<.�'�|l=�|�:I��<on���=Ћ;�&P=!;������<��V=���<�Rl=0��<b��n��<������햽 D��0o;*g�<��I=(��;���<_jl�:(�=�4�[䈺�἞u�<�E6=�2������G<I$��j����P�<h�߼:�<e�Һ5�.;v��<bу�/`�;M��<��;z�<=�a=��!���<+ڼJm
=4�ۻA��;���i�W<�� <�n"��L��>o+=��K;j=f�y�ȼ��v=�3�:?������ì��I�Ya�<v�>�k��_]�3��:�I�<�K�;)aG=�>���:���ϼY���/�u��=��S=|vl==�ּG�7�R�<&ZE=�x�<��M=��x=�,޼��ټ5�׼T�=�~5���<>>=yS=�l�
�9��׬����;���;�P����)<�K��L�L=��!<W��<W9�<~�������1�;�üy<� .=��F;�qU��zt<-T<�fl<��<����Q�:)/�H��<�g8��:=�p����X���="�����#�<=���J��%=��<$� <������<�~�y�:_�}�t��sޢ� �6���#=U��W6Ƽ�� =��;�L�J�&=D?y;P�4���2�q��-)�<ۗ4�2TU=r~"�C�=
�A�G����_#�<��'���k��EM�bnL��7�<='�<߰H<D�2=ʴa�{�==��ü�,==�J=�5������<�����9� .���;�y<[�8�ț�;H����=g�j=��ݻ�1=xdE�	�ü�E=,�_�qb�<L�Z��  <S{�����;��@�T�c=-`<q*S:�u���Q�5�߼ڸ��x?=k�F=6�d<�"k�cX�<tsF<a�9<E�i��"m�_0׼���<� ==&�l���t�<B�2o�ϴ���c<㙱����)�<�A�<�� �(Ԙ=[8(�8�����<vQ�<K~<.=�e�<v�=��=s�5=�b��e�9=Lу==8;���<��-=&���\�r�����<���fVӼ{v=���<�X�<�UU��=c�e����<����'���{=��꼌q�Y��o�E�h�=�wv2�Dʌ���l=дZ=�F���9��=L�׼*BμV��[ƭ<�����ټu�O�~a$<���f1�G=�'����L=��^�g=jĄ=�M�<�U4=�ju=��'<3�Q�@�C<E�;�R_�`��ġU=��?�|/k�>5�ğD�3P=y�M=�${��ߎ<�f`�U7���;k��=��n��%��/�l�)=�1��3t�<*P�<7�<okU�R�Hk��Y�<�x��ֻ�M�L�*�۪p�����E�ڝл�=W�ɼ!��<��t��#2=l�U�8��<�4��k�;���=��9��i:-=S�3��⃼�:d�G�üU��^o���z����<���<��<ت =�X�9�N�yk=� <9Є�
0=U� �f0=���<�\����];�kʼ!7%=��ڼǒ�����k�<���k5���K�;�L�+~�;A�=�dX=
{d���߼3�<u�
��,�Xj=<1�R<��:���<9qW<d�<4՗<a@=�r`��/=ϒ\��b�����;�ڸ;eL������t�^��<+� ��`����<��
=l?[�܏N=�IػO��;C]0=�,�;��X�e�<�ln�$<r4-��8�<����=��μ3����=�1p=l�S�(�=�F_���1�z�'����^Q<9G���=c�4=V}!�08;_:*=
+��bV��żr3��7Aȼ���<�-�:Y� ����λ �z;��������ݻ��$=+�H<���G��(=�o8=<<���<�q`<����!�m<p뼤j��~>^�t(�<�x�;a�M'=,X�<�<��V=Rݛ�<�<�ξ�F����<�Z;=yY =؏���X��;t["=�13���4:����ܼo���u=�&��q��9��<�h�O��B<fe��j�;�cR<�(=��?��w�=e�Y�&��1g����:���^�)}<nG<}v&�R=��<I�л��%������e�`�=���maq��b]����؀�=��B���L���t=tn2��{�<���<HJ���=�u�6^��J�>ͅ�v\�s�ռ<�ݒ=W�,B*=�]�UZe��Z\�.��<�a=Y�����<�Ď=�a��0~=@S�F=X{=T����[;��$=4h˼q?5=�IS:-zǼ�t���d�;O���g�Q=�FF=j��k�k(L�O&g�>>A=
v-�Y�@��mf<���<�q=/�<�N	�Û`=�8�6O��d6�<�!=B��Y?��=�<��<�}��� =s6 �6��<�k<=d\=�֥<��V=�b���e� vü�-{=��1=^�_�,�ؼ�<�K=��ݻ�:�<��<����<o&߼���;�����*�ƻ�1�<���;vo3=���<�: <�j=Юp<�b�<��<cI%��_g:�(0��m<�0���z�2ά��<<t$=y��|�[=��IcK��!�~�ͼY���� �;��G��č<7�;F��;��߼�J߼7�Q�]�乛�� ]N=n�̼����X�D"�<'�R�xv1�ݫp=B�<���<Psv����=d+��@�����U��"=�1���߼�'�gx=�>5��A��b�;�Y< c�:YX�S�K=	[�=~�	=�#���	^����<�=�C���=�c/<B�\��V׻6==���<�!=7I�<)7������J���e����<���>G=ehr��~=X��<�?<=�9x<��=D=N k��=x�?n�(�.=� =�*=�<�*=)�#<h�$;�L�=/f���-=���U3=9Z<�n�¼WL=��\=�-�-�m�+$3��H�=Wq;��"<^�=�R=�q1<N� =Ut���(�d��1$㼀�x��3*�qK�=�.(=OH�!bf<F0=f�;�=@es=Ih4=�<]�W�2�h	Y�{�<�#z���X=�q��!b =2N9�i=5��<d�����,Ś�fO����D<��K=�vȼ��ٻ��ϼ���<�u�<�a�����=��<!�D<h��<0\/=
,�� _=[p=;S���D���֓;2`�H�=���<=�h=��*��-����< ҅<ۯԼꭉ��J-=MT�<F�T=��=W�n<T9< ;T�}�
��;&��D�;b��<mD5�Y=�s߼�@�<��;l�><fQ���F=aS�4��|P;E��u�*=���<k<�oH<�<5����缄�:���zJ;��'�%�;������01�e�D����<b)�s�?�&0=ul+=��1��M=z��<�)!=ƌR;RT<ݵ���;=����<&�:�G=���<�����=�T�<+/1���\���޼YƼ)3��*���<vh*�Ϋj=(ʊ�9�z��	=P���]��@@=c9�;�/ <�e�;��g��=%:��x�<�W�<ڗ<�N8<�&��֗���<WH�<� �>I�ҥ��,8ۼ��^<F�S��^�;���<�lk�#2=7�o=�=��V=�딹b#�<8��� ���)�M<�9��$��<9'ټ��h����<H�&=4<w�<@�� ��V縒}<=����)�=ZLx<=,�<��V�<�f�;�զ�@��;&k$��c�Y���m6`=:�S�+�r���M�4>�����k��<iSL<e�Լ��c���0=m�b;��żU*�<? =�=�r��@r<nu[<�؆<r=>z�$
��U=�=�/;=��-��:F���6���_=
�=k�$���<�Ѽ��	<o2�@�+=��ʼ�iC��D5�����b��}<i-��=�";ܬ���I��x(=�)@�B[B<������<��< B��$E=�s<���_��5_��v�i�+�0�g�$P\�X��J�I�7Հ�~)���Y����_�]���(�QbR��9==��˅<��/<������?{��H�S�����:=U�=�4�<�C	;�x4=^+�<~�9�z�~YC=�ͼ
s�;�@=���<~]E�-r;�45=�@�9�< ��<\j9=IE�<0�*<t`0��D�<sk�<?�<�Kؼx�=����+.<۶==�o=�\��c��d� �TV��}<���<�����B<	���mp=�PI��Z(<����U�<5�<��<��-=O4�<��P=.
=mi>=�
E=z0�)}
<��ծ<�ٗ�Vr��qY����:�灬��(�u� <��<�7�;��+=��S=��Z��0��v򼼄�<�Q �	jԼ^<=5p=X���	Ҽm��<
�,�B>=��9=�6�;�˶<�2;���Z�5i>�j=��%%�<���]d<��~�P*�����R�R����.3��M��� =���:��n��ѭ;��`=�zH�Toj=>얼�aH=���;RV�D��<�X��!=��v=�m��= �<t�#=�󼇘�;1̵��<���<�t�<s�ӹ��M��?C<�}��>%<�(���.<j6�\�<�kR<pL�<�CS=^��<��]<b�P��{�;fH=R��<�h=�<�=~;��T�`]���K=�%+<�P =H>����"=[
`<83=1>���[<��_���="�z,=lk =-�i���/=x1��M�8ƴR�,���F<�b
=kF�;�$<�,�ƙ{<Se�����O�"��.)==��u\:O�޻~�l��˱���<�Ļq]��Z�]=�|/�p39�QH����/=b�m=z)��d�M�ּ����R==?�%�Ҥ<7Q�;Jz�;�.e�sE�x���%=�=�O������<L����<�;A�$H6=r�O=�O={f�< RZ=�^=u�
<��4=4kA�<�%<���;Aq�tG�}9��E+<}+h<ڬC=tIS=�l.� q���:y�V=V�f��[	=6G� O�<2�;i`�<�:�:�׹���ͻ,�N=����r��≮@��A�	����R=fh��M=#f<~#!=�]=��=Ԡ�=2Fȼ�R+;�a�-�{���$��j1����<@�z�H��;�~�հ�:G�A=d*i�n5�<8���I1���k�sL=�-e�$<� 86o=i|;�|O`=j��<W�Y=S�=���˛�<t�?�Z�˼�����L�H����L���1�)��wy=��<�aT=��<*G�.w�|�e�G��<���<6��EV=�޹�/�&��̶�7k��C7��<�Z^���YD�)=�C���=̕�<xR<�&=�T@=Ё�i�;;^���gP=�U�<�����a:��=5�@�IV=�~�<O�H�
s�<4Y<��)=Q�I<a׃=?~�<Y�<i\�<�{4=8l+=�ȼ���;&�=f�����M�=pk�^;8=2�(=)�E�b�&�8<��
�^��<���;�	;<�@=�����
lϼr�=8��<��ӻP;=�h/=�ʺ< �3���v�yy����=�.�<�X=e��<D˖<�+�c�d�����[R�V�=�2'�ϝ��>�<��=5̟�I�=!�<���b�4��]�����<��H=z�-=��<�+�<����<�U<��'=� @=�6P���<<ZX=�	�<����;M׍��e5=�Hּ�e��&��L�N�c�i<L�J�.�;�jV��D3�s�� a=�Q'�J=W}<�L@���fn����*<�<s��<qʀ<@aʻRyټ�� ���������6EH�#��d�<H�����J$=K@0=�x����<�o�<m�0<ayJ<���
�<��O�xSD=��J���<��=���<Ir޼�J��0��;�)=kT�Y;�%:6	=1O=L6<l
��	��Ef=�7=�]���kP�sE=��<x�ռ��<����+1R=�R�<;���5�g@�=e���=`g=�����U��ԅ;��b�<��}�݈1�41�tm=g�a<-"F;��O����;����n=]żO��<��A=ˏ�<�b�<�n$=:�P��b=�o=��5������;�A�I<-������i!���=�&=�5��%=3 )�	A=`�<Sȇ=a���'ca=�Oz=l�N�2SD<����P��,u=m�6=f��d=*}=�V#��YO�1cg;�d�<k�-��O#<O��:^U��g&��g�<+�Һ�8�<Z7Ɔ��%<p�8=�<�<�#=l��3�=g�<�9d=�Ȟ<��`�+O?�'�<��<�Ɩ<��1�*T<z��<�G|<�ț<�.G<�1��׆=��|�i�ɼ���,[&;��Ѽ�;=G��<.0<4�=P�9���|0W==;d#7���7=O�&=F��U�;_����$<VLݼ�/�=mo�$���n�����;x�g���"��@�< Bt<e�����B<kB��� �O�p^q=E�<1�<E�9=Uk�]�=qe��S�_�U&�r�G���r�N���%�X�5��[�<=��n�|���}=�4�ÚQ�m69�?������3QC����hE~��rh=6"C=��<<�J+=��;�,�[<��%=��k=�<�3�rx��Q=Ӽ��1<�i���E=x�9�U,'����^�J�� �;p�%�X��'�=�W�<�W=݇4�{�:���=eb�<�+���=^�u�Mr<���<TK�;F ���=�WJ<7]���\aJ=�g���ʫ�d��.t��{��/�D��/�Q�=�<�"=Z}=	��	�<nP:< a|�
�G=v7�=d�=�7:�  �<^~
�1$!;��;MN�-廚�,��o�<Q�3=�:%=[Y���Ի��R=H�I���Լa�<�_q�{l���>�f�6="IT��(缛�;�]�<�ʻ ��˿���2�5���lr=��Q=��$<�~����c�\q9���F=��r=�\o=��9<M�<D�*wͼ60�<2�N�s/�ŏ�;�Fڼp������<+��<EA=�&-�W�2���=��:an=�"F=$<�<n�;��I=1�8=u"�<1m</��<A9һᲊ�ܥA=q�D�6;�� %���v=O�=��8=�:i��6� Y9�K��I�F=���>*�$@��伛�!�!���A'����:���Y�<���6ը<V��1|ټ����rV�;��@�\�ֻ�}=s5<��:��<Q��<s��<ys�<$��U���\�s�S=t�˻�ކ:ҕ=�8=���E���b=9��;X" =btX���1=�L=X%\=�u#=�
Z<d_�Mu=6?���6:�P��n�T@~=��=R}x:�ؼW��-%=�#�;�P��;P���!��f;�xi)=�;�7�<�"=*)^����<�ћ<���Z[�rt�<`���<%2=n����d=!�<�y[<ډF=bm=w&��M�r�p�ռ�F�<<�-=��Ѽ^'D=��Q<�Qp;�-�1O�}�ȼ�_�<�=��C�<՝�"����ܻ�j���=Π�]%׼��<� �<ۘ���졼'!5<QuO��o^�!@�@p<�MG���.;�]�<i��<�:=UJ4�v˻P�<�߲�[=�ֲ��7a<��<ĝE=w�W:G<�$һ�S<I�Ƶ=�U�;���-�<�Q^��L��V=�^=��w�8(=��x�^��G*;���<S=�Y:��e=���<ֲ�.C����H�K�캥�;7��׵M��\`��Pt<�Du��<���Y=Ů2��'=�b<Q
F=������<"6�ܻ�<��=!3=��<��a�5쥼n�Y=~ׅ��xV�
Z���3�DL=�Y� �<��c<��9��>=	����sB��~%�3%�v�2<�뼭W2��
���(=��'����<S)������m=�续i%=�;;�=���;��(��=��+S��P��HL�:]�<Y=����W���;�� ��L<J����%='T=��|�	@6��|=Qc	����:�=m*����+QA=O���M\�7�E=ș�<iH[<>�+=z$`���N=�X����(=�IV��g� (]�C��<껥ϫ<U�'��=��:"S����4�=�*J��@�P��<����h=��5v��(�<ד�����<�;<���<^\;��B�����fy�j�<5]�<� �T�B���b=9�����-d=��8�,kT�=pm��ꇼ>�3=P�(<q��<�8=����7�x�O=n�_=�%=�yJ����f5���=�|N=��E��!�b�!�}GE=��wi��B��<L�"���<q��<%��;Ϛ2<��L�?X����<�����<�wa=��ż�e�w���R=%����P�N��<��:�"��p�8}QW<>���+���_�xs�<f�<�nH�q����9= �!=�K���l=�B=TB=�<6!���%�f�	��EG��\���>�#�ἐS<��B��������;�|7�Q�C�h���{j=��s<Dk=<�w����;��C�Hq�;�h=�!��a�}�;39��W�B�-ɧ�8�b=�SO=�=yS�<	U�-a���<x��<�^T���ؼ[:�<y���L�J�ۏ�<�4=K��fe���g=��5�
�7=�c�uJ�<������}�^L;
�U=>�ͼs��A=�;! =Nt�����i��'H ��rg�JvL��\<�x�;3��;,^N�o�<VN<,:=*ᘻ����`���ɕx�?�p=|�L��PM��M��� ���2�}ؼ��}�;F��������]Ȁ;Č��8�;��=4`�;W�P�V����d�<
h=��a{j<#��<f_���gW�Z+f�m�{=2=�\P=8��W�!�$�
<��`=�Ms�s3<|O-=8=}Od���<�Y==�7�ު0����;|W<=�_1��xE�tf,����<�4J��_���k��TT=��u=N�=���������:��m*=X�4��p4=��=��U���<�G�<ڟ!=�M��C<�X=:��m
��<z��= ,���1�;$?	=+i�=L��;��y��*�I=W�:���<�?=N�̼�=MO=\I���?��
�<�7`=^Y+�[�=�69;[b�;D�i����<�9�</3�<:(<ڬ�<�!x<,��Gy��A��ټ����U/<H��K�]=�[�<�BG����<�!�y<~;��<� c=l;=e�T��23=�5����:�;���䗧��j;�_=߬��#�O=��D=<wT�aVI<rn:���&�@��Y��F^�Eh:�9�4X ���H�K��:~Y߼��<�wm=�;��ա�.���镼t�i��EV� >K�Ï�b�<P�=F�<_��z��;�l�;.>����<*�:�|��.���@����@@=�t��H=N��m2���v�<%s%=>��<}>=�J=~��v<�T�z;=��%=�;o<�'&��@>=�L(=�H�2��=r�!�!�׼�����={3/�I;����=�C<����ɻO��xG�.�<��9�-���U�a{%�zc����D����<�����f�����B�&;����f��@=�3���N���Q���4��H<=�G<�<�ͼc8=ou)=�^:u����t�貼�Lv<\��(`��4�=���;r�=	&C=oR!=�� �m<�]<$�C=\��<��m���� =��o���:���P�P�_���8�ۻ�\=������;��<���	��nP=������<�K`��2A=yQ�<[h�{�=�W�<�uC=`�O=�E�<�y�;�)S=�<�cpü�;��U=q�q=[0&���`����<�x�<n\���h<�b1�r�=�A �f�J=��d���9=�z?<,Es�M�$=Y|=�͔�"�B�!{7��c��d�<h�h<�%@�[��v=]���4#=AS$�1�t�B��*�v|)=9����v
<fJ=_�=��?�F�<1˼�L&�#]W=�a����I�צ=��o<�yZ=�,��S=q/�<�N=�� =�G=��V�;<��ϯm��7�<�o=I��3o<6�=��-�=���9�<�J�{\h��9+�x��4=��=*�4�t6=~�<�YP=�5b�#^���<�26��A��Rq�jǞ�����btc=�r<L,��	�s�@�3��޹��4���#�|W�<�Z�;M�<�Z5�����8= -g<W3I��*N�s��;��=֏<�C=�u�vs5��C<5��������<6d�v(���_9�'���+N=7^L=�_�����3�R=B6����)=�.�a��<��p��@<kb�<�s=5'/=���{�Q$=IM;:�]�o����v=��<�A�<3�1����<�F�<�^�<Yd��L��=�=�0�<�-�:�V=��W���Z���<e�=�Dü��)�vp=��o�T,Q=n�5�;��<��Z<�ÿ<R'=/$:�F<��g<=�#�B�(=6�< u= "�;x�W�?-�U�q���<�N�M���R�J
��2.<�!���􍼥�M=@�<�I=��>�*ļ��1�m�= VY<4!��� <ѩ =��=�%#=���<El仐C���j�=�%��L�<�[m=>������=L�ӼAAG=��I=�'����L�<�	:=]�͹H��=��Ц=�d����;`�Żލ������.��<��y9��G��'<n8�@qQ=Mm+=��J=�i]=���a=9�M��<_��:�������)�輭�;e�`�R'����[=�-^�}/.<�P��2�"���;=C=�hs:N�w=�D�<�ԉ<��U=_�p<�o���j4���c=�<<H=#S<��0=�w-=�÷<�㫸{�O��?��)J���
��M�;���{0�<<��W�?���H<j���׹��׿�<sQx�&A_�-�*�%,�z��<7U7=Q�o<�F2���w�d�2=.�-���)=Dd8���j='�=ۮ�<
��*����1=���<4[j�y���6=|f�<��\=�g*=Q%~=)�j=?V!=A4ҼAD��S�=P�';[E�QC���H�[T	=����8H=��<��z=��<����P�:�0R�<j�c=��q=<�:����<1L����<��j=��<��A�����g�+�����������a�N=��[=��]<qT<2[�<
�T=�o�$ ��K����<�0�<]����d����c\S���4<%���a��<"@�0ie��
=��<��e��S�;Ww'�ŅE;��(���7(��x�5Nt=�	�;(�y�8�u?=���:fL`��	=�W=���<�<�j�����:4��<��l�Y��<�۞<:cw=����*݀���K=�CM��5=
�= �;��r�,� =y���Di=P{=R�=O�3�ms9=��W=��a=��c��K�;_ͼ�� ���=A�=�t�<5e��?��x�<<�b	���
<nO��و����g�-=
Z<����fT�O��:XL*<�K5={�L=Ys���(_���70�<QV=��˼��໰}/�%��@�n<��x�W�6��O����Q=]�E�t�<D)�:_�<�aA= �N<ȏ����μSn��e=s+%�ؚ
<��<�-�<���<�{�=�1g��?z��� =5W5����;�J'<�2|�T�i�Cy.��W�͒E��Jj���༝��<��<6�$=`}��u+<�dI=Qz\���<�%>��~�<4�h=|w=�#��f=YPϼt�<T�8=���3=3Z�<�#�<eJ���n+8��#��j~��e#��_�=��f<9�H=���; ���8�� �۴���=fN�;���<|�4<b�|�UT@�?�n�;�e<l�G<�\�<_g���=���;�(�hJ��R�P�l����'?=P�>;؏���e�J��;�냼�u�S�J�u�q�2<ĲN<�ż�d~Y��5�=���<L�B��]�L�G=��i<00�Sժ<�=?=���9�!��c����p߼d�9=�}��X�<�r⼫�<��*����A�L��� �<�BT=�,O�:�n=P�=��<�6��!2m<�$��	X�޸Q�u.J;p�<"I�<�=�I(=�<:�1/�I_��E2=����5�er= >�l*s�w��<=����Ȝ�<Bu=��&=V�*;��J="��<$0<POS=�n���Y]Լ-5�#'0��1���T��I=��3<��;��1=�����Y4�@?��/=�"-<��=�k\���\<>�!<����<��<�� =Io0�ceW=o�
=m�ǻ}��<�0*���Z� Hu<4�L�W=�n����.=Iʆ���=,r;(��<�n �{��<D^�� V=�n���<8@?��,�<G��<�6����;3�;h�����;U��%�<a%�Op7=*�5;��4��l�<�n2=(���]����<�T���������w��r�<,.�]9]��n�	��<��l��k��>�<9Kļ	jP�~3�<B`=�9k��Rd�� �F ��/?�<u$=�?@=U�<[�A=<�=�m���w�#LG=����|8=���;"`�9"�Z���l��O�=�f=�=�=4=a8;iC�;�`����ͼ�w<�<���冼�|w:4�R�4%�<@�.���:D������ �;I�;�V=	6=?ⅼ��	=�Wi����y�
=kE=�<)ti����<��o��
���R=��]�]�g<��伏5�<5��N��s���y;=?�����=R�	<M�Z=)E=�P�<��ʼ_��<J7=~tH=��]����<!+=�]�<���<Y�e=����/u�;θ�<�^��m�~<S�n<�;�26;!꺼�<�:Uh;J)=��Y����U��<<�<Yx4<Nr<Q%)���<�^R�3�<��<޼�[;E=q��o4=�w�;z9=,՜�h�;�주�e�<��<XW�� ��dɺcE�KN�us%=�v:=
�;N�=��ƹ��x������>��a#.=����I�K�-ݜ<'e=�Qϓ���h=�~ =Ĝn=s�3<N\���B=��?=6�W�4�W��X=�m���r���=��9�'=�2��v���L��\-<��u<z�r�NW���9�zI
=!�x�[�w���̺
�<�t�_�+�v���ԍ=���<U-"=`Mм�ϼ�Y=�>Լ��l=�Nv��R���8v��D&=bd:��^ ���J=sz��;���<H�k��n���wV=Ub�������<8j<��=%^p�RU=�|@�(�h=��<T��<~�ڻ��3����=6=����<Y����P�~�<L~!=L�=ë2���=�x�������R;=H�v�H?=����8�6=���h�\=��<}��<���<�o^=��q<�33�1<=j�1=�p <�j+���/��@��{�<���e����;�9�!��<`' =�Ь��`<�);=X�=���;��+�'z7��]��Rw�<HqB���<^�:}Un<��R�>=2�ռ<����9�Rɻ}��9D��i�o=��⼐�7��)<T�3���L=R�N�rj�o�<��8��#$�C�	���c�� V=� :�0R��B���F�6�ڼRQ��*z�J�k;�L�<�M�b=.��L�8��<!=�K��ԫ<���>�����bc��	� <�<�x�<I8=��;��< �=8	��#Ἃ�k<��;g�$���[��8�aU_��c��m<��<!m]�#�,=�x�<�"=��&=���<JI�< -��'���B�o�Q��_� ��� ��<ӽ ���=�W=2�]={���e=Kis��`r=̮(�����b$��+P��׻��P�#Br<�<3=jİ�^�=�CL=Ϥ�<|$���$@��,��+=a�ͼ��D���[���=���SU>���#=9��<�3S<��D�y�a<m�	�zK��^�<�N=�&=k?�*���j�U=ح��p$r:�4�;�G<��;��7=|R�<����N �\�=ʼL��<��'�=�v�k��<�8�A��=�tZ<{�=Q�U<�u�;�5=�_�RJ=�< �Q����k�(h7��:=1��cZ=��%�]fX;4X��`<�+�;,�<��<�\��=�3=w��b!^=M��|zq���<F��<ߢ�<��=Eѻk�7���d=��<�5���`�I���=��	�;ln�!��<'M�NDm�t�<�ț��-=�`����<w���i=��V��Ǽ�m}�=�>=/<=��<u���',=��<��<�,=K2ۻ`M=Ԛ�;Y�e=�&=!�=���<-��<����W=�m<=��;�@����0�<�?���-��+<`�� �ϼmC=b��U��<[�Ƽ}���>��2�=Z��<3a=���<&mF��ȋ<Ù��u=�[.�ߢ�;�����?q��<,=�ː��,=P�����<�.
�b	=޿��;
;#�Q=v9��]�<H�����f���~=��<�l0=�y-�S@�<N'�;�=�ȡ;35=n�S=�y�P��24t=�2=�;"��  	�r�:=^R�<z~<�1�<K����g=�-%=j=�N=���i'=r���S�ü�,=�9+=��p������w<]�
=7�R��3,��S�;���<�,�C`
=]�L�9=(*A��N�W�q<[W =����l��쭇<b�<���:���<��ͼ�N�<�"F�Ա =��=|=��;�мH*ݼ�5�<��R�v�9��|!�G7���*�!�@�_+m=��ɼz�<�l�;��<Sg���=�l�KP�<�K��F�;�!��K1��ӻ�S8���4=�H�����C9
��Q�<����.<z|ƼX�*=/���x=�n.=�P]=t9�<s�s<%0L=d�z=F�X:�)=���<�����N�̼B�U=��l��U�<�V�<������u=���\8F����<�w��Ǎ�=�|ܻ�w��_
<�KQ��x��d0�<|�?����;>]���6���+&=ۙ��O�=3e�G�d��:�;1��;�����<9I�?���^�Լ��d��G=�=�5�	K���!J���=H��=q����-;�t�3�X="	�[�j<�`��%>=������=��p����<�QH=d�B�M#=��F=�>���/�s����=�E=���}q����_���NS<$i=�C�Y=�����8���&C�ӻ���9ΰ��oV=
m�;w��<vl<�5�X2���<�`y�q�?=��<�����<��N=e��LB���<V�5����Tϔ<�,�;ȸŻ�G�<�.=t�;|�;=��<�<�D<1��8=�~0�m�<��W=O�:K��<�v�<oA��O���an�{�2�'����8<��<T�Z�����{�!����&<�b<D�#=M�[傻�K=�C=��Z=�,�4���c �B��<��4=S�.=����V1�<e(u������=�\/�M���{��XG=m	o<��f=��;���z��<HbA�S	=$�T��CK�����@<.�=�Y���q����P[�rCF�Wٗ<�0��x߻t=!��0����h ;2�����<�>0�2;p-8=��.=����GC<��=���ͼ~]
��O�#q��T����<�1<b4�B���q��^�l<�[�,j=�R`=�(@;(�<3l�<~U	9D�[����<D�z��X�
_��D~Y=�Q)��]�J�[<�3�<�U=t�ǼI'=<�6�;H�F=솫<v4����Q=���r8&��92��{�tBu<�d�<�"F��;�:9V���h�o���4O�l��<�.=�d�"�T=4�V=*H�<xO���ҿ��Q�<s� ��|`=��ػB��<r<5�&h��B�=[�=}=�<	��<��;Buv��Ǥ���}=T�d�Fha=�j<�T<)�=�V�<ϥܼ��E=�袼��8=��>=Z�4�wGj<YU=��<�k�F��<V׾��r<gͻ�W<�>��� =�Y<1�=�L�9i�=�L�<=�:�����?����K�+�Żt1<��м�g=�<���������'=�t<1��fN�;�=w��%�<K;)=�u.=M�X�1g�<b�;�DF�<�z=��=(�\:�=�57<�==S�5�s��B��#}�W�U��?V�ZW>=o�=S^=�V=��8���<AR<�<����T;�<�O4=����X�����;o(���ļ�J=��-=���;	୼WV@��~�;q� =b��:��'�����S��@,���K��==p��<��)=��E�oL��jT�'듻��<9,�qI��$=՞=��<Ԝ���P��:��D�<�#=/LԼ��8=ǟ����ȻTJ:=�O�<���<� F=F0��z�<g�<ga�J@��V]�ea7��<ޟ�;g�<��"�{����3���a�_�Z�m2�<� ��\a�������T�<�0=-<Lz�J��<��� k=pR����!�O=HK=#8s= �������7����I![=�� �x<�����+�T�z�Ӽc]<Eh<�8�;��=��ȼЯ�=�ګ;W�%=\m���$=.�Y�]�X<9�J=K
�;] �:������=���<Q6#�vr�<�L#=Á��i	!�<����+��P�<���<���<�c�<��˼	6:;���<Ut�<3D6=�3=Y=���<���]�V�"�:�C��ˤ#={�<v�����=��@�?򼖚=� .=n�R=R0;.[=� ;��;=�Y��rjx=�:T;��c<�)�X�T��3�p�<�=�� =�*>=�2n= �p=�C:��h�m�d<+u�<�3;?����r�W��<�7=Iq(=���<���l�1�5!]���S=����3W�;�ކ;�ti�|�e�I�L=�7D<��I���F��M�{�`�a��<�h��Hl<���<�@{��|�ɢ3=��u��G��RU3�ݖ����K�9o><v=�p�<��<��G<��	���;f�=}�2<R�a��<�,����<
�lT/�ԅ�T=K!"=�	޼ �<v�<)/h<�2<F�4<wFl=Q�<�⏻��=����)=r��T=@����	�<l�L<n[���k=��B��.
=��{�X2F<N�e=`�=��O=�]G�2��<*�-�9 7={�C=�l�O}n=XT�<3Z��<m3� �x���\��&���ҼP��� � 
�<@�Q=��(=V�����j��<��Ŵ�<y`���(�"�Ȁ3=�8�<�Ҋ=o�$=��Z��?=H撼`�=�I�;�0���ʼ�|��� �+�����H��7ϼaC�-�
��6='T�<� -<�Ē��j!�CG7���(���(��,=D���N2�uE／⨼�����S�7�n�`<�Z�=l��<⥉=�^.=`B��d��L�<G���g/=��f<�Ț��
���k�(+�3-:�y��<�a'��Ԗ�7���73�N[a��s(�����<~�[]~�c�R=��t��$<k��F���9=���7
���`=ݰ��Ψ= <�:.�I�Q�,��<0>=�@�:�m^��7�<U�=��]=�B?=A=[�&=��<�a:�v^=/�h<���<G�z;�����j�ќ<q>0=3�I��c<Pg=?d3=�k~<�9�<��!����e�m�� �<;u��C=��1��_R�������o�>k';�Ӥ<T
=����'7Y���<�F�<4�ϼj.K<ߍ<uJ�����<Y�5<��;Ô=<*��d�<C�<��=g�T<��޼dȓ;�F� �#��k�v��<fi:<�ٹ<��鼬X�<k�w=�4���m��k=�����>"N�ؕ<%�d�<�;s�>���l�<����=�]=�x=�oW�j�N��B/����<9c���%�;��FP��� = =�lK=ޤ|�K 4=YU��]mQ=t�D���,�\/o<�@=�)�[�8&=5���`�4��<S=�3�p������.�9�hE�����%\�j��N�==��=-
6�!�;`�A=ۮʼ�[�q�u;7� <��=�|/���!���ɼ�/�;G�u<	)��֔���發)iD��k�<֒��}�=ps��=s��<^�Ҽ7��<�������N�<����I=k���l���h�<�Xp��
߼�SD�Md=2���=�V=ې�<�vJ=��F�:<D�ü�c�<��ټ�s�#�к�Y��M�<���<��y<��<�=V=���bT;��<1�����(=V� =+��),Q��uڼ>����̼��U�zO���
��oj��!>Z�h��<����I*=�j�<�&:<x����,=6�@�#�O=��<��f�]��=��;���;�N+=�.��d����I�(W���;�
��<�q=��C�|G;w�J='�i��L�{f��0<�?���`c�&�d��,��f��>8=�p`�o;7;�򀽰�J=��<�@�WAӻ\�ɼ�kI<�G�H&ܼ���;Ork=��$��SF=rf�gF߻c	Y=�L=\Im={��<��{=�:�j<��5;rDF<nyY� �R=�)=i���
�A=\�:=ǌ���#:��t<u<��v<�:ż:y<��=�+E�Cr�䍍�y3��"�U<�aW=����nZ��`.|�4#=�Y =�H(=�(=pl"����%�g=��,�j	�<�M�;�\Q=q�<"<�)Ƽ��V��i�3tu�_x
=4=���*o�;*jH=m��KsҼR,:1z�<��y�F:���I�=PN�1�q�T�)���=��;/j�O���gYS�i�j�8��8=�D&��Y<��i<WV=� <��a=�2X��!<L�¼s��= Ӭ���Y<���;�e;�U�<��:�G8��\��tN=hӼ*�����<�Y�s��b����/��pڻv���B=`��QԈ=�G\=\@=��߻ēC<�)<X��<M�<���Zo9��XB=��>=?��<�o=�5=� =�l=��9;�Qc�"'Ҽ����#+;N���Dl]=lF��+<CRX�mR����8��*�'Ԓ<��G=�e!�n=x=��=��-�q�����R���<%��~P�;"�ƽ<=��T�Z�<�6=���;OT?=ă���c���߻��=����%�<��w�r/,=�_l=�=�<A�T=���;�<2ڻq)=��2;��<,�|=���<�9��*=�Zf��h=�ݡ̻��X�S�Z��`&=�}��If�;|�=*<=�;Y�[cd=��U=aR=��Kri���?���<���[=;m�<��o�}ᠼ[Y;i�����A!��m�<�l<�=��;�s=�N�s����;��^���!=��Gz�=S'�;^j���F���<±}�3��<mhi��ˋ��a�� ��6�<)�<T�=5yV<]q.�Ĉn:�|i����<�US;�%h;��Ի�u¼0��<�6�������<ˀS=N�`�V�$=���<��/�T�<���%�U��<��z�L�м�л}|:�7,1=��'����<T���b<:�6�H>l=Z�,���*�F�"��E�h_M=H��<T�<@꼊-N�3��oG=Ǳ��ST;�Q
��*���1=�Ag����8"����<V�Fhk�R�;}���b��Ի�=lY�����<y"����Q�!��OI<�ӝ;19W����;�L�=y�ټ��<��<uA�<�`�=����4��!=jBH�3G�<���<� ��x���g��Ђ�2�=6�����]�ÿ�zg�<�n���;6%?=��;H������i�#b���bP=���<#��8��|��Bp��h9=�k���F�f\ �.��đ|�䟿��q�<����$�<�a��T=3O*���y<��3�X=��7<�5�;�U=�xH�=�l]=Wi�;�K=2��<�=�@=l�b=dc=�r��Y$�0~�<��<�F	��u �������<Y�@=<��<K�ּ��=�5���M���M��z=��<��M���<55;=��3=���<��Q=�PT=��<A|��UO8�P��<'Z�<ң=qX<���;@��;��)��ui��K:��3��J<&� �;��<:R�<�L~��H2<���d�#��*<�L={�/��T���<�?�<��_���ի�<��;=k�=d�#=�&I=w{�<|�J=?�e���:^�y<֔ ��f"�$��3Ҋ�5����D<�V=u_�<֮h��AT<���tЕ<s!��27�����;`�����{x�֛��J9K=���;�ʼN"[���ּ,�"=�2�o5��*j�b���m�-+=Oe�<[4<=B@<�&���@���X=���<�;;�`���]<>@�G���Kκ���}�M�K�	�96[�;�<�F�8(�<����� U�Y9���.�f3)=�~�<�=ϒ��n�?��/ <7�
=�	���UL�1^=��;�=�<�͋����2����<X����[=/A�=�ҟ��QW<�'�s?���a=�6F���!+��q��]�:IM3��'v���}=�j<-5��c��4A�:�{=�MR��9�>��F��=�5/�;�	��߯��G.<�H^;]-�<����S�z�PЛ��Ӈ;�晼t಼��]=�-l�R���.i��3|�<�9�<�9=��j��D�;�a �S���h�*=�C=) ���U��:�:qz�<����)r�����p�<iޭ�W��<�ת<�޻�@<��<��.���=�:�<.yc=��<�vҹb�E�{[�@i��3$=f=�_V=x�g<�dԼ�q=@��Q<��јĻނJ=��#=fo=��H<>�b=ۻ�=?_=�+=�&l�(�<O���;S<� =���=�3�;�y=:Ȫ<Y��<��:;b�0���L;3 <���<k�:r�7<���t
=T2K�O0\��CR��P<w��=�1㼒��<�M8�w=����:�|t=���_��s��;��P��,��z��<��"���=c�:��o��[;�:=%�����S�1}��I,N=��T=�U=4��2#=�0ʼ�&�������e�x�N��I=)�ڼ58=Ѝ[<�)=�����*��Z�~�<��E�����+.=�3�Q�d�I���Q=J��<t`�s�t=0�<v�v<|ْ�.�Q��MB=l�{1�Q��:�=�ؑ����:k�9�{�5=�SH�q�B='���~��,��<S�X��<�5�<�M4���һ�Y=�9��b��
��N�W��*��m�<m�8= B</ż�]B��da�rn���;ڗ0�d3�<���<���<��	=2�}=�]�i�M�1�e=�`"=�o�<�ݸ�ں���;&���s�<`T��?<�����y�+��<?��Ђغ�⫼єu�ۍ��$�)�b_d�s� �:1+�IY<{�G=YC�Pȼ{-@�f�<�ϴ<��<=����tl���J=��<
e=�ޠ;�t<�d���V=��:=]O���cm=P;�:,�<�qa<��鼏nT=�Wa<�0b�Ѩ�o�<�p�<��1�d"�0'�W3_;��_;9�<�D=t5ּx��;K*��J��b'��#���k����;�"�;\��\^=A�ϻп8����� ��<�蘼bP�<��b=�~�<oJ]=��(�.!�l�K���DC��i3�(���G�.��üclO=W����:=B���zEx=v�,=`���?��P����� �<�=�e�=LX�.�#��Z<�"����<`b����:=J�_=��#=h$����=jN(�0E��(��"~&�x�����(=��<S�M��dJ���<\�K�ar= ��<��X�ۆ����R� �2�|�n��/�<-���Qo�hAؼ�s�kā;CL9��̼���W%���<�#�<s�=Me�2EM�_$=��;�u�ש��=N�=���:)~ּ-�9�?Ҍ<��<E���b��k< =iES=�'=$ '=>=�{F=��
=�)�;:+t���û�-��4R	�K�h=�Ｃ��=8":U�<�r������������i=���<ɯ��k{���F=Y��ZB�H��<�9�;�'<�� =dLb=��N<ʴ�OU; �f�*���]�v9/�`�R�YR=�A�<��!�b�u=cI���)���A=Z\=M&���(�F�<��ژ=�n=Sŏ��w��WI<,ü��<�5��K8�,�����9,�>Il��s=��'���'��==0���9��:�K,��L=��W=�Wp��fU<�䈸l�Y�X_ =��;Q����]}<?�ۻ� �<V�d��[=�{g��Y�<D�n=�?�<Kñ��ּ��<��=h�=��ݼ����:0�<O��x=�B�%��v]�<���<�(7=�<�����#�6]��IT=s��<b��<<�j����<<k`=�|�;��i��!%=g���*���ZS;Ǿ[=de���E=��<-�Ҽp�#=(:�<��+���%��\0=<=�x߼�~�Z��<���:]�<�g�� �q�|A*���H=���;*��;���<��N�j4���;�lj.�W�~=)`��!<�;�<QN:=�� �(�/�ʎ;����j=���<.<9�sYe����摴�������;3x��C�q��S��K4=�<ռ��ݼ��V=��<���RR�\E�<�T>�`�����v;)$r�&a��#D=V=��T=���<H==�Ge�Z��:
3=��ɼ�U�U�ݼj���C�<��c;���;5k�<*�̺�mA=�1=i+�aS =?E=�L��B1�W0=��!=��U<�����=s��=�n�ƿO=x[����?=�i��x�<���<���O���@�?�ؼ��?�t�]<�����g=�ૼ���N[^=�<̚�<��*��=�f=���<��.�e.Ǽ`rc����K�6%�<àm�؊���<��?�s��<?�'=O��}O��Y��N�;���;Vl�v�<1o��>��rT=���-�OD1���м\�(<7�,<DfI�$�=�j!;�]M=)�����g=���:I�7=+�n=?�c=��^�gف<�e= �"���?�>T�<���<���<3g<uӳ<��μ9k=���?%�<����t��0���{��1<h�&=]�:D8�<��=ǃ�;�^,����H4<��'�E6B��C�;+�<i���9=��;�-K���<o�<�E�d��<��G<�r�<V6ּ���d����b�t�b=i׼ɪ>=�.d;
�Ⱥc�?��j���Ӽ��N=o��;/��t<~w=��d=!��<�᩼��z�7~P<�=�!=D#I�O��;��<?����ʹ;6�=1{5=��0=hVs�o>��f�:��D=�bB=|��<��#�g,�<�3F�3=�E]�>����@=�,�<����Ne�
�;�2�<��˼���̼#����<;�ۼ�ۻ�;-;���Lp<�>=R�0�#w�<A�(�����2��$���<�^r=y�E���=�iG=]��#�m�2='�#=��N�fo�%�~<�p<�������c����� <9�<� �z�����^�G��6�[=�-=��YP5��a=2X2��[-=���� 	=,z;�������� ���%�d���f»+�O��o����5=ؠ�:�G#=��D;�.m�r����XV����B ��x=�o=;��=~=7�����A�X�����)���
z:��=�:<v䐼Ĩ7�˟Y��8�<1�,=�-=����Ի�*;�����V�S��}̼�=��%�
\=�t=x����;�;R=w_=>�*=s�e=7=-�;�w�/��Kl="-��JT%=[�=������y=�T�;��6=f<��<�Lp����B9<?�4��7�L�q�>� =����ş�;�'h�Qv<�26�Ɣx���h���=�0[<*t=j�Y��A�W��5<=I��� :Q�a�a�^��v=̓*=��:��󼭜�;�Ҽ���g��5?=s�)=gG��"����b�=:�e�c.m�>�=�*����j�׼���<��
���*=�&��������&=h�~�'O=T�-��B��)��OXR��ֈ��ռR�ϼ8B=�ք�>cZ<:��6Gk=��<.n���}7��p�J�������{�;f[��GJ�Ni�<���<m/�;~��<���뻓�R=Ev�<#�=<t�I<6A����;�{B��$=&:1��<�H��I@=��J�g
�x�J�"%f;��!=Gė��%I=I��<@B=}�e�IÍ����<c��#茼�$7= `V=��/;2�`�/�=����>�0�W�j�(�AZ�zm:=YX�<�,�<�/�<HS��'(w���Ǽ~,м-z"��pB���Ӽ`^�>^<W��=0���̷<�B��Fi���<��<Pt�;1���e��?�E=RR:7�/<��<l1=�A^<��=� $���D�4�]�MH�V�=A�E=� =�3��E��_=�[�<�Բ<�u^�<��b<�)仚'�;��	=x\��LK<l�~9�q�<F�J|�<����Q|<5�#�@�V=b�ͼQo�<��Ӽl���c`;�����<x�;=�L�q=<�y�<a�E=�m�C��=8�3<U�Q<���kk�p�"<l�<~�=t��<zS��6 �<W2�<yD'=E��<��>���,=䫼<�6�Np<i4=G{R= �\�r�)��==򮽖@*=9�7�4@)�[� <6e6��O���<��
=��H��ȩ�C�`�dE���x���%<�g$=xg;�6���o�4<�ƈ���>��#Y=e�E=ć��]4=彍<����oH��\�<IĎ��j���ȕ<�V���j���6�b�����5J>=��ʼ�VR��_r=kL=�*���Ƙ<{>�����HW�<�≼�5޼?!��㍃��K|<��l=I�"=�mf=3���!˼�ZA�ӱJ=�v��:����D��W;R=߸��E�O;=M�<�$^=�q�<@T����R=)p�YD�<��=� �K���Z��a�ˣ����4=� =D�<jPռ'/�:�On��f=3L6=�r=FU(=��ü��Z=��c=����]�/=�b?<��Q=Õ=�G!=Ѡ�<`��;�P;��W=��M��3`�������<LU=����j1=����ӼH��=�f�6��<,�$�h��[|=�^�<���|L=��<�+P=k��;�s��]};�kow<Re�<�3)�y��b¼�����U�J<&�B�2u��9=x�ܼ�?���=�A�;d����|�.�#�O6=iߜ�������'8�<�~<k�==���j���i���_=�E<��3�߻ļ޿�<N���Ъ�o�=";���d;��%��U�;b�y<it[=���;@1����<	j=N��;��� �*�ɚ�:�I	���=����?��
�}<�"=��<}պL�h=�r�k��5�+=�=<�%�qZ=�J=�����i_�C:���#=�l��m?k�0i=7�3=>
)�I��#d=��<L��%3=�
&<�z,�R�|�����Vƻ%'s;P�Ȼ��=K5���<Jb<�qn;yߛ���-�$�k���-=��(�o�`���X����5e��#���<AU�:�ڼLC���N�<qT����V�N:�6�<w�q�(U�<2=��^=_ݜ�n�=�g�� �����ͻ�⹻�ɼ��<�D=|�ﺮ��;N,(����;e\��<�%b�-�X�<�K���>=,Ǽ�׋<m�Q��<�Р<�Q��g�:m��B6����������u�<(�*<��h<�l=e�&� �����r��.+��Ѯ�WO�<%�Ȓ/=�z<�<��|��BV:=b�����\3��#�L=�M<dq�8��p=�E<�ږ�0�<���k ���x=��케�=jH=�Ƽ�!=�&�����b=''��.��M!=�;�/\�<z���'�!}����d���S��'��;B���i��<�����c<>���\�s����c����8=��w�%ro=+�=�Co�.=��j��ň<��~�	��B�A������S�T[ �� �<pg<�t�;�U=��=���;�6���<W�#�Z10�cQC��%�<����:#��{q�E�`��+=<Z�=���V�<�T�P;/��2gz=ɝ���L>�./�Sw����<=߬9=�yv=���ּ���;iH����<
0=�l�:NH�{��;u>\�E`���i=V�8��䒼�N%=c��<�+��
ռ<?���*S=輆�D����%��v��I�c=E8=�y�<��=����?=�(=\U<~��<ȶk�����h@&<�F�;q?&=ʴ�a"c< �a=��:�s�<�6=�1��h���=we ��N<ٸ����;q =��C=~�ȼ(�����}���;��;I@���)v�+G+<���J<6HD���O*=#�ϻ:t)=DZ�<�XC;T�A;�v�<=��<��W��,=w��<6電��#�Y(I=��&�̊S<�]K����=�1�Q��9G>;=�;=m��^u��I=-��<�g��	⇽7����<��<w�<�$=Dbz=C�B��8�-Zo�w��Cq��/3=r|�;8�r=����l]�=�%�: R����<a3^���d=��(d�<L�<78$�rx���ȼ��J=4o����h���=����b�\��P=O�`�Dl���e��U��M��j7��Jۼ�<=b9!=�r+����C�><�u=�c=Y�=7��<��+=/�*��=ә
=��%�]���H��:�s=@��R �<n5=��,=�*:��ܰ<�J;�n�J=3�6��9���?O=�����:��f==ϒ��'V.�p�"ݼ��k�y�y���2=������*�����x�GVp���<K������=t����d=Di�9-�<��<�T�=M��K����n�<�+���#�	%�<�J=f<%~���&=�� =Tȍ��o;���<��<��Ck =z#��z��=p�<V����?��5J=H�=��Z=���=|���Ќ<����Kl<��%���<�Z=�4=qA��g�<�7=�˟;CN�<��P��2�8l	�FV���,=\�A;X��B��rK<|�=$JY=�ς�U��;���<���<Vu=W�=kH,;=L��]<E����d<o)[����==����C��Y��LM =���}-=A%P�s��<)N��/=���<���;]�ۼ� X=C�<�-U߼wq*�å�<u��g�i=��T���=�E������`�����Z�<��r�m��(�g=��<���	缧d�:r]%=�@��ݶ<l�p<���<=%=�,��O�:�C໊��<]�����;
M:��+<a�T�'��d;�ܐ���:��/<���<�Y=��=��=<)��.�<��;j������N�ͻ��X���=�zY�3��M�L=�\�0����I��(c�$7�On$�����5<��޼S�~�{��+><�(:<2����B��d2�3�?<��C=�S=ei��OF�<��|<e�»�IT���$=2���9�<�])��,e��)ʼɽT��!�c=pWJ=�A<T"=�`Z;���:p@"���F=j/B;�5�<
��B��:e̼G�=ֳ�=g�<��<�;�<�V�<��=�ɘ<+�<dΆ<���< �L=<R�������7���O=y��;!7�;�Ũ�Њ=�Q���d��<�ü䐽!3:=C �*��Y�<��=s�0���]=�G��3�:낼�"C��i���6���r=Ӯ�<z�@=�E�;�����#���T�曓<$�2=�#�F�<=���_k�~v�=tE��%Y|<%��=B�<�*%���8=+ҧ���=��ļ��R=G�<9��NBW=���V=�c�K�<���xl��R��ae=�����5��O7<��g�y�'�%�C=�=`#0<c�X=�;=!Ր;ub��ZD���+<B��<��,�i[=[v�p�7=�}߼^I �>��:��*=���C�q9���=�=W��;�h�<�/ƻ}Z���,=�o��=��X=I�<�}��.�����<�hS�&w���<ݲ���{<N��g�&�/z\�?�<��X�M�;�;Tro<�>u="�I��Mʻ �;��<��=�"=2������4�;$�E=#��ĊR���<��U�C+;5��t�=Z< =�(2=�={Ć��F�=�f=ϟo;J7<�zx=-�����N��
=��!=q��<�{��$�a�[�U���@=^Ʃ�_�R�z ۼ(��<�d�;l������E�`=s�=}�P=���<�M=�]=-9=-�b���X������Bϼ$��OM=�=�<���ɻ�񓽅5<q�=u;=`��;w1���;����;�<��<-&�<�uA�: 4�>9�������<�~�<����|=�g%���q��wU=X�_�d/�<MT�<�I�;έ����<G<F�;�F����;E��<�L=N��<�--<B�6<"Z=���<@� ��[C=�=Ty��\�����37%<��:�' ��9)���G� �< ����Ƽ.6�3�������=��!�'u�������b��by�� ��u����K;\<�h缇�<6=.��;��A����;��W=Ȫ�<IZK��o<+�x<�uA;$r���=*�=&v	�v1A=^��<q���<y���`�r`��� �<�6=_I
�Άr��UF;uCt=:�.=4���ߺ��m�=����t��j�Wb6;n��<w{=���L|=���<��#�U�s=��<gU��Y �����
�<k
�<���,H�;�3�7RX�LG*=�NL=�zݼ�Mx��fh=t=�Zq;_�)�=)󻮓���/�<l+=��S=j�s=C�=�E:%����jS���`��&�lB˼�4��m�_=�bO�a���j��<��=N�,<=�I��P=��<
b���<��<=��5���<�n$���F��7]=JiM�V�<~W��A��y=X? =ǶZ<��<mL��w=�R=��<5�T�O�y=���<kh���h<��@=�!5�����#;���=i; �<E
=!�F��C<��9���v<���S �9I�{��mA'=m;<���� ���� o�xLr�LH�g�(��P=�2=��� ��ͧ�x��/�	=���Fqѻ.*�� ���Y�<+�F=�n/=�OD=�W���-P� e=�JL���*=�4��jb=a��<�qn<�D~<�_��@S=�9Z=�}[��4ȼ�=6uڼО^����<a#⼮KM����2=���;1�2���= {�<��<�i)=9J��~����_�?/�<Ș����_<����%=(K�;���'� Ɛ��"�v_X����;)�;.�~:A¼��4=�)=�;P�%��6U���1=&�^=���<��8�� �	M=8�ܻ���:�3f=�o���;�FT<c�6�6f	=H�����=G�=d�D�;��<�I=�9+=}R����O=J��<���2m=�=1�k=��<B[�<a�'�"?���ü�¼l'�j��i�2���=2�*��N[�QQ�(�����<��ȼ�z=��<è���-=㈽�逽�o��=,���j�<���;@y���l=Ɯ �h{�<0ۜ��'ܼOm=̖�s�s=��)=3o=��;����X�u����-���0=�>(��=
���.�=�*'<I�n��6�<X�k=(�<K��<�ͼb�N<>,d<\@�<��=�z%�l����g�T1><�񂼥�C=��!<3�=�~���z
=g��:+��Y[���_��m��H����",<>��Qw=>�L;��˼?z�����t�(0�<©$��ޅ=q/D=��'=����av�<�dz=@��;��<�%=��;�1-�>�b���s��p*<�̆�%�<V�K<~�;�#V<=G����L=���=��=0�h�k�+=�b��s���|?=[C<a5��+T=�I;�/��
�&=���<�|�<<��<�(C<��=��4=��[=K <>N�Y(ܻ�<�H@���<{D��u=� *=A{a�o�=�K2��SZ=���-��m�1=���<"eS=O�=&����=SS�=`0f�yW+=��=��Ӽ\����o���,��;�:��<�;ɢ��;Q.=fx�<��=	�<���G�9=>��<ɛ��!���M=��ɻ�)<�i1=yH=臺����<ܛ�nr��fA���;�8��{��<�=��=���]�z��;3m-�Z4=�<s;=	6<��B=x9=0;���	<�G��ü����W !=�������x�M�)�K��=Z�	��*��v� =G� �a�W��zz<��
�� '���)��<���<Ϛ<L3󼽭�<H�%=�E'=�%�:���
7o=i;Pż����ď�R�i<�*A��D��i�<�7[�� 
��k����N�pѼ��@<p퍽٩���hO�����^.�d�A����<(�<9X��1=p�H��v�;c�<I� ��<U�1qH=�����<��~�u��<n"漳01�<��:.1��W�$�fӔ�)9m���8�.�+=5=��8-�<�j"=��B��C=gu/��A=�9�w�<_��~I��,=�;��
<f9�<
��;��v=�4u=?ɰ<z�
=���`֧������W��0J=r=3<�u=��é��Gi�b^]��~���ͯ�B%D=�A=_!r��i<���;�m� �<.ލ�"�h=��J��I�)��:�A4=Lc�<�f�9S;;����9=���<aI�Q-y;�9="�:��{�� ��D=w����<ޙs<׼e�� <��&=���<�S�9PMr�F@b�ƌ�;K��<|aL<֎�<�<���<Y���J�^=v�L�q(::�<9HJ=+O�4�b�����@B�����*�h���h�<¿C;��'�j�l��R=I�f=x% ���;���>	���μO����]�c��+�K�ܼ����J��<,�,�|C=�	�D�<��=�L=6�p<�D��!=;f!=f?�����=Y+<����fK=�72=����V�ƹ0����T�OK ��1<�@�<���<w]�X'ۼI�<��F�71��=�I=�_�e�|�q���L5F�^@@�	��;�Km�Du1�ې�<�	p=���<�uK=�Ч<7�.=�D=�FM=�L��h��;T<���)��1����o����o�<v��<w�#��w�;�����L=���[�=a���k��:�`=K6�8�+�;a�c���<E�<�h����̹l �c� =�g4<Ԁ�<��j=�9~=��]�ľj�tI<�7���lD<Y��= �<HHH<�?���&�=RJ�;o(�l��?��P<�ʆ�?�<��ؼ5.��g��; +=GE���v����Ӆ=/���� ���׻(n�<�5D��)�;�S=r��f�)�
�I����������E=������N=�<�x!���=ʍ<=`5	=��缇�=գ��:��sJ�~/%<���<����B�=�H�0�?n�:Okc=�S�=��������A5�#͑<t�o�3�żS�ͼ����4;٥ɻ7pI�����@�q-=/Q-=!D=(,=�:�;�G�>�绮m�ˎ3��jP�u�'=B�ֺb*f<�h�=����R5�;�9%���.=̟h=���9�8��)�<�Dc��r8=bsA=s��F�<k�j=\/<i��:w�=���wV��{�;~{����b=��<mqE=�
��_d�)_I�I�"��/�C=k9��=C���u�<�s��*�<����T=�mJ<�O��P�;�A�<.�{��P{���x+=|�:��LƼ��h=<���Z��<N�����3=o�u=��<N�,=� �<���<��-��v�<���Y�=i�n���=�}��,-���\��A�\��<�5ǼdD=�]1=���5�$�<Q廼�T�by<�]=�;�3�̼C�0<�=OID<��9=� �;�ļ��
�>9��e&<����=%ּU#<�g>�e7��咔�iW�<Ul=��V<b<�e�:��$��ɼ��q<�b7=4`=q��=�u���#����<���<>#Y����uH���4��A�<�<S=�B=�����6�Y�׼�~ѻ���<�t���k���w9=����=WlѼ�I_�젼�Z =,�;"����K9=�\H�p(a�2H��]"=�P=��=0��<�!�Ȥܺ8Ș�KI����=h��J��*祿��>�*���fd<C3��5�:2빻e?�<�����4��<,L=���<?��9RJ�S��<�w=s�;���;9�+iҼ��f�1���2Ҽ*-�<7Z3��<v��&�����ļ��)<�E��\v�
�<7巹�U=�mż�f;E=����:��6۪<U�;J.����<���<;�<m����nP�(�.�>�A=p� <��0=��<P�ּ�<�Q���@��v=7 ��<v$F=��<S=�
�<������X��]2�ɼ=��q�x~��,G=xV�<�d���<DZ=��������=e��<�[=g�����h����%�<���$1�Z�Ӽv{d�HN�A�	�=�j�6�T�� ¼�~���5�\�$=1�4������G<��=�6�J�<ﲍ����<$��;�K:<�<M]'��)�j�e�gh=� ��{�<qc������'�c�&��<�bR��?=��=	�<���:p��<Dj=���<�m=�=�聼8W2��=�|/�c���`1��Z=�b=�؁�*�=�������;s���E�<��ݻ���9Pt=��i=?��;���<�t�< �:����q�<��@�DQ�<�=����U����;��^<��'��F�<{�ȼDM�<s^¼z��S*V=)ks�ZP�<wb.����<i}�<��<=??Q�,$j��?7=z'�;���0�g�j=J]<�,,�,=`D�;#��:^�=?+O=��+�6<��!Y=�l<3N=	z뼥�E=F<[P='��<�v�z���W�<3�;$"!��~B��V�<L���0bG��e��dq:Ϭ ���<�D=H.���a��[U�<���<��O<��{NM�q�,=�=�Ǵ<ki<���=�6�<�x�<����Mֺw�.�3<\=�B����<�༱PS�eP��2��<�&3<M��<�D=:�T<�=\_�;~i;�'=Tˠ<�A�5"�<�	��j�<�:�%:=nVv�#�`=��=-#<B�K=�U���1�ژ<�fm<�?4���ּ���<TK�ɺ�?.<�
��U}/��v<[e�<Ɠ��񹻡��<�R���@�_ӑ���=z��<�8�ג�<��b�v�;�b��
���WƼ�B���J=����0���F��9�{ZU��;k<҅-�I��;A"=�-<8=���<���;'�O����O��5a>=� ��<�#U��+��7��դ�3�=a*<�S�'����Ǽ�/���*G'=��`��c̻N�"�/�M��x��xl=�^R��|T��� �ށ=�L1=�]�-�<}`�
�	�o?�����𼓦�;�)�<x="�N= (ܼ�=(���WO�<��ܻ,>=�T=�-K=-�k�<ہQ=���;Ծ=Q3��!�Z#��*�=�ǹMWӼm{<U.��V1��[���"�G��<���<��=�!�R̆�>�:ż`���f=w��$�=Rj�<	�@
=2�<��T=�k!=ʴ=8P0<�;w�=� �����$X=M�Ἦx���o����<��+��aϻ�|C;��%�Fy�<Z��;���f*�;>dջZeU�H��;t�;���==l:j���������@=�;lʓ<C�P�]���2X���_��Zq
�*G=�Mu=(�*�U����<�(<7�;S�w��l$=�a�<�
� ���4z��	D�e����G=� = ��}N"�Z�x=c�(=��ü
~ =�躩(���9	���}��%�<F�;a����;��<�Kh���2=��k�'=��<[?�;3�E<�	������#D�߃���4=Y�R=4|�
}��xT<�A�<A�
=}O�Ѯ<g�����`��v}�ܥ�<�22<�_O�ȩJ���ռ5vؼ%q=~�+<�iE�BK�<�!<��`=7ؠ��+�;��;����D;�7�;H��=P�>��a��>O<]S>�@]��4�l<x�G��W=��$��ˠ<�*���<��G����&<p&�<<7+�i T=�{==�%=%��wY���
3=^'���$N=��;o�<�$"����=)�y��:�����`=L�ތ=��q���;=��?�!�s���\�BE��"=␐<��F=sP�<~�΃�L�+= K�<v�=`N���w<N2=c�,�;�?�6gn=���<��n<��3=H%�ٻU=�Ȣ=4N�=ڳ��=�"��H�==n�w=�"R=�ԁ=����KɼL�=!去�"=$�=�e������K)�9_/�(X�D/�vK�=꼐
{���=��$���=W?C=���<�Ӗ<�@Ҽ�2<"nQ��7�q�:w�<�%a��|H��$�g���D�==p\"� 8=�e��6c���*�v(��.Ｕ�$�ş5=�k�;4q��=iY=�8�<����;�M=�ü�L�:Y�=�K�&��# ���<W��<��L=��=7ű��K<�Q�<�p���;�����O<f+r=׀�;MZ=�9Q���=�˃�:,6�~�a���y<{$͹�q�&�0�WkB�WZY=�i=�:��K$=:�
ƻ�[Z;~&8�%�����
�̣=�\����y�/����zL����u�ڼ+=y`��ܯE=��p�1ȸ<еȼC6=#��<��!=�n��jM���
^���4=XiƼ��H=1#=�n���L?�u�<���<� �+�7�ֹ�����qq��s|<�b꼄�
=3��<��ڼ�O���<O�<���T9G����E�P=��<�)�=�Ϭ<~(��X�� #=j	1=ڛF=��=�껈��<�f�(�z��_
=�~v�zo*=<�2=�]G=u�¼F�.��_<0q8��3<)�="�j�y�=�%�����<p�M:�[$=<�^�fi�<\�=Q\�;�ռ���<���;�;�a;=Rc<gݼ�~4=v �O�<�=�RY=gv��dZ=��;�L9= �x��hR�*����a���7������*��Sֵ<���<^�4���7{���V=��_�����[���}=Y�-���Q<�?�<�ȣ��8����<nV�;$�< +	;���#��I�ּ���<'�ɼ4�E=��<=C9=O��&�>�d}�<��7�Ni=����
������V��<�P�ǡx=<���pM�+b�<	>=����].�<�o�.�*���=��I=Y?J=lɣ�?=�D��2G=���=B�<k���fu������=��1��}h=~ӡ��2���9��=k(���G9N�<��8=�h&��;���P�:�Д;i`�=mGo�
�"=%��<�.=TSN��N�<���<_� =��;�1<�8"�2��;"O�<��F<��K���~=Zo���-�������<?�"��(��ɰȼM���1��<.5�<���p��<>��4���{�=R���w�6="A�<b�p��S�<4�?�E�.���F�Q�H༗�ܼݵ��ذ�Bg+=q����1�V
:�>���=��#�eR��&IE��A��-E�@�<j�q��4�;�%�;,9�w��ȏ;�,��#�\Vz_���=e�U=ꮏ��}#=~q=S�2=��<o۴<�>��L��3���=Y�<Ա��ѽ<ZI(;p5��w�=��4����<,k�$Y~<��>��<
=i�`<�2���5J=��������w��%A�l/�o�=gXK<}�4=�C��N=��@�{�L�������\����<^f=���^�=j&�L5Z�:��;�����R�=�d�<�ur�� ��+�<�=H��5�=YR��ִ�rL�牗<7�^���*�
|��i�W���<O�L��<�{�:g�<���=t�����<Q@m���<����0����?S=>��;��Y=����t����1�Q�|��;�6����]���^0��M=GE����p��b:�٤<$�S���Q=�� ����;�z�<z;o�E��9��Լ]N���I��z���th�<=�v=0�$:	��K��(���99ڼFH	=����k�ۡ���D8<�x4�n�,���w�$e��S���
]:��2�н�K�߼NC
= �ϼ���<�!<��%=mz��2&=��=�Ǽs�&=b�ܼ��ť=T:��$��d�<UQ��>=�-C�"	<=�<:�O4M<m�*P��3 �M��q�m��MϼwC�	܏<N=�s��j�<�߈��� <1�=�)2�m���F�F�<���9V=�0=�tx=������#�.�ʼ/��<��<��N=��T���¼�ƚ<��=�A��m�<�T<F�Q=
�/=�>˻~L�<n/��02/=�`�<C]=�:�H�;��r�	=����d���nY+<�*�M���ly&=�uJ<q�MR.�#[�=���;c��<D�%<P��<�}]<�輎u��}\j����<�=S��:?q=�d,���i�6=�6f=�Xv=~�,=��2�s�<t��;<~"i����-uB=a�������!�0���V��� ;�����g滢'>�9/R�g���!D/=�3q=*o!=e/=��;���f�μ�1=�ڼ3a˻Mm�<5�^�{MQ=�>�ۦV�2���ݽ�<�X�Sg���E=���d����g�<x� ��S%�x�=�/���ۼ��>;��4�(�<�g��<ÿӼ�7=�� =2ڳ;�S=�Ɂ�:�_<��=�=S�v��oл��o�r�<"=흮��7=�O=�j�2�r<�).�O&~=V��of<�:s�Q��w@��pC<��=�R��`5����;}�R<KB��͜<b�<E=d�+�V�=G�<$��hǼ�`�u���~�u�9��<�b�V�漾��;�����Rȼr���Y�A=��/=�������U#R�B�K<و;i-���w	<]��`X���[z�Uo���2<��q=�����A�<��8=c��<�'�� i=�<K�W����/���<n�����G=�5���'»��-����:~K�<OE����W=���:f_�7H=�GG�N_<c���U~	�Q�)�4K���<�&U=ě� �\=���<yϤ<��Լ��@=�*D=�o<�)!=@^Y��N�<z���v��k��l~<�&v��@B�ij=#n=�|�2E*=�#�r�=HM�<�����TC�պ���;��+=*��kN�=��=!�V=��3=N��<��j�����mI��3�<7.���;=C�t�>�<6=���<��8<��=�`��v;u�T��ؼ)��<A�;��B<��}.�<��<��<��j�B��Kg=yӈ<������ʠ[=���<hGƼG$Q=E8���%���ۼ�rV���;��ɍ;�5�<��@<��̼�"�<,�I��
Q=�/��l2���>=��#�z���R=0䊽'ʼ;?�m=3�;7�q=0��<3x'<�-d<|-=��:s��<c4��f<7��=v)<=�ت�0h��Fb=g�p=��=\
H��#l�~h=�s@�G#�j4=�f��{�<M6����L�G<��/=�̀<d�=J�缎m8=�(H=}B =e��:�%=��%�_~e������=��w�=*h^�t�ȼ6�UJ���=��
἗�u�`={��<��j��-���<{�:ohU������<�4=��e��<=H��<�)#���ͼce'=n��<W�V��j�<����(=O���~UE�y���*�|=��E;[=� =�/z��fV���=U!
�!ib���=�<���g=%)�G����*�<�l=��P=(IW�H�C=���;���<(�>��B�� BQ=�;����q5=e�K=f��<��;��>=��<�U=��R=
H=���=�~���=5����<�s4�N�G=q��L� =�;��$<7� �q���=�/#�H��<kI�<�`.=�K�X�K=-[=o@u;��=c����D���=�:�<�yG��B�<�^$�K�N� ����L<Ln#=��x��;m��<���D�:j�;��޼t�!�b�<D̼�:��79ּ��=��Q������"*���\�!:<��<�A�<�S6<ΩH�Tn3=>GP��n��_Ys���l=�I3�惎:Ϸj= �xo>��]<�;��T<җ�����@�;ӖV;��Ƽ��=�s��F<� C��
���-�b$����'��1=�����b�9Sݻ�. ����;� �%�c�;��4[]�=Z��&\O��פ;�c��a;����<�,ϼw��<f'�:�Sh�n�@�7�`=�M1<3G��P���S<?����Mj;P"��*b��^==�����h=��w=[S�;���q��<�1%���0<}�B=$�=Z����`߼"+4= =kӠ<U�<�L=t����)!�z�?���%=/.M��b��h%�<�<���<�\a=g��	�;���<
��N�H<F�����<ud��$3>�E�b���T��E|=���<7��<�1���	=�<_�<="��ڛ�J�F�+7=N<��d+;	B"���~;o��;ǁ4�]��?�;r�ۼ4l�'�k=�l\=�=��;�t�<Djļ{������<A +=��ƼA(�fX�<��=�O�<��<9�Ѽ�r{��a�<,=���<5ne��N�;�< ;�#��-i7�`w���=�<�k8�2i5�"C�:�I��m�*<
.�=K��<�)��.,�:�Y<����"7�F�h;����������<��j;���(j[=z�C=m.�<<|��H[=G|��(�;���9�9�w><��M�@�g=�m���ۼ���N=��[=�d=Q<B��Uz<-0=eڌ�?N*���<�,U<�m�:*��b�[�9=�����)�6ח���6;���8��Yo���!�q�(<F�0=~�i���q�T^6=�x���$���<$G <�P@=�=͗�<}s#����<��<𤼈Կ;��y=��<}r]=Y�|<R�8=�8��$*[��5�Ll���;��j�A�i�3��Yt=�������<}�=���<V+=ʦ�7�<��T�oG�lH���mf=z)�<��ټR��; S켕s^;��������q3 =	0j=S��<�2�<�Q�K�A=��̼X뷼T�U����;~��S�G=w��<�wc�����fü}�I#��z[��X8<�e_��	�<>�&�֒i��NM=��<�\;=f�<�:�<j>J=�ڣ��p��79=�$I�ZO=?]���ʼK$��aZ׼��	��u��i<//=gky=� ]�\�M�t�ͼ6,N�v)�<�FƼ�j6�=z<��Q�P����<����,�0=��p�AA��hx���=]�����K=^�Y�t>=+f�;���IR�;}������<����<��e�U�?��B�4���bDp;�`L<���9XA9/�*�u�;�(D��i��p	?����<7����\��'�d��5ڼ��ʼ��j=���(�mƃ�l��P��&;y=;�/���4����@�W���<'�#�=<~�#�1���|=��Y��3&�$�r<m�=ZCF��H =�+�þ���&=�;�#ϵ<��j<��^=��;O�<�a���-��t�<��)=eI��g9�.�T<8�6=�=8\=g�1��P�<k��<ld9=΍U�}���#p�<ߒ&����;бf<���<�d;o�X��S=�E���U�8=%���o=mr=��𼲚�<�OC�[�=*v=G&�<zB�9�v<�zN=(x~<�2Ǽ�"���b
X=��m<_6˼os��&^�:�[�:t���f��%�<<}v=���<OS�!?���i�� ȼ׿��7.:��]=E ��8i�VVb;U�<���^v�������;6��=�|���4�[�U����f��M0`�"�<��=�l�g�E=�ي����$�c� Y�=w��;��ļ}ż���"=�V<��<FM;q�d=��D<*�2��N<~;�fڼ���<��U��R=��<B��<��1;3���!���K=���<~�O�Ł)=���;��,=K�Z=qf�=�=�� -��컒��<M�O��q=���<�/��e�2��KW���>���5�j�y;�'/�r������T�<��q=�@׼�.2<2�=�3<\�J=�͕;��f=S���*K�Ǌq�r���Qi=������G�g�1�=������<N��'�D�)R0=��M=�lt�؟�<e�N�:mS��ɗ<�5"���8=4�*=1�;�nN�Ϗ�;ô��m�#G,=Џ�<N�<���wh]=���<�jY=���:x�R=)�g�p<���r��o���v_�a.�<Ԋ�< ��<,�h=c>X=�h�<��.=��$�D�ּdl�<G��_V=��;=B�<��=l=o��� K=�>꼛��<s�j<���<3<�rS�ϟ=�y�<gF�Q�;²)=o��=�<��2=�uK���
=e��U�ռ$���;B�7�r+��Ki;��3W�<�2��پ�P4m���<���<�ܼܭ��ؼA;z�������Ӽ*���^�<��ɻȏ�� 2^��B`=O��<g�1����7=�k=��=){Q��-< xc�z/H=s�����ֻ1e<p�軰k�<��-�Ƙc��Հ;B�N<�<������ü�g�2�='��7G�ذx<X?�]�D�{�=�����=��:�<�����3=P�ۻbo=��P��J<K�޼u�8���_=���,w�<*;N�&��u��ˊ���}�7Nh���O��?=�U��N��Ύr=N���u��<t/� ����D�ݧ˼1e9�Y�_�W@=�%J:��<o�S�m(=���~q%=,=O�:K��<��6�K�6=�[��K�1��|�;o-��ky�͢$<�򼰓̼S:�<@	a=$����_¼9B��<o�<�D=c&m<�:<��M;%��;��N��?=�=������L<?��:�R=��<��
=w�%�X+�;�i�;�7�ny�!]���퍼�6/��X=���]=���<z��;�bo���>97ݎ�M�<v1��#�;��<���<��̼LΝ<Y�6=��<�qW�K=vЎ<�Je�|ҋ<��=J����E��u�;0�="�����`�+=s�_�,��<h/���^4�|��FC��2��v�F�8����;�&?=�ͼ����J�<���s=2���+'s���<���<m(�z��<.��<}0^�
Y�=�[G�R��	�=��;����8�.d��O<�X%�K_��Bu�<�<6�
�����o�$� r�<'�B��fo;�n�����<�b �Я�<V<3撼z$=���y�8�,uz;�4���}�A���)䞻OY��7��<��/��^=�x=�9w>�<c�m�t����#�S	t���=n�ؼ����N�H��4D�1�&��$�<�<�<?$��>�9;�E����ռ�g�<�@��A0=���Y�����i~;=r��<Fd<�"�;3�<���<k=�<-�ͺ��<
>@=*>�B�1=H�#�>�$�Vk%�$xz<�F�<��׼H���S"�<�vZ�Uqy�'џ���V�z�}��}T�Ǽݼ�`���N=f�<L{Y�f�n=��a=�U�<�Dǻ��I<w�<�������c��<4O�bٕ<9�<���<�5q��h���$�B�h=$f>=b==b�h��k�<�w#<����s<=X%�;zV<�M���`=$�2��;=�p)���j=;H=R�#���-=~{z<o�<c�<�2a��a���H�0�<-�̼r�<`�(=�B=])=�1:=_/;0�s=���{�~ μC�'=�#=��W=[Z=��G��:�<j�C=Me�<!�;�^="��,�{a��?.Y�����4"=E�l��2=�ֻ��b�P� ��#=5"�у������+nI=yR �6R���<�� =.N��� �<<cB���7��v=Õ���=<�A��m=���X�6=�8	�(�D�Z6n�/=Q!=��=;����= \<�6=�D�'��<��$����8.<��M=���<�h<���<$ �I�<.�c�,�]=/�,���k�v�R�3������<0�P��	�����<Z��:0�<��L��ؗy=!n�%�Ǻ"�0=;�=����=����Y[��M�>=�K�k��}���x�<�׭�P<�V˻�:��@��c�����9)�m=�%p=&�<��R<��G�Tڼ��K��)O���<��<��H:7�<���%x
������-=����-<��m�g�=����;���d������^=����>=�Ts�@�s��2���Z�<��I�U�j=D;M==�Y�<�$=#��⼎<���<��<=Ƅ=9�伙�a�7�Ҽؼ=o�6�#��#���P=,��K4�<���������"w==W$=$"���`�x��<s>#=d�F�GKM��8���%^���=<(i�<�_���+���`��� =�f���<g�3=���:���2<�E	=���<������;�&��V==X�)�<J�]�<�h�Q<�h=:�t�@;��b=:�	�W^=/�=�ש���s����<�]�<Mjy=���<~#@��.4�c��S�/;*�;�,w'��B�<�9}���_<�� =�4=�+�=sƼ\�4�1�1;�*�n�=�jJ=/�����O�Ѻ;��6<X��<v��?=�?=�cX=�Q2=T�C��j_�a$��i^=(���������qm<R7=��|��ر����<ͦ1�3�ȼ $U=J�$=Pb������m=��={s�;�RA=w�<� �;#��<���<#�e:�i����X����w=La��^e���~<7�Ⱥ�;��<�<�F����<
D#���<�>W�<e2�,���@I���
����<Cu�룬;G8���k<��=�ED���6=��<��]=�=����<1YC���D9ܑ/����;�y��mo=r&3�/C=F�|�A�=�F*=5�ѻ;�:�[�=��-�e���'��<�l=�a=��<��\�X#<=��=�VS���!��@T=D�����N����<+�:=̀�E�=�q�;�?�;����c��5���6�P���pۼ��m����7i:c���qD��z�<�S��t=��=��s=��0=��C=Y�����<�}���l�=�/=�����@Y=z�M<2��<έ9���>�D�<��:���\�$����-FԻ0Pڼa�9=�,=E�+=z�~;g�[<���P"=�)9=7-=�`C={��b��<��;=xN�<��I����;��1�)攼��5�(9��w�����;���W$H=p
��:������ώ<�&��μ�����ܸ<��L��Jm=�t=�� =K��<h��w#������zT=���;��ͻ�~n;�����/?.�Iw�<�<Rg4���<���A�+=0S�:���<r�4<�8=�7���~4=\<=o�:=�<��<^v�<ؙ8�*8�z���%Ո�5�ݼv0�F/=����\u�<�<��ܑ�����|=2�l��	�e�=.�0=�B�<�;��`��P<�~���<" ɼ��=(�Ӽ[S����[���<�oܼ�X~��e=b#&<"B����s���-�/���(�0N<���<Fg;=�JH=���-4:�������<�X=!#n�-�
�N6 ��T�S̢��<�=o�8<Y�	��M���=��<�;�Sg�;�54=x��<���<� ���sR�*[��+�3kc�˅=5�j<��A<&�=A=��<�c��P�&=��<誄��(��h(��������Iz�<�4輎�a��)6<U�<A%����M�@�<��"=m%d�� =���;��޼��A���W<�6=�e=��:=(�<��<Vi/��m��Z��L6�� �����<��q���C=�lм��=��N=_=�x=+Ō<e��<�ƈ<��+�a��=�=bn�<P��R��ޒ4=��'=^9=�B��~s���Q=��+���K=X�h����wA��Zڼu-x�-C5F�ԥ<�AҼ�����Xr;ڳt=J�]<M`���<"��-��<��:P��t�<*BҼ���<������:��"�,=�b7<lS�v�R��"
�F���;�@�=J�<��j�R�n�Gn�h��h��<6#�; )9���a��1d=/�<�	#��2@=/&6�B� :V>�<�zݹ��=�|�<�&��A���DK��)�<�܁���<P��\����	�<�Ա��=�<��Z=�r�����i����=fh�<܎ =��Լ��=@�V��ǆ�D�=Ya�g�ＭnU�[օ��8y=}�.=p� ��e�{���D�%R����<�ǻ�Ï��/޺�kl��c�6�<}�j�j>��O��=}��<�đ�V�<�����1>�<��S�����pO�;�͂�/dJ���W�{

��=�;0=��<���}�<3�C��*2=Ƽ�V�;j�h���7Q��&�� 1�bJ��O�ݼ�˝<�,����;� �<��f�L�	=t�����<�/��!=6�x=S̏<G��<�i0<��R�;���q6��#��^��la�>���E��<�:�w�d<������;M���F�[�)f�<�vQ��,���=8�3=��G<�iX���<�tC��Q�;�o��}�<�yU�=@ɼ���<F�%=З�<�Ot=��"�U�;�x�;)�V���	������-f<��*= ��<l��<�p:�儼��C�4��S{�<��{�ɹ�)1;YE��X���������M�B�<O�8:��6;N��;���>c4���ƼA�u<�@m�J�-=��;�n΢<�=�4�<���<ɝ.=?&=�K=��=6�2���<.b�<��;=������V|�<&�X;ՙ����ߨg=�kE��x⻬�<|��I�!�0�#<2=��j�~� =��4��=+�<)
=V�>��!�<T4���5q��z1=� =��w=+����;�g�j=j��=D\��_�S�����.��&��<D��E�?;�"�}o�q��;N�\<��R�.���s<��'=ꈞ��� ;|t�<����:��ʻ#U=9�D���8�<�3�;�!߼n(P���]>=,��Җ=�-=��i=ޟ=х�:�R���=��p����<�L�<��L�P�=��7='�h�����1	�-�<���by8=[Nn=�;s�c�;�^�L�$�.��K,<1����r�0�C���<���G�<<RK�][�=z��T�����~3�mM�<�ۊ<'m=$����6�����<�{\��=�P���+��\�I�����6=��Tr���,����;ȱ =@l̼���<�H���N�At�<�Q�<9cn=���<Jw:Tsf=򳓼J˰=BQ���e=þk;�#�<r�;D�=�<3 Y=~Z<����<7�R�[�;�&W�&�=�M=�� �.�(�
�H=�D��_�=�и;��s<^4�<�f��|<��f����<�đ;�=?�M=�$��
<d�2�x�$�@_=�r�:������"��qp=Z};1u�;��;�t�&+û7��<���<�<m8��+�;�V���'�<9'=�a�<~m�<�軛�7=3�d<��<\��dG�<CO=�� :;mZ.�TPZ=��ܻH=�Ձ��t=
��$]���9�����lo�ʕI=*�3=�Ft=�X�N�=?v�<�"*�;8��0�-���f�<>=iU�<g�<�F=𶛼.p/�Jc=�|����?J��O���C<���;�s�<r]=��=[�Ѽ����Z�~<.���py=�~� ���������: �p���;1=��S<���*u#=$Ti�^�=�W�����������<��<���<:=�<mhX�'`�<B3=��<0�ٻ'�a=�P==_�'���Ӽ��=9w`=�c/��^�<a{��D἖�ջ�ċ;=t�<E�F�O0 =-[(�b��<
�\=��'=������<�;=VKǼ��;�t����k=�� �$ze=�՘�;��v=����u��,�=U�U<۪U=^��P�6=7E�z�z��YR<q᝻�q�� �==�7=ج=��i�J�;=���?Rռ6J�<�����B��k=��<=�3=)H@;��1��/r���2�q�<�6=��7=�ȋ�K佼g]�<�l=�U�;@���zB�Ed^=���;��5��<p�ܼ���l�\��?�<�J;C��T ��ƕ=8μ��<���]Av��(�<e��������;��*�ߐ>=�zD�5+�<e�Q=����o�#�<1���=�V�<@R���F=5
�v<�˹���;v�����,�8q���~�9�껬&}=��J=Q{Y=
ס��
!�|_!����<ڋ��(=���;�-��h�;��=�\���P���z<N<�/3�
=���	�
�M��ʹ@�����^=vC��WJ��-
=V��<���D�<�f�(<\���-<γ`���ӻ��ݼ�>��מӻ8��;N;�;�_}�sU�<Ѯ���@��3ሸ�o�Bf<�|?A��=�����;����|������;]L��;F4=�E�<n�8��%<��6�%:��<�y3<=���<GI伀p�4��`p��]�!�㼎)���t�#;��U<�o��\.=Xn����Ó#��42=�>�7C�!��3�?� [<�}���� =���_<cϻ��;�I�<(q����<��`��2��a=�gF=C���T�<!�\�4v�6<=5	<	}�ԉ]<�:�Y�M�]�(=\�0��55=zM;=n�M�A��<h��<�EN��xu��k6<��(��BҼ2�ż݌ʼVĆ;��8=b1��a�;� =��<��<A_�<�M��&����<�����[R��/a���<gȻ�\=�{F=�G=u�U�1I�<<A���/��.����)��`�x#�	�Z=fh1���<��P��N�|�u��=��'�/1���;��>=r��@\�< 
I<G =D~�<�6&=��̼%�;�`q=��<��<#h�<G�Oͮ<��:'>I=�A$�2D=	����;ou�<�Et�
�>=�?(<��<!�<8�g�0ʯ�F�<�HܻJ��<�\!�0`��v'=s#׻�̳���F<p���qK��7'�U��,m��)k�<a���<��6���J<�e㼧�<Ǳ���L<ͤ<���=��K=��?�gD=[00=��,=D%<XV���<=\�u;������;�� =�j���Su=vU���^<�K�<�`<�c;��_=�+��*;n�<�J;��<�p�<�N=��s=��'=�DR�����W¼#s<W�f;u�¼D�:�*����y�
B��O�<y�V�W/����˖�&R�<�ͼ��ռy�X<L�w<0HO��;g=t�=�oV���J��� =,9=���;�Po�y��<��ú����K=2��<��`=Z�M=��<�Z�<�G�n�=�=(=o _�}�6=dqR<�>P=B�G��>>�)v�<�S�;XQ���
��K鼭;M=o�8=�Z��-����@��m=9?N=^01=8�<�߼��=0Kr=��<EP��=~Kؼr�뼤Q=��_;
E�<}�;��	�<&�1=+4w�hW�;��%;RJ<[�4=�<�<L�=�K=C'��eq	�Bc=�&�->f��3$<S�=}���q/T�����p-=[k><S��<2&��o
=�����8�@��[Y��)�uX���f;�;=�ΐ=Uz�<�|F=`��<�=����4�<s���_��̈́<�9��Z�='����3=+_a�q�=Čp���4���;�9�7Y�<#��<Z!<��<9X<����M���:=,���Kn��l��$�1����ڕ���ټ�6=��;�D�;y���:V<��;c|����:ڧ�<& һ�Z��ua���<m�S�K?��8�<��輩=����~+=�,��cO=��&=+=���<ly=6���1<�s=г	<E@��܇w�l)=�4v��1=����r���<wC>���Q��Y��D�=��<础:��;�ܼfߣ��h.�����=.�F=h0�|$�;�X�<�,�����y�T=
8��Q�]��.��<X�ټV;����K=I9��$;��<=�HZ=<�;�M9=*$=�ռ�_�5:g){=Ġ׻�1%=��R�><���/�<%��<��<��6=_�b��9)�(c=�S�u�v7����]=�h��<b�E<͒�=�	��x%=S��+&�ҕp=VP�<ϐI<�kP=�V=�#'�n-=��<��@���%��պ;!PU���$�Ig=��2[����<��p=*����w�.qº9|���5=�
<�)!�N̼�����<��N=:g=�{~<]�j<%�=i[��=^�=�<�cA���9�����:=V�\��ZK�`�=P$=��4=q]��&�(��䪼Y��<g���Ա���(�<�J=c���󩯸����	�<�x;�ʊ��������j��j����"<*�k8��R�[=�N�8�#<p<�<�=,rC�Xߥ;�Ft=i��;_�N��b$=�=7Fq��RU=�H=ʲ��s����<���<2[�<>�M<
�<R��u���$O=��;�=��'<�oy��.0�09���FJ=�.�<�~=��ּK�o�x̸;�Z��g��L\-�d�j=ї����B=��_=>�"=��v=�B�|/�<�<��g<&o.=C~u<���3G=�(;�4=W���0�o#�<��%��/�O4=6�[=��=��u�����0����ݼW`Q�,�W=g�:�eP"�b�v����;)qc<��"���
=sl_��{���#<���;&q̼j���4=��1�RT=���;F#l=n����Dh��%:��	=qE�;ހ���P:��W��x��U#׼NT�<�L(<��j=,����UT=L�T�6�G=�[r����<�{|;Ѯ<����<�=�Y=���<z8 �Vz��U?��p|<M⛼e���s�]=�8���{�<mͺ��;h	=���oH =��b= 8�nu <�?�����<!�S=(��~�<�3�s=ԇ�<��K<9%�<��Ӽ#wd=ԩ0���<(�=xb���8=9�-��u��ڒ����d=3�= 
���v�<c�\=uQ��G�C=��<�1=�^x<޵�<�>�=�[D;�v��J<���~�\�==۶&=]����Yt=́H=\�=��6=W�[���e��1�<L2= =��q���*�(%���x���&��Qk���WZ��ϗ����%�e��<U0�<zw�c�j�Ͻ����<��)=B�,�Gnּ�o�;R)������������u����~�f�-=�l�b�n�qo=�\<�$����&��Xc#=Oo��3��5�<=�4P� ���<c���%Ѽi=�����O��B��<���<L�e��O = �d=��~Q��sw=,>=�|���gB���<�_�8�	=�<.���H��:��t*=�0�</��<�ԅ<�eO=z��`I�<���=6�]=~��;�c=#�:�/�<yY�����<�/,<2_6��!3�!(<dC��,�8�K�b!=m2|��#�<^�C�~@ʼ&b5��,_�j�=��\�SA���<�b��3]=�ڻc�c�ȑ�<��=y��Km��<6��<����N�ANH�
Qܼ���<��c<R�>=G9��:m��xW<_�<��%=	O=�|��8=w!=����c/ռj"�<�!=��=�����<c�g=��D���9�q=<�=�8<����S=���<Z����>��h�='g�<ۼL=/w=��F�Vw��ǉ��e 8�
�<�¼Z �
���kN���)=+����";%����źl�F=	�I�-Y=k��`d�,=lE�=�����.;�:�����J<d���pm=&��٢��-�=�?#=����=�2�<�#��ӌ�����=�r=ѱ=�H���G<��<��8�WԼ70O��|K;ֺn=U�<F���I<bB���:�SF�?j��'�</�_�G���;���<3c~;�kF=�]/=J.3=>�"=O0�<�d��ێ���1��ė�4�<(�<�;��A����ۼxJ,=J�$=�����f=�Ł=�X�jv[����r���5=��X��n]��_<���E=N�==��T��g���M���˼:[_�|Ef=��H�� (�t7���<+�(��8%=��1=��<��K:C=�V���Q=�Ѽ!r����#�/<Q㤼�_#<(ha��xg<��E��IB�v��*�G�>W �D|�;C�9;���ߖܹ&M�;Bp<jj�<34l����<�w2=�N=5E��F�$=��߼�D�l�S��N2<L*#�{WO=of0��֓�U$���A=�D0���<wh���;�Y���go���9<��=BC<��֤<:S��X-(�b�I����ֈ�^&��8R��x=�A�{<�\L�MQ�<�!z<���n1=�;/��1$�ay<:f~�<�,�J�����p��;�L�H�=�R7�MSV����H���$2�{�i���!��##=w=�j=AǄ;�q<������,=�-̼�ֈ�k@�<�(����<���jD�;P�Y�2׶��݈�x^='g=={>�=��N��y��<1h`=Ji�;q��Q
;��l=��^<�=:�=1x=S�黥���{�����!	����`O2<��n���;=��"=t�+�ǫj=h��<�_�|�=�n���=`�"�K����<F)=Q%��C&�3��<(�8�5sɼ]�3=� F��n=�8a��d�;b� =�n=oo=��;|%���ٱ<��^=��q��C;�m��9����"��U=�T�]�i��M���g<_�+�i=}3=��*=��q<3�C<V�Q��`P=,�-=c���󟕼�==e.;3ae��=}u�;�_;;F�(=
�n�oD;=#�����;���XR���=��]V<�@��W�;2m=�ȕ:�$
�����I�<W���3޼��:f�Z����wH���"=�e@=���;o�x��%�<�����I?<wL������^Ք�'t��7+�`1=��f�JB꼖z�<7�|�Wg��D����/B=��n;�>�<�+;$NN�N�q<�ad=�	m� ����X�x<Bz�<��J�����	����h��}��m�;uR�<C�4-?����-=F�߼@�=6�<-�Z�#_�;m�2=s��:�t�;�*=rY.�ψH=q�;�2=n�<=�=�?���h1��%D�=�I=�=�k:z���5��e��Ɵ(�T�=N75=��?�!��<�����?�uv\=~%�<܇ =C�*=��H=՛�'	���b�<Ո(��Sf=.�9��B�1�f=�=p����=�<�O��!�#�n���9T=�&8�e�˼>;;<q�K��N�zs���<-N$���i��CN��RW�@��@A<9i¼2�;<2��ɼi%�<vK�No<<�Nˍ� 4���߼'�<��a��*@����	!����=�=�*^�C�<�N�<�Ks��\==��e�7�^=#�:�y#=_���a�;��z��K������m��:^�/(�;G�M�(�+��)����~Ca=s�;/��<��;<O(=�6 �L�R<t������E#<��;˲#=vX]=k�f;$=�3��=a��<WTW��<��񂲻=F3:%#<��^���%���/=�#8�g�<`=�<y�<uG=�#�������=�,����<#����V׼���dc=��ʼ�X��{��׊M�c�*<t�x��;�w= �)=i�=#)x�?pV=���<��m�_�6�`M=�r��$�Zԛ��}b=ռ.j2=�=�^%=-�K<TG ���(=�g���a=;�<�A��� =2��Z�&=OG��K
�<{x�<��r;�=� ��ׇ��U$�M��<���Sۻ�[&<�mؼ���=Ll��Y=D���u��1U���v>=�[a���-=|�=o�a���O���=W7̻��8��߼R���=���<�&+=�l=U�1<i=�=��=$�<��0��;�l�<ȑ�~-�<mzE��:�<؛���S�\�6�E]��v�A���=U���XQ�<R�.���<}**=�ǻY�+=�A=h�	=8�y�� �<~,x<��f�PO=w�I<*=��<��a;@%t��A���.����<k� =I�;��N���F���'���Լ�B<<�y�������S�q׎;��?=/iY;v���{>=��:=0�ռE����j;�h�\Z1�JJ�^�� �/����H�=�)�<.!��-���<�с<I��<&l<BѼfPs<M ��o)]�"��;2t�<PC�w$���0��7J�ݛi<	9�<��$�N	=CE[�oy�<��{��`O���(_=O2K� @<C 8=Qж��%=5�#=Pq�hd����<wf\=Ӌ�:�s2=����y��r;���?��2o;/IC=R�u<	; �Fɐ<9�;d�!��� ���E=�p)=v<M=�b=G�]=6uB��'����<%�����������;��m���5=ņؼڮ��;=��0;@@=ud��\$2�]s�<�)���?�:�6�<�?;=2�e=1J6�`�Ѽ[�Ҽ8�7=�C.=�j1���i=Sի;��4=������<`��<O:4�S7<f\+<e溞
=x�=�=t�b�F^����fX�<'^X�ҧ`��̻���<���N���	G�:<jG<hC*=��&�;��<����0=cӸ<3�Ǽ�>A���d<Tuw�AX;�U=��[n=t1N�(���/֙�0�-�\l�<��{<��<�X=G>=��ۼG7�<V,�;�򜼵K4=N�<����A�=��q����(�&��=�<2���6<�-C<�EO=ڐ�;�����u��$��h�:��=�XL��-��6�5�\�O�i������w�<k��B�<T$=t��=x�G���=l�<�:׼���<�ۏ;�C:ţN� v�l�=RG+=U`�<cm��ba{=�̻<�2�<�8S�I�Y=C9-�06�=]C;�祼C�:SQO<z��;�T��e�p�s<�}�;�
 �%��klżC=K_=GZ<5u<�2�;�X�<	�=��[�~�=�G$=Y<�4�R���?t��,R=�q�<�d�<?��<��<d��<��;�n��O	=��ּ�� <߮H��e]=�Q��ߑ�+,'�<��x���Ф��n�L�KmJ��D�<A������v��:���7��<��O�lj���<��o=Zi`��nH��J8<���}��<�Nq�����K=�Ի� p�<{��c�/�u=��W=K�/̼��=ʼE%)�|ҥ<Ժ����<�~=>
<���%#n�p8;<./�<�7C�Ͱ =FL�T;���p�<�� =w�漨�3��H�,Ћ=hi����Q��d��Ѓ<�:7<F�;Ajn;B��=�=��<�<�]<p�;+4I<o��;��"�E
����+=��4=��=�L=t=Ȟ8���N=iq:<��P�� ��F<utt=i��<@�������=c����=���w.���p=�i=�Y=������ͼ���*5�@�d���(=��5(t���=��`=��7==s����+|������Q=�鎼y�R��F3=S�+���
�ż�<�)�^���n/���<�$��)BV���=2O�<�O�;*=}W�<��5�8��<�(a��^v=��<��<�t;v��<T5�<��<�(r<�G�~d
���t�o;j��;��#���<��<��Լ2�C�: �=�>>���ּ�tv=E�!=��<n|���+�;�7q=��a�N<f0=�,=�æ<�c3<k�ϻ =�ǂ���4�Ps�;�2,��A���׎=[�=6�$�n�b</gC<�%��| r=���<[ƨ<�Y̼� B��F�q>�<_� ���7�j=�IX����M2=$6@�]k;�3`<�5= ޗ<3�V���=��:����\<BZ=�����˺�Ih��§<# =�<��=�,F�$Q�)�==e��>��<)m)���=QI&����;ݏ"=����d<������%�/���:�Ԙ0=��:==�x��.��aS�����<����q�(�j���ge<i�B;�*��,D��_=����QY=��<P���n�qK���9�=#��<�	�<[S���t=�q <�*$�zMV<V��gU�<��=�j=�
�0�<nc��W�<�Ns=���#�==��<�����j<����<EA�������;?=��I=-O#��!������;]1�rF����\<0(
= (�	�=��1���j=�����8�R=������<�]�=��#=�!�<��)<�Rn������q�<#�C����9�n\�ʬ<���<#�^��3�<Y�<'b�������$��D1=�^Ｂ��<a(!=%�V`��6=��=hi;��V��2=d+��q|ݻM��;�D� ���|4E=d�=hO��A{�<@�<¨�;�<�W�zֳ<�α�o�O=�B=$E<$�ݼ�="�k=O�T�����C�&=?��P*�<�����A�%=�8J�W�&�F9=&��<q<���U;�M=l򻯻=�w���Q��¯*���?g�<������J|����;rU�:^�L=l�=���W␼X�j=�<�����ڻ���uI;��ͼ�`�<Z���	s;�
�>���Ի�)=\���U;=���1��9<%�	���G<nS�]�P���=8T�<�w\���c<�v�<�p;�T��g3=E�m���@��dҼZ6��H�4=#��<V�<_��<�+;$/���!��O�<,�=�K=�=�8R=�]����c���8=u��<ٔy�z4�qXŻ�k;��<�E=��:�����,������Ի���*�<)Z1�����<�<p�(=8_�<���<�%���V�`-�;l���}U�<	x��u<�2��Jn��T=���=.��1@m�ε+;�.�)��<�u?=��u��<A�]<�vH��K==�c��u=�(հ<�L�����ԫ�j�=���U�=��#=��;)rX=8�&�!��=3�;S;�<��=.�=Fݺ.7�v��;�;���U�o=q� =�$*����;x����(�z��;��d;ӻ��8<=SFa=B3�;�f<A�������_u�o�����(=��-�o�,=\t.<����:=_���0�=�O=򧨼%���z=!�_nS�g��x�;x)�<krּY'0<�߼�0h=��';@��j$=Q�D=��N�E2%��
�<�T�����<>=�T=�����K�:.Q�@<��ż�6��ѣ�y�P��㵻��<|���ּ�]Q��2<�|Lh�XՖ���=�fļ-"r���8��:�<�<�;�g4<[x<�+@��,x=ˎ
����:���T;*���Լa{=��c� V=�H��G?=p3�;]�d=n>k�^��<�����=&�<����΄<c=��<��/�aN����@=-:t��*�=jH����;Z�L=μ��<���<�И��%:��i3=�������:�^���[;R<-�L�ټE��Q�����<o`= ��F�p=�oA�)#�;��:�
�<w��6C� hf=�)�;���y{�	G��"�,=�7��A�g�U���,=������S���^=�z=��M=3(H�񉥼8�=���1J��!�7'��<h��Ӫ<�?$�]}0��5�<:=��)=�T�=�良�����׼cJh=
C<F��~�<c�7��� �U�<�c{�u9��,����Q����S<Bg[=�p_�cs�<��?�f�a=��K=��9z;={c^�u�<!�/=��/=�='&#��/\=�y=_�0��<м	=f����⼨�&=d��<�.�<�K=�6c<J}V�/���F-~=��=0#q��˹�D\�K�A�ݨ�J�ܺ���3�4�G��<|A*�vd����f��|���Ѹ:y��<�R<�a�)%�^=�7���ļ��<S�<��<����Y����K�c5���<�4�;e����w����f;~;��=u�[�\=\8Y�6��<'�=H<�?^=�7�<�h,=�����`�2��<-^M��S�<�*4�Z�0���<�v=�F`�S� =��0<�C=r3�+ �<�1s�H�Z�,�༓�
=Rb���!ټ��V=f�<L؅=C�̼s�ƼH�l<��D�3<<OҺݦ��P�����)���)�<K�;�g,<���E�(={�8=�v"=huD�!0=��\ <(O�9��<ۨ���0��b<=��
=٥��[�hKX=�H~�y-��;�B=o�3��:/=>@J���[=����&(=�����u=�<�!�������5�<�V=<7-<.���F�qK��n��ڼ�hO�������;y���v��( ;J�غ��ӻ�N�=\�_���t���5=���; �A��5F���\=�y=SS�<m�４�M=��C�=P���U��
��<K�Z<�6�<f���Z导�H;���-l<N�O�� 9�J�<�;���u<��~=��q<Z~��X���i=���<���<mRἉ:=kN,=$�-���x�Vު�}�<wjټl��<��_�Q�=<�9=��;D��<�9s��O8�i5E;%�мkj�6��<	=Ȝ]=K�\=f�<p�[�*=���<�r&=��=`wZ=u��<����{D���B=�a=��<3b�<�d�� ��hn�����w�m��e<��	=@r��=��?�f������ 8=��N�2㼷��Y�V�.��|��<�B��XW	=���<N<2<�&�<����䦺94�:��<{��<��;��(���<�C���ػ�w�����a�<�?M�W.=%^�<��]�3<=��=��&��_�Yo����]<a��<�s<�UL�pDJ� ��=4�����=T�1�5��<v��<��%=�y=��0=5_�;�b���=�2�9��<:E1���һ�<DvT=��Q=��D�.�y=��5<��>=�_�<��p�=��μ��=ѻ7�x�7��;��ݼ�{?��f=���<�Z�<d1=�(�;��
=2��<e�=�`=�\�;�C=��{��Ȃ��`�<E�k=V����U���\3��[a�f�伀UA=" .<c�E�Z�J�r�����9�gf2<�@���<���=����*Z<������=���<QM=��ٻI��hc�S4��-�<�0(�V�;!0~=l�
=m�1=ǿK=��7���R�3���F�'�X�!�4>,=�d�:�9<�1<h��r��8���<��<��20=��8��6Aa;�b\�G=񇾼\�"䟼�.��b���="�=\:=����J���x�g��[�{\=�;� �"�����m}�N�c=��=�
��E�/�R;�f������}�<ܺ$:��:=a$�2-���V8�<�J=�M:=b�[=s��<5�g=����<��F=�����;쾣<��<���<=�h�<�ݼ6�/����</j򼛿��� ����i����*\Z<0Gq�0��<-���PW���<���<i��<�s��0+;�6=!�1��ƀ;�����8>=$�d=�ކ�hN�=���<���=yV�<�Y� �1W<�e@��%��q��#�U=U:�9c�<�z�<�>���i���<��9Դ<2�=�� =,Q�=
��<R�<#O���=T�ߺ��8=/��<[��}�<0����N=�Ǆ<��m�권= yf�?�6�:���O=%#��Q��<�?���t��[;q<Ǽ~Y��� =�׼�"�;�0��\�.=黁���=��q��6=ˑ<���!I=I,D�1�e=�E=	L�o!@�M�_��z�y4n�F���SY�:[�=�V�<�"<)�߼A?�����<��<�_9���C;�<���g�j���B=��м��D��o2=�eO�/&=!cF=�,o�I��<S5���=�n��e�<�ļ�Pa�K;��~=�=@�=%ܲ<S�V:��T<`�5�J�<�6}<?��:�#G=xn��p�=΀M��4��b0=v*��Sּ+�� *�����]*p<�Bj<�A=#⼼^>�N�.=w�`=Ҵ1��&G�l;��==�Yn�Oσ�H�4=>Ә�8��<<A=_^N���+����<���ڃ/=n�g;r�Y�Y,���=:�mT<e�һ-��<uw�%[��i�S<+S=�=(0l��;Y��iJ=]��;��&��=C�мTw��� �}׼;(=6�k��ز<�ֻ�ɲ�[��<� �<���<
J�<�wɼk(=�*%=��H=�d=ع߼a�*�C=�{�<��
�crH���\�S,N���f=S�==)���=�X=k����:=�8�2=E�M�<��;��/=���$�N�Ռ
��dJ=�ݩ�S���`=S�J�;h��ųH�+�=��$=�<���Grz���N��=j@$<x��JYZ�?�T��W��o�a�F,Y=q���=�H1�(0~��]��A�<���<ªR=��=<������8M<y��U�d8�q���9y����ռjz<����$
���U��(�<И������Ӻ��J�d�H��S��g�t�i<�N�<�sA9u�Z<ǂ?=�T��XzD�W�:��A=}p���=�4d��տ�RfN��-���!=�z��*;�P�H�(�a�A=E�/���Ѽe<��?<n7�<qă=e%w��M����<�b�<��<y�g=:.6=�[^�x¼�ft�yҼ��O;��9���;@5=D��\�B;\�y�U��u<���v<u��"���jz�Z�B<�tI�06g<��=���_��<A{<�7!=l�H=�?@��z���A,�
-q=&Y��ۘ<$:L��>=��=����<h�<$s~<:�;�3=�-λ��I(=��O=y5=n��<���<��=B&B=�ڴ��#M=�@��\=�GX=��P<�!�<Q��=	7=f�W<�1Z���K���R��u��o�:����'����</B�X�y<��;��;=��/<2�><M�<�_2�D0��4��e@<ٔ���r��2	��<�]�:�2^���=?ǀ=�>���^=vE<�=I'��C�>�0�`��F=OF�<��'�q0=�?F=a?5<g��<w��;���<��9=�|,��xl�k1%=�4:Cl�<������6�D"=,�D=�N��%,=�90=j$p=����vĵ�����i���V��<�6$=dJ�<��'=�'��*=��8=�m'=�	@��˪��@����;7�ټ�:+�W�m<p�����ּ����(=*�g�����W�<�Ol�Y^�:>-^��[��=�=76��=|x�:��F��Р;�Q]=���<�p=����)=Qf�;U�#��l�v �;Ƌ�<6�Ƽ{b�<�z��-p�<�7=	�Ƽu�e=�M ��C��&��7Z=?���s<��D=G�c��`���nE=���=ǐ?�	U'�����C�cR=�;=��;�5)���ڼw�-���E��G��$(�`+{=����T���Zz<c=<1�:G���Z=7���վ<�j�;�[�<��?=M^�|��xQ���⼔�<T�b|=25�;����]�39�w׻�;��׻
���� �<�&y<�%�<\\/�"M=�$W<���<M�<"����T�<��o=���<Nz�;�u:i<fZ=��<BF9<l��<��b���/=HxJ��뗼��k��i=`H{��5�bd�;�Ǯ�qn�������L;^�='��-�4�j���Դ4��/�<�N5<QrK��=�v�����N6��iC<�8/=��=E�ü��6�i�&��`c=RQ/�B�z��"ż	��=���~<���<��=+����J�<u0Ӽ���|��<V�G=��<�G{:-?<�,=-�:�����
�<w;W=<��������l�C7�<�:�<X�=/���q�<��R�����঻ʡ���ܼ/:<<l��� � ���@"=���a��<�A$9w�A�v��:�2=T�_�t7��p B��3=@�3��X����H�t��O���F�/= �P<�6p�C�W=_���� ��><�`*����oi�'�'�32�<7c"�/��ŇڼR� ��,����q1�<���<��f<�=�Pd�Gw+:s�=F&]<�O��#H��Z	�~c�.|��=�\,=�H=EQ
=�ڼ`>�;'�d=��^<P�F=)2��Ժj�<3��I��_����<�y%���O=�����E=`-=�5=C�H=H|����}<�ջɁ<p]̻��<ԩ�<�,�;�1�;���K}һ�o�<��'=d_=��<��^��<�4�<_�<��]<x�ż�Lx=�H�<>]"=[�<Brp�	�=ˤ_=A2μ��=LD��T����<r��<�]+�Զ�<@4�<� =�'��s]=�-=�n������� ��D"=�J=�^=�¼,�Z<T�=]�N=񚧻:�J�(bu�9"�;���%?	=�D=�Ʉ<��<��o=�J"���R���':��8=z��<3�V�!�==*���/��8=�к�ͼ)x�9�H=\��=v�˻�򻊜��}<��4<ҡ����=��&�2����������tJb���=��{=�86� 	μI*����o=3Ԁ�ŝT=��F����pV<#�;�Wf���8�!�k<@4��Q"R=B[8�~ƀ��V"=#�!�:����`��NӼ�zI�Hڿ;���<2�.<��=�E���,�<�� �&��2p=�|C=H�Q=�8=ײf=aY:��@�<Qr=^�kW=Qs�<����-BE=>����#��ש<�=_��<�J=�3=��<P^=G�� ���<�N����T��N==�=)�=I�;]���q���<�p�=���<�J���H��q�;�-�����D��<Q^�p0��Bx=6�;�����)�<l�;�,��K$=�[d���#���<q�<�.=EE��[= g�����
�<W�=�="�0aH=0qQ����'1=�L�7*(=�R��Y:=P��<��.��}"�r=�H�<��v<��/;�̸<p�=B�l=�=/c<3N=Z��e��c��7��������ä<��<B�b�5��A�һ�a��9M=��8=��W='��;"�<`�<��4��@\<��=%�8<��Q=�� =죧<��(=��<�}w�jIY�j��;�С<���ȝ,��)�<5E�<M9F<�3��l#6<���<���LL=����_a'<s[B=�~=dp�<�,�=oI�<'��<�J*�!���T7�<HHS=���<�\��e&p�+�/��:��A�N�/:^����<%my�6�¼��
�������=�
��34�-<F��
-=�z�V�)=;����7=�!=p+a�"��<@�r=VY%=�����<C�R�<?g!;�� "�z������+x:<�-=�0<gX=���=��u��CV�3���,-4��K��~F(��ѯ<ֈ��+�W=�h{����:�h:<�<�Ɋ���<e��<�(ȼ>�<ɯO��0+<��m=�
a=��
�?X-�f},��gE=-U��^�	���	=YZj<=ᒻ��W=��S�<}���,��0�O�]��@$=k��<8�=Jc��uyX��<`�=��:Ó�����<��û�;o==�<����=H�<�;]�d�=IM�?��N<}��<cg=e�f=��^={��<H�='w�<Ca=�7�<���ث�<دm�jus=�;�:���rL���;�MZ<��=O�<�;Z:ӕf������f���o�<'�l� �K�#�2��8+��̅��`<��-=�U�;��c=ש5��=��8�@�����<(��<���;��<��	�_����C4=5<��B<���<H�T�7c�:��%=���U-=�CO���i�p򼫊p=&�#��4�����G�e<U�-=��=��Z����<�M�3J���T<#�0=62��	<I*�^�@��P=\ ��\
=��<'�M��u����<C#�<15=�� ���'=�t*���>�P�B�-=��i=����$=�s	=B��d�
�<��;=��)�-C(=�G�LQ`<b�;V��<n6c;�{�<����F��;�@:��5��I=tD�=yG��6=�C�-�1=���<��f�������<Mҁ��Y=��<� w�xP��v��컽�T=�W=�fB=�g�;��z;�~��Vj�t�*=_��DN�;LM�.�:���Y=Q�v����<ƫ����}=gΗ;�i�<$'��8=��==1ې�8kp=i:��%�ϑf=�!�LF�;-Ր��&�<��[=��H;���Jƻl�< �_=}=�T;=V�_=�*�<b>�;+�%=�<�kb=i�<9��<���<*k2<WB�<�V]=w%O���:W"h��_��9�.=�G|<^W�<zBA<�^� e=��:�^��<y���8��N�a��4�.l�D�I���3=��A�|�L=�g[��׃�m,5<�Ѣ<{Ǽ�<L.J�"T7=�G�<�ԯ���;~���fF���<�\��ۻ�[�y{:[�L�n<�_���e)��t=9��<�T<�-���<q��'Xʻ�Y<a�-=�<=�:<8�=�V=�;=��:�*@<X=#�y�M��._=�L���x=�I�hT���U�ז�<�g0���.�Ē�;3�'�{SP��:ӻ�*�<Z�K����<����N+=��?<,!���ռYR=.u=)3��S.=�
�<��0=�ۂ<5�A��1�"=R�W=�I=��<7JU=��<��H���<��)��9(���;��g���c"B�ӼL<N$L�@�!<�nU�b��"�1�r�<O�����7*��ʼ��=7�H�qM�U��=q�h=��<�����<���i�V�=<�&����xs=������ؼ��/�/3�<Ʀ%=ƶ"=�R;�E|�<���:ઢ�)�Q��A=*�<K��<�7=�W�<Ea;�=�Ҽ��ϯo�%=���<1t�>&#���#�u5�;;=��<�[=�i�<HH-�o��<t%O=�׼%G==�EP=Ԯi��qi=��8�:���\=�i�;�'�֘�'�S���߾q��.c=�_=��<�t���=]�$�&�7=�V�
���$J�#<��C=��[���;��=Ҽ^=X;�ei==�=��!=q�<�|<��u��Q%=��}���D��^A� ��<0(�<���<;�i=���<�����|����;��<�ʪ�}�r=h��pm.��}�<vq==�=���<��?=G��uho=DJ�/�����b�%��<m�d<����<P1��/��'Q�+�<�#^Y��ŏ<�L�<�[i�^f=�p	=7qe<��<Tc�yS�d9<�DK���E���Q=�i=�3���q;�7ռ~�<�5;�MD&�x�<�F=a���Zp�wI=ռX=�=5�8���$��<\f={,޼���D��<R�<��:;PwE�^G;9��<2bv<%�=i�!=������H����<�r=nk0���	���ϼ��O��{I<86J<�1= ���	Z=<H�<W� =f���S�o�/;�!-=���AN����<�=d|=�R��s;��_<=B�f��<�<_8=Gh=���X�ɻh�<;�����<W�=G?�2e�<)�<8�w<H����W==w��<p�=A��<69{:~Xμ:)�Pe';7���9G=�ġ��r�9ycQ�@��<��L<�g�<���:�8=��=|����Z��<��N���T��f�C	�<��`���_��c�9�z��ڨ���R=�S�<U )=jЖ��W"��OE=�2��x-=�O�i�=<�V=x�}=¥$�ԑ�<���<���<ld��(*z�`����Q=5���<w�)�t� �}i!=
��<b�M: :����<�Ѽ��1<�
7=�{K=�|��� =��v������-i=8��XEb<+��<�����}�d$����G+a��=�����û��O�{�9���==ف�:C��<���<��=�HҼ�O=��<���<�r�<��<=G�.��\E<+�;��j�,��;�sp<'�;��<�i��ג\=.����O=��=|lG���1=U?<MX��S=��v=�+l=�(�� =�g=E=��G �����&����<�������y��;ᰂ��L�c��<�^=�J�<�} �3��@f=Z�=i��;]&�Q�B=��:!�2:
��D=��	=�]<����]�;=%ֽ�)�]��B
<� =Z"=�)C<|�<��V�P�\�o�<4B(:�)k=�'��mc=E�C�3��
=�9� �#�W׾<��H=�x=���<GG��S�����<�S5=�O{���*�ݦ�:)ӱ�v�>=��<f�1�]�<��야�<�6H=Q x���ûvOT=[���D�<�@�� ��Eߥ<��F=�]�>㻃�_�A�?=�*=�9���Ҽ�"=9s�&�c=3��;Z�==����'����܈R=�l�;�:Z�ďQ<��9=9��0�j���<n$����<�-<���#=��� �<	Z�<_Av<˗5=/P�<���:޻;���;�\���#���<�@(=ɱ�<�sm��-�MR�:�0t=��~�uT���6="Ζ�j���1=��'��1�<C=�3�<��=`�L�w/f��Z��pA���� �IY=<��v�#=�f�;��N�_��(8��S3��Z4=7��a��<���<�D��_��6=�G7��9`��VC=z�㼘�.=#�<P���(��:�f<LP
=�qK;��v=�{P�)Dw�|m|����<�9��6%=)3��Wy�<�gG��<݆�;�d^=�	m=(��:�؎<��<-�=�G�;R���&a=��.=��,��<j�;�H�;4T<����K=�����<�\���0=JD�;0D}�c<%����<�t:=o�'=v6J<@�D=^���k�85�=�7����<���<�%�<�ۼa��b�!=�u�; <���]?=���;�˶�M;�d=�-<j[R=�;=��*��iF=J�/=�:�zt�S��<`_�<AV_<��ϼz�K<�G̼�3F��<�< +��THc���<a9=E��"��<�_d������l�M"<�j���U:�<A���/d�~���M�D�ϝ"�*"����<QɄ<fo�,�u=祿C�ؼ)��<��=����>�����;���<�l ��A���2��o=��9��Е<)@�9�T����<ђ�<,��oK&�N��<�<�<)`����<�C'=�"=���<@���7μ����	�������zC�A��|pR��<==vg=g�x=���fp!��`�<��b=� ���ɻ��a�jH=���g�f�vWS=!�J=ߜ\=��;���<��ռ�W<��i<���MB;!�ͼ3)<i)��� �������<������ =�`=��~=�an=�1�l���a���Z������X�;8����3H����;���<1ta���+��ʆ�#ٓ���=�Z.=2�b<�oI�6�j��
��j�V=eI=��޼0�:<� �<��<X�n���7�<���<�@��{[v�A��<��"�=�w<�eM�U�<��5�*�<	�=pٻ�t�����<�tA���x�E��<i���h�;�$��<�Q�x�=U0h=g�l��LL��� ��i���z�<�=��i����<D��
Vl=}`��7��<n	�G��<�5���=��J=i��#�+���
��� =)��<���<Nz_=�M���=xˏ���J=�Lۼ���<���<����J�x;�J�e�@�r:<�b@<ͱ$�I��<��^=K3���<r s�8�:���:c/��4=S�@�������	ؼ(��~"a=��=r\��bt=�[�<��"�V�A�^�=n�=G���=@�6={=�w�<��} &����;��V��䄺7H�&	5=�B��Xa=�c��Fy�I�=���;=�?����>�PW�Iw!=��=� U�a1�� =/��<<Eﺪ�q����<�Q�<� m<�'���T=5ͳ<��6��?~��r�<*񭼘RF=�������31��ϊ�<�����8Ҽ�����"�a�;I�E;���"�<،G�C�Q��ƅ��J<gw缬�d�a�F=S�J���4=j]�<��H�1�ͼ��>L��<�y�<�
�F��<FW9��K=^�7��(�L�N�<��=F� �Q�;=�3\�6��:c�<��	����<���<4�d:f�����=�w=s�'=�;�2b�<�=��,�ƺ�<��<�G�򇫼��<7��0�ܼ}T�<#B���H<�)� �<w�5=�VU���<��	=uT�<(s����J�5�<�K��g�<�N�;��B� T�<c�:?��<M�"�u��<ݫ��L�=�<O;��+��X=�A=<��<���lk�)>�<I<L<��#�P��+U#�Ԓ�<�!�<��>=L ��S=�p{����<�~F<����-D>�H�;��T��-W=mF̻�9~=�F'=*9��O���#_�N8�<���;��<( ��_;8�F��m���&=��T�<�$�:�<Ԑ���?�<Z\�<�{u��\����'�I3��β<�2;"��<��="˂=2�N�)N�<��<��l�H�?8���<���0�ߵ3=V����=���:�J�����8�J=��=�
O=|\��V_H=.��;�珼1�Ӽ�:X=��=�y��0���G<`<�yF=+!����R(=��I� ,S=(�=��?�BA	���g���]����Q=�H<ֆ�ݰ��6�==����:�v<�>���ټp7<�'3�*^����H��g�<�U���<A<x�?=�<=��8��h5=ee=ݼ���=����f�\gg�<l�<��=��<�+=�xJ��QU�J�r<�w�<a,=� �<�����1=��������wa����;a8H���<������;�=����<����<��b�.�6�C=jg�:�\&=z�M<i��J=~_/�!�z�&�ɼ�l=&�9<D
T<�|]='���0:=x@��5�:-��<�Ά<�!E=�����k�?v=���8e��ṵ�l}=v�&=գ�'�n�k��慼��-;1��<jA�<e�<���;ǧ�<�k�;�O�p�=��*���"�s�;;�/����<q�?=1wX=�ԺF�9:Q<\t���	�<��=x�=�m;��NB��,!=o]Q�RZ�<���q��<mU�6��<,~Ǽ��)����Q1����B蚼��&=my=B�[���A=�Q<sKu��n���p�kmO=j�T=�i�<5���ו�<�<�p=��X=�{=�"�<iw'�Mv=������=�K�&�鼤P=7�뼌0�:&4��?=�=����+�;�@!=���iI=Wԕ<Vn�;�~\�h�h�����<�9F�#�=��I=���>�;`�o=@���D���<����e�V���&<�=nF�.2�P؇=�!=��Q���"=�&<~��)9����B��!ܲ�9�?מ�M�+�+��G=�f�����"i�2~5�)4r=��<��<�jQ:���<����E<��Ǽ
�=<w�_�>đ�gcK��j-���M�aw�;�~A��$9��,�w� �%g��/=�*������D�އ;=�.���o̼�7=�����g=����]����<a=9=IK�<'��8�L��t�;�C��=�3�<��<������)��gH=�	�<�b;=�Ĵ���=�-2=��U=A 5=4=��A�	�W�vQ�<6�����F=yDؼ���������	<� �<��v=�-S��.=>;�ָ����j��<y=aQ<���<�-� ��5<oC��c�9�W���]=ª=QZH�=�#=MKƻ*�\����<4�U=(,�:�.�=�M=sK��	�9�\=�
<��&=z�R��/=��(=�pʼ���=�#�.Ȣ��;=�>�x����;����Tټ�DF��t���5���`�ra<�=ĠT=܏��t<+<\냽8,�<o»"c�Pd�w{��<�G(����}���yUP���<�M9=�5�k~+��=U�ҹ�<�jy�6��+u�81(�x�����?=�^<��r�f��,����e�71`�]^�<|�s=����m +�$Z-�R��;�Jh��!6���;�:��U��;����\?%���<i�Z='�%<�Dټ��2=�CؼU�<Gʘ�y���Ir�=��N�?!#={�W=�뭻t���>,ɻ1ڐ�/��շ�.X�:u�V��®��y<%EQ��/��B�F�U���d�\<��~�a�Y,�aC�SrM��rz<���������=B��<v��<lW]=p&B=��ۻ��<W١<�^X��*ۼ��\�66=U���o#����;ޚ%��29�
ʛ�ޯ4=�Ի��h<�]�:�N=h����;\�<N^W=V�ᘫ<(ӱ<v���Y�=�t�<&�h=��G:Y��k�:<����K�ؼF�Y���� �5=4A���Y�͊#�8�;�~=���;}��<�ڼ�ZW�j���#=?&)���7;�8=��>=��L���üx��<*�̐�<ɫ���:�:>����2@���x=��<B<=ot�[��<-<� ��8����[��N8���<3�i����J�<�;=q�z;>Rz�|�<=��p�?jd��E)�;�'����<n<�'gt���R:h��5�=���<��w�OWT�᛼����,���<�#=��l����:�A��Uͽ��=F=�JI=�ż<5?ҼGG��5&=�/�;�c�<9L%=��h=�'�p�Y=������Cd7�[W��/<u�=���|����o=�d�����`���F�iN=S�(�:������Q�r=���<E����E+=V�<�{s�jl�g����޼�.F�����m����;A�s�S�v<�!��?(�ЕB=��;sQ�<�&:�>�<Ĕ��r�ټUJ�<_�|��P�k�f=>�F����d�[<{r-<q�:h�/��^<��	���5��:i����]�<����,;\��<�����ɼU�^��_
=���<��)�R�B����<6&=S<�<̹I��M����4�}:F�
c�<;�T=��c�3�s�8�U����nu���B�PKB�
��<.C(=��<���<�>���4�e%�yip<��Y<sH�<E;=T��g��<���Mt�<b�J="x���9<p�<�<ycQ=/G=Zk)=�0)=���<�y����(:�s�Y=����wQ=�b�<i:���K�����H�)�O��<�d2=üI=�F@�
�<ݝ`=���m��<���<'ټƀ�<��=+��<��<����0�����N�g�Ӂ�d�X=�&��k8�� �����Y�N�N&�<��~=a�<�_a�'�x�jЩ�qJ��kZ��B�<�]�<2�>=r���F��|/��O�9^���7=Eg༜Z�R�	�������<)ޞ�R^���Ѽu�<�źW��=� 
�����\P=��ȼU>��2ͼG�<��6;���;^�+��s�<=1=�̤��/Լ3�޼+R�|*�(���$���k}��0ټ�=S�<��;MP���λ�mv<p�<��<�w|����-��k��B;L�$4w<����:�Ly��r<�_ͼ�7ϼ�=���=t!�Z��<v	�(���~�<U������<�ۅ=R#��<={=7��O8�vV%<P�r�%����5W=v8<���<�4��`]<.å��HJ��rI=��j��B�<�㜼`uݼ�Lۼ9�����-= |�<��9˗ͼ#b	=}KQ�F�ʼj%�٧<}	� �W�Bv���c��f�_��BL��������:蹅��.������i���<k �<�Qj����2)j=�V���C�<��<�;�5P�;�#4�[���c,��P=Uk�<�P�;�=�<��<Z��s��¨=���<,j%��w�<�H='�=I�=J]F=+ġ9}� �)��e�L#�:�V�<�����=u=����:�+g=��i�A�=Î=U#��=Zuh=��+���<���9g�5)Ƽ��\=��0�-1���DA��K:@1�<��;=x��ƣ3��kt=��S�L�+����{=��;������=�/.=Ia�+�P��ְ<5���T<=���<�����Q��uN�V�<���<�N =�ZF��>u��b0=��=�'= פ�SG ��6�%�S=��<#�6;�������<�ķ;TE=v������=�� =b�'=���A=a
'=B�:z�=��u��b��2ݼSj����0����ڨ<��<F�`<��*��L8�}�A=I�n�4�)=��$�|$��e&=2k�<`;�<��+;i�=�<=:$���6�$B8�dȻ�W��{�<�*�֣<�e=�%=�K#;�>=�h�=��:�a��I��5+��vr=Uwӻ��;�@�JP��,���sa=�ff���nv0��}��&=l�Z=��f���Ǽu��9c�<��<`�<��I��e�<���;��'=�\b�h.<���<V��h�^=���<�/'=!0��zK=Xu���8=9��X�=AXw�L�9��kR=��<�=�5
=��;��L=y�ּ[8��=��NI+��޵< B<�
�>4E��v=t�<�]��hO=Vڤ<���<��;SE= Y��4�H�Z���ż���R<#�c��`=���B����)�6*���T="�G�&�����r=�b=$�6���ȼ�!=�Z��ų�<�b��w��<��8�h�<OY�<�?/=�2¼Q��<d�j=�	K�8���͂<ڥ�<�c��ϼ�$��<=k`=aJ�<<�1�,5�;q�=�1�;�0D��ZK;IVV�"ͼ��Ϻ������%= �#=sd�<o�ٻ�0����+O=ƒ= ��;3»�7=W,�5�N=��=��M�ƃ����&<|�n��ƾ<!R�H�����:�=��r=�Fk;�kJ���+=)f^�Y,�y�<���;�i;��A;"�<̱�;4�ƹ#n=�a��Z1�RQ2=�"�R�2��'P��=-�L=�=]�a��.��!t��y��	=�����;	�E=�v��!��Cr��Jz�:��t��y�1�I��V��z��\�7=c�~j<c׸;8l���ȁ�sE�<Y�<+~��w�Zb�:�� =���<cLP=r�����]�@���(=`�Ѽ΢�=F��<pDq�+xj�x�`=U?n���<d!l�L�9���7%�\j�;�x�V����< �;0��n����d<_�2=pO;i=��wX�<�#9������c=}����b��ּ��@<YG�%]$=��(=:=;5����<��ϼ#�=��D*= W�73,=�l�=�r���-;��94ہ<�li���Ӽ�����6�a�A=��J�L��^�9=s5=�%f�UV>��+=g<=�勻�!�<pټs5�:��M�m*T=�P�<q�lѝ<�@�OR=W1=h\���~:v�����q���r�<�T�0�G�P�D=RK׻����~�=v�=�8M<Nټ��:��:��+�<&�f�P�]<�<�ȼ���꼽5�d���)�5�S!�<J7=���;~���M�=~wF=���;}����<��;�G��e��X�L���==*-�a�<��%�d6�<Z%=��<��=<r�<�yO�mh7�X��;=�z:������!<D�=��!��S.=;@\�;��<j)�<�$b=Sj�<�8���ҥ���żI��<K�<���)���d3��i���Q=�A=�F��<��x���~��J�s �xN;�&�:< ���c�$,<�́�r�>=M]�~�2=[	o=��=��+<s=~�=t�<�.g;K8!=C=h�<J=���<��<u�@<F]X��J�H"μ����Uꄽ�+��";��<��K=��F�֌W�x�K=Op�<D&�<��u�d =p����;=�0�<i4M��ҫ�������q�߼�;<=t^��L��a:����;ttP=��b<J�<# ��M:��Y==G�gU��w;���TNw:�,�<���<��	�K��}�;I �'�"���<<���%�K=��Q;�o껤�q=��=��\�ƻ��<gJ�<&Hѻ�u�	ǀ�����!(=&	
���#=P�H��Z�e,�2��<	�=����3�L.=��;��<)�"�-N׼6U=��q=��g=0>��9m\�����<P���Y<������;�2߻��,�r�=WOm�JBʼ��<��w���F�=e'=�{9���!��=��0=m#�̋<<Lڼ����&�<׈D���j<�8=%�a��pe=	A����=��<�!��c����p�%<P2<� %�0��k7t=MG<=��8;'f=����l�<DK<<��T�<O=��_�𩩻��<Y1+���C���� D ���`<��弎7̼��<c�;V
�=v�y�z�>=8�<�/�<�#E�Trk:Iм<9Z*�F@=���=�=&��<��<�;= f����(��4�oᨻ��\���N�D6�<��;��=K�ѻ��H��'=	v��N�=�����H5�$0���K�p>&=G[(<@��<{89��>�<`��!N�X��;x�3�:�-)�<�B%��Q	��/�<��1=��C;�|:=�=��引�=���`�����<AV�<�����<��ѻԃݼ���<aqs����+)�
��=�Dݼq�=y ���W"=�5�0�=�(;�����\�Yk<��м�����#q��4�O�M���T�=j�Q�� ��3��t*=��K;��'=�� �=	���k<��+�:��;�oW�f�.;.ذ<��^=�_��<v��d��M5��%=�e\=0�=*X|�ɺ�<�<�b�6;�q��<�.h���N=���<���;`(��[^=��p=K����<�`j�^�E��Eʼ�M7��e���i�<�չ;'���U`�D<��1_=;�=ޔ0�g;��sD�c=m
�<ZH^=�柼�w%=;����;(��<�%=�\�;2Y�=��Y��:�G<s�;F+���>�<�	=��w��]���y0=���̄k���=u^D��qU�U�g�(�����u=N<Qn4�/�=T\=�T�x�V&=�=�R����%f��G6=��/=/x�ꖒ<I�Ļ}�;� �U���0˼M4�<��A_�;��U<Bl��hV��;�؆�j�0�yu�W=�Ӏ�)��;��s<��:='V=~�5&'=؛V�e
���=� �=�J1�j��~=���+A;�]+=\=Ż=pa<��$=�$L���<+Ț;��g<t^w��h�9v�=ȵP�L�4�K����Z����0�_*=E��b�'�6Ke�o �\T�<	�L=�R�<�ǼW����:@=_�$����<w;�eּ�`�v�<�<�RP��X�;�$4<ѡ
=�:�x>���o<�:}��Qv�2XT=����¼���<7F�m�==_�<ud��Ğ�<n��<t|7��=�<$�=nH7��2�#�c=���Dﻎ���2�<+X�<"���Y=g�-= �ѼNc�<�E"<�9����<�9b=���=��й��:=���3H���K=�6�6�O��m<Г*�s���:<�o�<k=�m<=>"2<��	=�W�d��e�W=� ;=
W��D�|�=�==z�_��h� m>=B�j=���s�=�Vj��w���:=7(�zPd=O(��]r&��_=�]=���z=������S����Dه�ye�<N���˺����<Yw�<9x=;l��K�;�;�=�T���<����I�:������E<B����<�^=8��<�.t����;kc =�2�O�;r��<J����<�K9=w�，I�<A%���A��P<�[<�m¼����k�<���<�E�yo���<B=}�\=����D��lt�1#L=�{<Lb�� =Yn ����<ߪۻΎ=i	5=�'����;R��p����n�z����Av=	�W=�Dº앻�1�;��Z��Fx<�\�<����ٛ�<s��<�d��mW��o�hXZ='�o�	��k�<PW�<�)����e�P�`����iwT��9b=��=��<�/����I�/O�}�$=3=�m���]��*=唲<J����*=K|�<�)��ü��O=M�m�`�=!����VA����_>��6��B���/��<Xq]=�=�;p�������=�ô<�����@��2M���	�f�0i=�����#=M�� <
��!=����=,�����<Ҭ����=U�:�����87;�"I��u[;c�i�A^<���7�4O��ђ<�f�<�9���[ͼ���N���=�<�������敱��������m�A<�_�P�:�3�K�=���<e
컻~�<t�<���s��Z�=��=�4i=�q���q�<�!#�[0<<t�Ǎ�����<2��<	0����<?�(�
�����1������<V޼��<��=�="M�<�����=��M����;6�=�6�F$_���E��=�]�<����y=�2=�s�EA�<�����&2���+=�j1���:O.�r�F�������I=��Y=t�6=Z���w=�2޼�.�<�B�<��{=iC=F�=��-��?:�;�к�LO=��Ѽ�6=۔=���;����9=�h�D��>%��xY<yY�����<;Cټw>��C�ގ�<T���2)=���� $=�w=�
;��=��=���<�b=��!;+<����{H$=�{
��Y8���ټM�;�Ɓ�Y>��h_=�^�2��<QiQ=�j)=�弼M��<R������y�jQ=�$���A=�{����;�}F��)=�:($?��4=f&;��^<ʚI<�U�������;�vC���=)�J�m)��⼇����<��aZ=��&�&Uc=�΂��E��>t<��-<��<s��=�B�V0��u�ް��u��4L=�������?���Ճ�W'=��Q���J�n��x-����B���B�"���<=�8��\;�5�~���=<��==l�<����6>=�u2��#R��jF��z���Ƽ���<��=��=�`�U=�<�7_=��o<yX3�{�Q��m�<{�#�4	=��=��+�l=o5=���A��<Ր&��=?�;�nk����<�D,=�+����|�ɖG������
I�;".=ӥ�<:b!=@��<e�=?�G�='A=wj=��=�������;v��L�<��;�$�.=��<�/ =���:��%��	�<S[A���;[��<�O8<��P��vy��3=?�$=��=�t�<��=u�i<?���<�:�M�<�b=x�üČ �:D
�j|���-<x�d=b	=W��o��4�< P�=wz�< ����<(�&�C�;1����=�z�;�vi�*.�=ü=M��<��s�|�8�:�|;.w�;��Ȼ����~!;��s=�S=�P����P�q��K����f<|;��q=���<X�C=9j�=;�"=e�5��?3�&@=�z#=4��8ּw$	=�$f���?����Cr�_�}<{�<���n$ۼO�&�5��<�.=~�C= G=K��;ݲ���x��/t���4������T�<R��<�#=�K.�v��;�i=OQ9��t<�u�<�d��y���m�=�)�<�#>=�m-���m=�w�;=b�<׼��x>=�4=4�Q�u;=C>=��2���:=.-,=`��<��D<�n=M߼�ԍ��n�<�F�<�fm<��-=�0ռFUԼ�Q��d;�)m�AR޼'�"�#�zsb���<�S�;���<Y,|=���<�i�<��/=2�=�z �4���]ƻ5���ɹ��"=Ҏļ�(=xڎ���c;*i=��<b��;���3ۦ<�9��Sm=�,X=�Z�l�������{��J�<Ɔ&�rE�;vO=ج6�Q�j�Jm��O3=����Ax�;0�<4)�<J�=����:<?w�eË<o�k=x5C<�/a=�p"=iXB��[\��G=�^O��jO��%=�:1=�:6Rټ�0���*�X]*=��˼�����Լy��<�8=�L=}=��ڼ�"�4=���WF��*�M=�f��=�<�>;�)�9�Z�<�Ƚ��a�<�Q�� n���Q�<)D�K�;�C*��k<�cIN��%ۼ��|<��;۵�<NG�̓<͇=l��_{�~�=}�-=���<�2�%���o=�ՙ��1�;�%�<%ݖ�Ѕ=B�<B�0�Hq=�W=~�ͼ{w$:�ې��G@���<���=V=p8�<��pq��u
:�Ȑ��QIX;��6�ּ���w�<%�V��m+��>#�v�=�{�<1�s�x�����<0�8�M��aE=.²���� 7v9�M��zH�*��<��\`=�!�<-�y�Fb���	�Z=١9=�l༿VϼIDU��L=�W=a�����ϻ$ҍ<W�8=#��=\;��<�i��`�m�O1�<��b=�S�O�r=�?�<��;I�G���*=!��p��<,���c¨�K�_��f=;�<�c�WG\=����S�<�W��W���.=;�U=ߨT��l,<�w��������ğ�<H�n�p�c�F><=|l�<Ex���:
S<��W;�󌼪�;Di=w
�<�� �-W9� �"��p����x�z��u�f����<f2���=�Ă<��N�H�<��9=y>������n,=�#�<50_<ZI���M#��{�<k4�<Y�=#�	��T=��4�.��"8�<��'<r�|�frM=CrU=|K��V�<��n��d5;�B���(=�
�܌��8=��x!H<U�_=����%�e<��<�Ɋ���D=YNr�v�L��k}����<���J�=�,<w�T=��x<>~=�W ��<�v����<I�T=.�<����}t<�
�<�BU������ 1���= �4�k��;�7�m��(��<�<6�R=霥�oj�<�z�;�s<�!�#]a</g=�XG=��g�Sֆ=�-6=xӼh+R=r�T=~H���yg�&qǼ��\�mIƼ��ϼ�N<�'.=2���%�&< =�h<v[�< ��=�iJ=�d�D��*�I<�)���L=F�c�:`�q�=NL^�ZPT��1M<��^�H�A=&9=��5�e�I���K�q=�e;�ې��q�M����<�����0��)|<z끻���<��\��c���b"�>��<&5�<�eλE4�#�#=׼ J�<c�ؼ�tt�����;a�c=���<VS�=<�3���G4j�&;=��i3=$.�<z^�Z���N�<�Q�(�(������c�;=覼��<og���;�v�=�}:~�C�&�P=!&=@=pv��s�V��=قQ=AƓ�J|b=����J'�;��=�*Ӽ�%n��?;��=z�4=�ؠ��H�>{���N<�}U���+=˷ ��k�W7s�{"o;�,���:#W��Z͛�\�+<X�;$p�:���;I{Ӽ�>��$c=*E1�|��;Zi�.�X==h�~�8=�TH�1��Vց��6���<�Yw��]��F=Y90��X����<)�F<����J��8��;�?	�P����L��a@=5�3=AZ�<�1C<T��</l�`�<�>�E����5<:;�<HR�<>�=�����[=�'d���/=�ָ��%=��߼q���qr�D�6=�&��ɠ=e￼�hZ�+" �$$����s�ҹ�;f�o���2=����"�
,���]=��;�uy=Dr}�D���EZ=~��<�v�\n�����<��_=�ϝ���(:#�<�}�;���`�.=�-<�_��23=�ռ����{<��F=�1��ۼ$�ؼT�G<,1�;-�~=�e:��e�į�<�J�Y�<��H��?N=:�L=~fW=�d=�Q[���1=��R��U	=��=ܒ���o=�
=.eS�\�b�*=��P�̞&=2g�;�@�j��<�K��w�lh�E��;.�ؼ/'=�cp���=�D*�"�m�?���һ&s���[�NC*=�һ�a�7��<��k���hq����h�5Oi��s��|�<	��<���<��<87,������W�<��'=}T&=i	=<�;?���d�;��v<k�J<RP��QVg=g}g�+j���x��(S��(Q�r�?�������@�hբ<ZO�<�h��F�<�0*;ɝں-�<����N4a�o�b�Q)���"����;kS=Q'�3Ew�!���b�^�U,�;��Q=J�u<�tb�7K�=I"d=Ǜ�<��w��@ =�l�<�5���;Ap=����oH=ɀ�<�Z=���8��Q���G;���� H=���<��	=��Y��K^<�!R���ü�ߐ�}��<��ͻ7��<amT<�tɼr���W���V�<�iż����M�<�⼠!���¼Q���'<"0޼,[��73=���<�Ϊ�s���$ͭ<���<�y;L���<鬻D�=cX:<@7)�3�=��z=�A�ٖo��Z�B�%��I=z�;�#:<tt��P-�Ղ�<�#�.�<H`�=�k=g��<��c=d��<K4p���<ӈ˼���< ^ϼq�����u���r<;��=z=&�0<���<�d<<��J�&�]=t�a��/X=M�=�pS�Q�k=���p �<���;:���xL�;�;&�L�����#�ZR=}y=>Xi�hUF=}ŻAչ�7��?v7=��=d
:D�\=L��<$����T@=e�;�>�<"��T���<U�<b���<]�L��H</�-=���E9� 5�����;� �P���_��;-��Ӌ�<�o�<!�I=�$o�hI����h�/=�F<=�e��#�l=��=�N�A=�,�*Rk���λt�����A�#$<5�u=�=%}V=Ml���"�|�S��2=w$��s�t�n=Q�o<�=.�D��(�<ʵ�;���� ���?;�+�<S
R��ּ�(�,g���
����< �=;rk�L�}=6�<K�R���~<qX���'4=i�W�=k"B��:3=:����)p�g�}<XZ0=!�/�#l��	��;a�)��0=��=�"r;�.�;*C4��¼��<��=�s=�M�����K<% ��׸ӼӦ1=T��;a�����;>�<�.Q�KF���B��Z��!�<ju ;�5=�=�d�)�5��U=���<F�,=Pd7��g�<{��<��=7�E;M��<R]�:�2�E��ACS<�r�"?=�Ǽ���h4���Ci�<�^<��Y�36����<�!�<�)���=VN�<k;O=��"�������<���x��<F��<�؉�Y�=�y�j=[+��ao"��1^�ҫ�<�2 �X�-=�t������μ�=G�}�(�q=|Y
=vf<�X|�3��i�g='c<��ּ��N�/��;|-�(��j,��"�l#E=����$T��K�<�� �ߺ�,=��Y=8�=Eg=;�<��ټ`�/���V��N<��n<��
=6�d����=��>=��=�HK=>�=�"<�(�����.]N�R,��`=���:�C��żN�<*�<e�8��� ����;���N����k"��)���Xe=�r0=Q�A�-'d���Z=#B���nͼ\U*=>@�<)� ��^�*�r�Z=���q�G=w�\�����5Q<M��3�<=h��"<M��<d�D���<��\��t�:X���P$���5=�
�<�t�<>+��_��A(�;G}�<�C���<Nt,�m�R=����Ӆ�<S6�kC���7�<H=��l<x��@y=��I=��������E=�As<Y��<�;��&s#=��=�6�jF�<:<W�@���W9�@e?<���=�;���<u�n=8g�X��<��<az�;��պ[�b<-r=qCG���4�A�q<I�'�S�RԺ�Vt<$�2<QGX=�W\=|#=Կ��M�;�ҋ���ڼ��G=yw�:�[�q�B=0>�;Aֹ���ٺ��ɼwY*���=�1;��Ｄ%=�����U<�"<3���8���T=Фɻɡ���<�뼊�a�9�=P�<<�6��=! � �m���j��;s��VE;��1<�62�+7�<9"c�m�$�gBE�u�&=
="�=��޺��6��Ko<��<����Ż�O^=��B=��==?Y��o<�7���=���<|uP��؋�W56<Y�����f=�ة<˷�<��,=,X==�r��\�5���ɼ�o�<�ִ��_���<��-=[�K�~�<?]<lr� ="=���7=9/L=�:s��  =ΤR;� a=w��<�<�wv�ߦ=u,C<�@��A4<M�{=�g�hW=�$'=ȼ�F�1=�(7��x���<ݼ9jA�B�+����<����G_R��]�T�A�+�[=�Լo
�<��u�K���a;�&O=e�����ռF�����k[�n^=�L����7=�����9��!�<?�D<���<��<{p�:j�5=��O<?,��n�#= U�<n�c�6��<�Hż�u<�7�<ggm��?=^=�r��R���6��j���e��@���Ն�!�����5�{��<�⼼��ڼ^���h7=�G�;q!l<=�B���=�E=�2;�M�����<`=�<%#�7��<m�d��ڷ�(E���z�M6�<��;��<��f;����Q�U<-�2<��P=fF=�[=��;�|���E�<<��<=;��l=L ۼ۟����Y� ��|<�-0K��:�:
û��<�����*=�og=$��;̫q<rq�<֚��$=v/Z�bH���ϵ<~�(=�W=jwӼ�l�z�.�!j=.�H9-Vz�c=ǯ�ܺ4=-`��ῼ(�����<T> �p(8��k����<�(��gY<("F=��<e:�mc9�/�N�d&=��4<v�y��o���6=|�a�I�ܻ��!=�D�<0�<�:^�`4��@PW<��7�A�O��$�ɣ)��.{��>�:"�<�b�^�����#;�(�m*%=�%=m�9��w�<ЎL�=2��Ŀ<�D7=�Q��Z:<|��,��<2��\�\=%IM=�$���<�>4�6�l�a�N=4� <j�)=���<� B���;��߼+�	=�X漘�Z�2jƼ�y��z+=��,�0;s=U�=�t��!�8�N<yR=��<������]������C���n=��<��p�<���;*2=�K!=�i=/	.=�P=@�C�;�:��<&�S��T�;턃;�Ng��q <=q;m	�<�fK��D��n�;x�
�/�0��ɢ<9(�~.B=�����_��B��+<��ͼ���ee�ͻ3,�����@=p�j�1�=@"(<�BP;�<��H�JɊ<�t���.�w_��Li9h!�<$k��c�=��L�q��.^X=�XL����<�:Y��)T=�4=q-h<�e,=W��<�7��<,�$G�<+�!����;d>�����<>��"8�H�y�*_���-�A�<4|�<�ᅼ��<\t= I��NR#��m�<��ʼ�U&�{�"=�1a�L*&=����I�<f�;9v=��=�|��`=k=һL=3`�8�<������<p�m�ǖo;aD<��=��=��$�!p�<��u=���<�x=�=���d����L=ַY<����F#r�%�7�8X�<���0h�G���:��h̲���0=�叼N=��=��=��!�j��Y- �� ���=��Լ��8=*��<��:��Dyh<>4��[��=�9��D���=UE>=b%@�gW=Si���;(�a\?=�h�<�D\=q+#=�e;�������4���,μ�|<h'�8:����`���S=�W�����=��<NL=�V�<��t=jL�@Q�<�=R�:=mF=9ļ�g�=��H<bY#=<��;�f;���<�a<�@��+��<�j&�5��o���'���z���<3�P=4�C<E`R�����Q�dF�<L-C�<�x=�F�<6n=#��<px�;$����!=���yѼ��<�^P<��E���3=5�l������{����=H��<��<&�\<�mȼ�|=��#�=80�(�\A��ʂ�+�<�
 ;��1<޿K���ۼ��!=�y=Z:��!ٻ�q!<��"� {��$>���8�_茻�Jd<��ļ��3�i���U=\�S��,3��.�;;&/<�Ň�̉-��U=o�=�//��]<�x(< Ӑ=^�=S��<���;p�;�x;	�X��ܼFrJ=��I�i<%����<�dF��:<��c���@=��9�Q���㎻�s0��_@=�� =7>���껗�2�Bw�<~z�<�=\2���<l�<�f<	�=�9�s�p��@ɺ��=���<�M�I�׼�V#�%�E�X�<�a�<=X�;��S=�\A������X���#=@�<�R�=7�D�-�l��G�%=D"�<}�|� ]K�%��<�$����<=���<�:=F6=]�E��!Y=��ж�<��k��j���R)=슺.	=!T=�ĝ��#����X=����<i)�sV�;�n��ʏ<�b�5�{�"=�&�gbO�Gi �b;;:�;!h9������[�<�J�g��<�C�:��+<���<�X,��u9�Pω�t]i=d��=�6��=l��}5��Hg�x��������nb�<��$=��@;
�<�}"=~7�<Y�7�/z��[D=�=�q=x?�<��<켡D�d�����=�'�gr=nBO=�i�"0���=��� �H=��;���2�6��Hh���2��>�4i6<�x�;jW��E�Xv
��pd<��:
=;dE=}+X�#�6��=R-/��U�b�r;��
=�w����*���O�k�i��!=�y�<y��������<@�?�7<�zR=���;��;��μ�x@�	�;N[U=�=KD�^�V<�ͧ<�s={��<�Z��m��<H	n=?�k=X�.�����
�טl��/Ҽ�B4=dp:�+~�=�V;��SL<r��<�Ks=5yT=9rt=Ւ�<]�<8`����q&�<����˻n�����u<��<#�����%;�3Q=�#�{{�;7�̻�=�?Ỷ�
�8m7<]eȼu��ݪ�o� ���/��"�<��=*�����=�(c���
=���<��<.�ܻo���8�����6=�K��l�<w#'=����}������7=W�<��%=�\ռ�a=�hx;��r�yؼ�~.=��6׌<c:g;#����`\��/��Y�_��C���G�;p���ڻc�ͼ�Ee=�{��̶�T8�<�(������}��>?�5G!��Hм�F�<f�&�Gʏ=��.��ɻg}������~�<����6K>=|�\=�M <�~e��[�]��<��;y�	<�z;�ϥ<���kC�;A=��<��;ߺ����E�e9�<d��;��T�^�$=O����$<�M=�?�sζ�=�����~t�:�1=�J��W��=����5h�;�n=��#=�G�< �R��n+<���<~j�<��U��7�<'�l��bۼ�/=�-�<��</A=4:2=8E(:���������<C*n=�D=9�&ߺ<�\��v�<�Y�<ilJ���%1?=h5���=�D$���<��=B:=�<���<q�E���@=%P�<���_��<�U=v)`=_=l�O�r�Լ	�ʶ�d#��p;28O=� ˻S+<��}ļ�գ�h-J�h;��:[�9I��<;���y�,��X<�E�<�K��%�=�&;���<!�<"�=)L�;w><�p��7���<0�=����! =9��O}p����N�<��G<�*�<ۻ��:�i�� h��P�L�<=tc�민X�k=V�r���������.�g�0=��(� m=�ɹ<��oqW=�?<�oM=��:q�'��\=�ud��z�:HF��h�3w�=�q߼$�;�ƼSu1<�NA=� ���6=��_�+W/���N��K���<�& ����;��=�$=Ѧ_���@�	��<�N.�������<��`���B�V��9}�;��y���<�[��������Զ�.4=�V�.X#=�6<��a<�:=�`0��Z���۽��4�d�>�R�?=�,��"V�S�)�(U�;�A��E�"���;���<�"=�H���ݿ;?t7<�L=��=���c��J���P=}S<ӻ�3=���5���<I�1����ɻB-=�RüN�6:�8�62M=��}T༂���#Ȼ��>�D�����"���O��5�8Ca7���L��V��!=�o��fI*<�.1=�a�����o=��<�<��p=�M��L"<��";)V;�$=<`�u=E<T=�����<�&0<s�@�5��;L�������6`��nF=�n*�N¼T�=�H����h�V���0%�q�q<�U�<w��������2<��-=1Y;�D���(�97;x��5����=��&��Z��#~��2�;��ļu��<��<�H=|�=D.��|���Wc�;�����<>�;q��S��Ѹ<=�)����<�E!=-�F��v@=��*�o�=P,��ȃ:��4=vEj��Lb���[=G�����:�;�<9����?T<�7���� =c� ��t2=(�;�
4�^=�=2a=�:�<���!=F2=`��<����`ż�M=Is;)'6=)5����� ���F�y�x;e
=tn=�\���Q�j�:;�缝�b��z=_����y��J�ڨ�����vy=A+5�p*7���<�n&="��5��9 ���s�Η.=�[S<=P:���*=@�+<��-�p�P����δl=��<��ټ_���e�r&���=��<.�N�)=}B�׃=��h<���<�TL���=J{<���V�+=���C?=�f���1=��;N�l����y�;��;{-=ye�Du��х=�LS<����(=�,�;�M%=��-<�)�<O���C���c<R�<��~<5�+=ϗl=��=4�<�#<"�1:̉�<4 =�T
;7=�a=�#w�B�<�!�?�=l��C�)����>�<�g���a�<ev����w������<���L�f=���<d�F�h���B=��:<�������=�p<ovݼ �A��ύ�R?\=&�F���b�m�1=ܐ����������4�<1Ki;tf.��>�Q�r<H����}K������X{��,>=��L<���?b	��5�4h���_=�Q;��f��ᮼ��9Z�<�V��f��4��ۚ�䳀���{�Nc�<h漓�!�Okp<S��3<v��<�R<g�����<مƼr~,�#O=��T��l=��e=��=�ּg������G���<�-H:��<���<�6���u=)v����8= �t���Ϋd����F4=�Hm��W;��=����3���_=�A�rt̼:_���W�<�u�;m�6g��'Q��|f=;
�<C���̐J=��W=��-��[��;��_�1=�^�%���)�gt�ߒ�<�6/�R������:I��"v�V ��s�<��M=:�X�s��<E��n`��y����;e�=�n<�b����<�<��=Ӗ˼�ղ;uq�<���p�;y�<q�5�E���=<�9�k1���(k���d<mM��'��;]I��^��B�:��.=I_λ���<�����J��|�<��S=������:=uL�<*%J�l =��B=���y���㼖7�0�e=a��P��<_��<��j<�=����+Z=䠬;���<y�=״B��*<��5=�h��mz)�=���M7�<l�H�GJ��E#�KbN=��';�S=.i(��F��_69����<������X��ڼu�d=� ;V�[<]�����8=P4,=*�P��l�<�ȴ<���`�F�4Ő���f=�B@�G�h�1:�;X��z���+��<�v��m�<�[�$N��ּ�3�l��<�o��t���d���j=�����3=j=������<�X����%��j�����U<yѻ�v;�Z��"�<���A˯<c(�; h�7�"����<�wݻ�̻��?=�Np��}?=xl<�0�^8����;Ң���@���D�����g��j�#�R�l�6i���gd����<2�2=wM�= N���<e��:3�E=|��<�_��x�<��B���8���$X!�P���#i=�2-��L��RW=LZ�<���<�k�<�H`=Ի1�C�y<�,�;DI&���8=�	���̓��y�<i�#��@	=ЌX=B5U=2�k���,=�\�<G���>=��օ={K�<�ȃ<��ܺ<�ǽ���=��U=�ӕ<9�<��<���&�C=Wo�<8�h�|���_=,��v���	�ٻ侩<��h�.�����;#i=��= �H=�!�<���B�⼎�E=k&�;L�C��� ;ٱA=���
r�{�;�=�jV;@s=�6�<�[=s�����Ƽ5�<�]��~�<�UJ�ro>=�C?=���<�¼�t:=���<Q��_ڼ�y��,(=��$<_dؼf]�<�k��ĩ�<�,��L/���b=��<��2��t�<JS=E6�<w0<�����'�Y�a��n���=�t�<c�c�P�;Wca=��(�Ń%��ϐ��y;=�=�;7�c��(�;F)���=L�S��<�`X=&=&�8�"m;�13�<Q�^<V� =BEd��`�ٳ�</o�ԏW���G=�N=j��)hd�^V#<��Y=����t=K0��}D��y)�g���*�<J\[�iz�������L���r��iG�/X��d+=O�]�S�����󻺿k<�^9<�5�E#b�d<��G$�iUͻ+�u��,3=cd�������{���!%��x,=��k�<���;u=�<�m���;gg�a�n^=�,2�.���Լ(��<-=�ކ<*�F�B�[��-�;�z��I��y�	���	<`R�x�J��ڃ=�7����<�}��J��<�R��i��<^���QF����5fq���o��w}<�SȺ�X�M�o���=9 :��<�|=�卼��H��;�s�<�!P�i�� �;7p��(�v~=�`��<9����sg������$.��
�B�"=~�Þ�:�bL= ���4(=� C�z�E<8HA��L�<��%��+[<�p/��i!�=���R��<ۻy�A߽:�u��6?<5�$=�o=7�	��"�N��4N.�- s=�;y�м2Ak<h#T�JJ���=S�%=	2�</�<�Q3=�0h��7�<�[u��~o<I6��ǅz����<�C=8I�`0/=#�=z-�;��!���,�G��:�!f=?*�U=e<�>�<�nb�au!=�L�ϐ����$�;����)�fÖ�ߏ?=���<Lv��w�D=E$=G �<=|m7=L�<��ļ�p�<�\��:޼����� =)^]����R�<t6v<�- �qZ9��<��=��ຐ4=��+=M!=�C=�F5=�t��S�����Ny��y��?i�g�B���F�"=���\ڶ<�=j9�%�=�ݣ��:���u��F�<��=��]��^@=QM=rn<KB=~�#���P��tS@��W���<a�=����W%<n/�6~xY�~���^��<�(o�epu�k�K=�k�<���<�S>�4���΋=����tYڼ�] �Qjs�j	���N��$�il5=?d=��=Er=��;�㼲�;�t����]�P=_�=K�o<�7�</����#܋���<=��<��@=�L|<yn=�4}��ET;te �Q�<���=B9$��t#�3CD=��ۼ��V=���&౻r�G<�[5���̺�़wI%�l��<�+�=d�=�e��x.�Ƽm=�=�q=R3�<�zɼ�0���!��<{��<W^7=���P���<�A�V[V=!�Z��!�<�w)=���?>���l�u��h	���<���Ɩ�<j�<X���Ct=��#=��3=�V(=FcO�i�&�ε�<_x!��=��q���ڻ�=iS7����t<��M�U@���==z���?���|�<<L=�o
���<û���
<��o<��=����T��GI�<C�˼,��<W8k=����d=7fG�m��a0�j���-YS=^�Y=��=�N=��=u��<l��<U� �M��<�,�<�=o*Ӽ8�n���=*u;�;=�����<��%�;F"=��<�%]�O�4�v�<��d=�y!=oC<2� =��:����<��<W�=��T=i������a➼9��@y���㼖��1�Y�(���Ht�=9؉�M6]<���o9�<�C'��mǼ\�]�9�=�V=HMD���<�*==�=�ke=�CߺN�D=z�d=8[1=$=��g�:fq��9۩<SE=Dq��~����;��x5��и���G#��(#�L�t<
�n�q=��Z=�K�!؀���d����<��_�+�f��_V����;��<�2=��0��=�=*�x��(���G�a=�$A=�������8M�h;:%	�W.��м
�Xn*��:�y�H���!���\<˞k;���X =�X����<�=�K=�za=�b9�(���ʼ�7=n�]�El<&G�=|O���j�?$����1�1:!=r�⼩�Z=",��C>j��;����뼪�<L,1=vQ˺��x�J=O�u=i��:i�=>����G�3��G2���<
�=yW��1޼�u��:�<��<�,&=_B:�6Ǽ$=uh»�c�;��ݻ�V�=xj2��=�uR=R�<v�ƼLj<=�w<��_=������6=y}k�$�G=��<B�o=��:<]9<��=*�7=)3?=�n�<D�m=e�<WϦ<�k<8<�T!��$���V;-d�<���;����:��~
=2J;ԋ	=��3��U�<_�n<��<�"�=HH:��A=H��<�i�<�������5J�z�<�_K��.�b&5�t�<�s1=�iR<�2����=�<Y=�[�<�q<�a�<���<�Y=D�B���;��$G���Q��U�<w�h=�Ԇ<�T=ѯ�2�,�<b���U<zD�<�2y=�`h=��)=<�w��Fg=���<�\(=K�N�ڣ��2[�<ʋ�l��<�R�0ϻ����׎<
��2����O�<__Y;�=Q͹�P��w��-��/�=��<��h=+!��H�=@ù<ش<�!=q���
�7�@��WU#��d�<*�<����K������^=GQK��	��7�<5n)��1/��D��NH�Q�<��~=*��^�]=��m������r<��<��`=�L2;FB���B���{�qZ<�5����/;�K��	��*����Gb��R�;n�C<�"�"#]<�`:� = S���2=&�=��<�^n�<����o��<0�=�h�;�
,�B*�ro�@Hy��M=t�5��u �NC=�Z�<(Wl=�=��]=��q:G/���<�E����<�	�<��=
�7=��r��^��ь���<�kڼ��A�F�μ�K��*�D=6uԻ �-�j�̼Y���nY�/�~=�?q�E���*=��=�:�<�WH=M�o9���=l�<xf�x�=�.��*���l"<w���R����u��<�=&�;(ia=��$=O�J!�<�$=[cɼ4�}��Iؼ�c�<�譼2 ���<f}��r=L`���tl� �?��H�<N¦<�9=�'Q�oQG�����m�<�XԻ�=���=-a;<D���i=��!��z=N�=�ļH��X��<��j<�Q�<��=$�;J=E"8=[�<�2="�<�+���\�<K�¼1>�;�]#��0=�>�<�`�X�$<�
�C߿<�μ�';'���*�َ����<0�7�DK=�=⼠�=�%=��A�	�%�5�L<P"=�Q�;e�Ǻ�74�r�F=�;�pO==���{"f=�G8�Ox��	ǼG�2���=�hh�+t�=���<$>ļ���i�K=��=�ﻃ<�D=L6��C�\���^��ɻD\]=J�"=�u=I�3���缵'@���C����;bl'=�O�<��<�LE=��8<�R<�=hz;�L�<]�;�?����?�s��A��;��ຆΒ<ϳ=������L�=<�ᾇ<���l�-=C�5�ڃ>�� 7�0�6=�~=���\==W������އ�����5W�L�������X���<��<�I�ܱ</J��=�*���$��-N=TP�_w�<f��:S�>=3��<oz8=�.�,I��c�W=�2<्<u�ϼ�Â<�m�FD*������<(����u�E�=��<��y���H=�A�<�=X;B<�(м�M<[���V�=t�I=�� <�c]�< %��ZC<�P=��J*<�{������O�+�8��Q��x��<�Q_=��[���U�|�k<��*=�r-�Z$=]:��K��|8�2�<�=��|k�(�*=���<�¼�g==}tP���<�̼���<���;�"6=M6	=�`H�';P�C=�Gw<:5;=�:U=�]�Nۖ�Y�;Hv.=��3�x=��q��y'=.�n=i���� =V�=�u���<�<n=<�c��xDӻ���<�  � �h��쀽MF<��oY=b�Z���ʻ�6����<#��;����!	<�f�*D�k�Fy�;ͫ�W�w���ѻ�o���ּ�� ��(�A�?=�5���-
=������<t{�<v�=�� =��'��|��<��=�<b�<��=�L%����<�S$�p���&Ӽ�����񖼜f:�ʊ=MKJ��z-�3���gP���";��!<�$\=�p¼@�Z=x�<�(<&�9֪=|5c�]Y<V�<��=),5=��μc�W=J�=�)3=}S��޻?�Ƽ�Η��y5����p=3E=`><�,�D�"=6��<97�$�<"n+�M�=�{�em�<:�)=r'<� ���1=+�)���<	�<�C�<�p��Id��7��<߷d==��<&Z<&_���8=�/)�8�R=�j��G�=�=�;����x=rD��S>=��I� �6����C(��I=03=�!=�W^=6��<�7����,=�����E��<��ۼ��S=�?��p;��=[�����|;=E�!�����O6=<� �9��!�:�D)��L��y9<C�2�����b�;��D=v�(;��<�^<�A鼆a���,�J
ʻ&U$�3=q�|<�X�\ͱ<����-��Jf�<%�]�h�W=��0</��<�%B=YS��Q<=�cx�!����7:��<�3	Y=a�<Z���z�=kZ�<�o���I=�UQ<=�����;���k:)��2=��V��=K=��)�N�<�q@��I�<L3�;��-=��`��k�n(	=�-�<lS�<������Ἷ3=P^����}�.�̅L��[;�N�J��x;���4�� ��`�Gd�<���;�a�<�S=��<�FT���߼Ee�<��~�k@�<�qh=�������F��;�f=�Ԧ���3�SU`�{i�<��{=3d*<�E-�.~���j�KC�<L�n<������<��>=� �<qR���:��	��u��5'���|V�K>�bc]�J���t:��>��&�=`J�<1O�=j�;O���y�ȼ!�.<��+=�U:m����;(U=�R=t�=�������C��Nu����<�Qt��"<y��<�D=K	����
<'��9/ %<�eӼ�)��J�<s)N=�a��ӓ�;ɸ�<e�=S�1��o�<(�N� J���"�<���<���<�Lȼ�,a�a�;��e�<�0޼�0���o�z�=0� ��D<X6Q�_k&=�1�-ӼJ��;�rY��R�<��+�m%�!=Bi�����鼞<{
=�CR=���=��;��^=D^��MH��ٓ<���;�輼�W��dV�z�4��� =}yo=�f�<��<O�<���?g�:xKL=C�G���ؼ0�<�@v<�֞������=��<�(ʼe-`=�Ӽ�H��<�|P=��l������	+�0�?=mx=�a<��<�4=k�G=�����N0��C��n��#=ƚg=3�=6��C<�?���I=���<*<�;��a�e����<L>;��=X���Z�����J�:=s�fw�;n��;�4��<�.���=Ҽ^	=�.Ѽ��O����;��\�E��-��;�����&;��̼�Z=��v�Kc=�
�ֹ<��>��<�_͸0a��V&���;=��e=	�V��ͻ��}�;�ό���	�k�_<7��<o���sa=�h<�����1�6�=z�=2A;��=���=����Y<mC����<t�E��e��|ȼ膞��d�;"�2��m(���<��M�b0�<��$�a=Su�_�����W���=*�����)�~�<CAQ�Ĝ��O����T=�(������<'�A=��λ��0��:�<k�7���s�g��<n�G�Ē����c=����m�S�����i��Ѽ�A]��vż><B:C==�ȼLF�<x��2<-|�:�n��i�2���,=2�=cX��Y��mR�_K��hd&�v���Y��E4=����ua<�e"<�d,=��Z��7��'$=��%9wQ���5��Z�<a^�<��R��:��f=��"�"��=�e���A�F�U��<�;3<�=5�#�;K�=��=iF���q;��Z��;98�;�K�q�=8fZ=��O���c=�=态�'F�<�Gb<�I0� �j�a-t<�u��8*�\�'��|�<�/��O=v$�<xy<a�=J�	= �u����<���׃<˲<�}�F�;H)N=��ļ��<�01=(��<�M=�@.�&~��H<=�ZD=3a����~���A��}��;���<s<=s6=T�Q=��0=�`=t�c�z�ڼT���O�{=߼�<Տ�I�5;�����;�̼�
<J��?;�B��<}a4=�D=�Lo�Nc'��#=�<[��2�����"��Y[<��n���x<��6=��b�h�������<s�[��cj=+�;�л?Y��7�\�xT�=��e<<��;�H������n�H�y#D�6�>=4>=mY�<�T=��u=?7���=_�P�>_<����0��<�e�;[�d=>�'��u<*�o�i�o�<w4:��)<(%<僚<DU������
+=���<��E��eo�+D�$X׼��=��^=�p�08��57=�0�����=(?�I�L�m�=v���4�3.:y
==e��>�^;l=&��ܱ�& �<�S������<�kL�h��=�%<Q�r=����ܼ�ֽ<��p�ۀ�<��&��_��9�=�:ự�#���1��D�3���=os��䫼��q=Q�=�A><�wh���p��W�<���<�P;�G=�$�Wf��f��;��o=��}�d���Q����n��/}�IF���>�Eμ�7U=�!=?<��<:�0=���H�W��g�M�=����e=�w<���<�C�:��E�U�<�L=B�2=��j���N��Q+���!�_2<?b<:`�<�s_=C^H��8��(�<\!��o(�e|�քѼ	c"=�A=���:��<��<�
l���m=�C=�n)=29�<E�<|�o=�G=����l�<f��;>��>�)<pbr;I��u.=�{n��OR���<��n<�����	=�8*=��6�x/ʼ��3�H]�����;��'��5E��A�=<	�==tS���7�6���Uռ$3�<Ҿ߻;��M�$=���~7=�M�;cM*=Z�'�o�1�u?�<~��â�<PT�<�̡��~a��頼/�=世���#���<���<�;���z�,<�}
;ʯ�<��׼39=���<jR�<����F0�X�>�=P,�<&s`=D9�;'�G=?;R=L=�n8=��	�]�= ��;Q`м#w=�Q��y�;���<�ܡ<�i{��
�|��E�s��̶�U&ܻc�<ˮ߼���O�;@����[J��ۏ���ټ���T(i��=�O*=I��<���P����=I��$�
=ń<��Ǜ�<y�$�o����<��lj=�z�;�_9=�k=&�<I_E��R=3�编-��e{��+�;�R�;�#�U��<%\)=2V���Y{�����_�?��;ג=�g=��<6��J�j=e�=�)Q=���|�K=*CU<ݨe=ФG��2b=��`=5�+�(�<U��<R��*�G��G=`%�A�=��<�h=��Y:�t�<�o�V<��Z�1Z2��}K��ؼ{�X��{@���z��zN����:n"V<Ƴ�<��v<���;�NübY$�8HG=+e
��6��rs�?��`yf��]�<S�7<:v�<���8=Q|/���6�<�[��Va�S==F��;�?<']m<K�<�j�<=���*��f�%���=�ԕ:�Mb� |���<+�o<�t�<6�ڼ4C	�����֬�<��^E�<u)d<c��<5V��`<.wV���v=�0J=���qu=)�<�Y빊�c���j<�S<PWݼ�3=r�����;Jk��,��F~�s��x<_'����7=8���<_�=�P�#�n<K�<D,�dJi�U�=Ƭq�GB=6üH�
:#HG���&<�[=���<d?W=��;��d=N=<%�;�<�$<�,B����<.H��
c=��8��V%<@=��{�m#��'��<�,�]��c`�a���`Ǽ�qn����<A�ɼ��D���S<\g!={Ӟ<	�3��<�?3�SO=})=�,�<�����m|� /h�Ezy=�t=S���$=�㩼g�<@6�SL�V�j=�y<V=�c;���Kމ�*:Y<�9��s���<tm�?��n%ϼ�;�<%Y��2*�<�:��P��j�[�<Qd2������u�z��<���S=3㿼�,�<�tA�(��<�JG�'y�<��'�;��	��e��p�=�4�0�N����<Z�h<�����ң<~oS�t�<=����Y <f�%=�2��	�.�<"��;:E�LS4�T��<,�C=��!=�$y<@p=Ŏw=��+=UW��r��w���n���̏�= �X=C����Ƽ�=���<q�	=�MƼ��=�	�=�XG�P�ʼ��=�� <�F��������ϳv=��`=%�k=O{+�t|ż\�׻�#�����Sq��)?=w,�Q5(��P���=���<�j=��O=o�{�=|���,�$�Y�
��~	��+�<�B=J�r=5Q�-D���r<9tѼ�R��� 7�艎�$m����=�D=��k�ks=N<-?,���!=s�<�0�<��P=e�&�o�輌ኼ�@���N��(�<��=�12���^��8�<e�K=z�����ULc=p^ �����<8N��[�A=��N�̼ۘ7�<�5n=�5��w�Q;��8�*W]�X�y=D��E�H��hj=��;�>��;A����B��=,Q�c���b�D<���ש���:=��R�㧔�	b(�CNѼ�_=��!<��U+�<�`���<��D=<`�<{��<��%�OE�e���9='+�]V���.�O��ux�oI�3�=�����<@29=>����H�=����+��`=��k�Exg=���{8=0�]<�,�=Lj=��:�@'=l@�ZX�<A�L��0=���;�"�<3V:��*[��d��to��B���[��E\F;ު5����<�4����<@��<�}�0WZ<gʨ���:�e@�<iJ��(���U=�2<(E��-<��==���<�7����0�m����M�<5vD�ΛH���=��"���Y�h�ռt[@=�I�����f�= �:�bB��&?�
��;~Ƿ��c%��e��1�<fO��5���O=-��<�*<����%K�<�Z3=��={�F<�'=��?�o�6!=��<�׺R�
;�v;�[ۼ�O��A=x�;x�`gA���"=a*= ��S�<�4;d�e=vs��<2�&��3�'�[��N=ؚi=�������<�l6�=ZE�������=9�(���/=2ύ� �A=�Dۻ+K"=�iG�3q =Y{<�=��S=�#����<��"�)�H�L�<���mn5=<�s�>I=:�<D6Z<������9[��o0=ߎ1����;��^<7V���:�=�`=��=�=����B��;0˴<��?����"�A����=�/�x��<fVd���z<�a�<�v?=߳<�]x��Q=�� �:�L,��{3=j܂���=&s|=`��f˛�N~�<$)�<t �;ٺ$=uj�<��k1���J�g�=�sd=�/?=�*�2X:�VR=ME�g��<P|��=�w;꿖��U=R��<�;��y�/=Rzh;e�;y�.=��%��=FX�<�W��$�'�x<���:�^3�;�T=36=�I�=�O����:����6����y=�@Ҽj��{�<rO=�>�	���-���_����O��`舼e4:=Z,:�T�<HI%=<v����<�f��]�� W�;�^�<�RJ��=P6<F�o��?��>�<!�<�"꼍��;�ٹ:�\�ɨ�=ֺ<�<��<�80������C'<��ʼ��4��,=E�2�sG7�d4<��<#�<%p���!�H�ռ8>�!��.b5=�2j�~�ټ�-����9�)u9�aé<s�n��:û~FS=A�<I+�<W��<�m�@�X={��>��<�q������]���X��!R�H�,=]�𼓷B����}��n�=l�<�>���J���;=��H������y�=�g�<"gK�Ss�Yѵ;D�e���0��Z��֢�< )=5��;Y��8������v=�=I�<6�|���*���w��<���'�Ճ<��պ*�d=�*=~\=z9=�s=�0==�P|=>�==e,=��2���x<㈘���b;_Jy�P
=N�=���<�G������=9�:���=�<���<������<�X�<�����=$�_�<[=��<Wf2=�Q<�Oܼ�XһDi�����\)��`�;���=��D�O7���=���U�@;h^�<b:<�BD�ճ�Zo&��6`=7�?�)u �>�8���D=	�)<���<m��<���=�Wv��A�;rq=��N<�=k��;�<n�ȼ���qKW���;=�6=���;��F<���<��=Y���p��=TV~���=f�T��<<����o�;�}Y��`=bj�ӹ��餇�YF����<�l/=N��<�K�N,������<��=ëL��qa��H��&6�"�7=��#=y�Rּ��<�|�<�%����q=��ȼ� =2o���f+��{L���ü��)�YB�:8V=���<Z$\=v�<��λ�TM�f�B=ZO<�Q4��Zt=��D=H�(=�} �,a<��<`��
`������0��vS/�Y0A=x1���X=2(M���x��A6���L��]��S�n��b�4�#;,e+�ק@=p��Ǫ�_�|�$���>μ�K[:3=�f��\W��mԼ�We�bV=��@=A�(�B�1�Ց)�B���Wm��=���:�t���9=��⼑�ۼZ7 ���/�{�/==D�	=�.�3�a=�60=�^��B�=r��F<rr��;�����d���<rLq��=[�چN�؞=��*�	�{=z�t�3�׻���<۸#<�T6=��e=&�~���W=�������'<=�G�9P$��Om}�����&�q<���:�� =��_��c��2��
=!�D�吓��}��ͼ����0U<BT=��<�7<�2���N'�3pQ=�E�<��=��g)=���<�x;�U�<�ػ�z��Yf�<�.��81;jI==Ю)�;�,<v�.�@����X�:�B��`^;�tc=ZZv<`��<;�<�=����<�	�҈=}��<���<��b��<�q�;u�8׼�څ�Ū���;�/�_�_;�?���t��'J<v�;�^�[[G=�4=�
=/=k��<�Ge���E��M-=�G@<��=�%���3<�N���$H�2��L��&�;G�=�T:-s.�*��<(*=�EU� y;�i�<��������r�<�rt����;[|���w<�<�����m�� � >����ܼ�9=�3��޲�{��;�vN��=B>O=��<�C���2����1�tVn<� =b<&�=�>=�ZE=k�<�^��?�K��N%=Q�<�?=�I���Z���lͼ�<�y=φ�;�S¼��;^؍��5����;��t=�H<�8b=�9O=zl�<Qv)=��j=[@�<��	����  ��%	��s�=+6������p:��j�{�{h7=,�H���=8�=T<�<��l�F�k<ހ��޳9�z�	ỻZ<=�=F��A�/�����E�g� �#O��1,m;V=�=/=�Z<ѵm� ��<@��<�[�<G �<��v��M��(4�	�K��(/=b�"=�s�<�u�<#AV�s�k��� ���<����^=��a;-�Q=�a����<é+=5`K=�<0<���<h:3��<��<�ӑ�y#"��e�;�����$����;�=b5��0c�W6�<xڐ<�4���*=Z �a܍���=� =�B�<P�I��W=X�� ��!E@��c�<�3�������/K=��&=��<�Ua=�?^=�0=c�<R�M����^�(p=>�H=x���T�O9�i<#N=���������==�0�=��㼅B=!��<��4��UI��&�7g��;���� �=9M���Ҽ�|һ��ȼ�N�1�	=Wn�<r;|<3%F���n=?��_��	����=�J���u=`���=:=w�,<�P�<�rF�)��k:��N���2<�ȼs<��@<村<�)�;�F����&t<�Zʼs=����;�<��1<K�=�xZ<�zT=(J�)�����<ůK;�8#=|�Ѻ�,�-Լ?��c�;X�"y����)=3}��86��=��0�����0����&�����U=dP=���}=��;������
�0>��p�l��� �H��<�ƃ��`=����"E=��A<�j=�T�<D=��:XV;k���꽺�F;�����X͡=Mn1�;A}=�R$���	=c[=%S==(a=�{�<�b9=���i&�;�+�8�L�g�<�<�P8:���<�d���<��@�2/==�"м=�U��eڼ3a��>�<�m;��*�5z��	x�<��2=�!�;�-=��<K�p��U=[#�<v葼0����ռj���"�#=6Lw�Y�o<`kT=ɣ<�����9����>��;˪h�A�e=	��<_/��W=�S;�,����=� ���O�<k}#���<��=Т�<�.=��X��1W=e�!�H�d=�Z�hdA=�ՠ<�n���n�,�=��ܼ�=@oQ=�|����=@=_���5�:����܀�Z��<{��z��=�L=��}�m�溆�Q��u3=�s���q>��Wμ
l=B�N�#-<��n�F!*=y�E=SNJ�K濼>�=I�K�������<�;=+�=���|�;�$�b�}� �#��I�<�q��:[<�U(��S:g?���4=�K��./�;*+�<��X��Hۻ[� =9$�� �'�~�'<`�'�]�_��S~<r�<�"{�;����8K=-��<��+=lN�<\;����.=���<��<��<�	�s*e=���<�5�z&�;"-<����\<$a<<e=%�5<��D=~n���=`b=,N�<�0ȼhļ�=gY�E/@�%�=�1f=�0��X�n<��<ԩ�<{����L�<NaY=�{;]!=ܞ�<�!*=is#���p�<90=�<
��:d�f=�G���<�S=���<��g= ;��F�}�;�a�|�)����<(Rͼ]�(<��;�F���V<)�;� Y<�:��n+=�E��ŭ�:f�E��"���%=�7����&�q�<kkD�cx�;�Yp=�C�=<l�s�=O 7=�.=QW��O@=�q��r��@��<!�Q��='�����<��-=>]��a�gN=��n=�����Ļ�`�<oz-����a(<�2�2�]��/7=t$��Y�=�=�<9d��fF�<��}����(�<�O:<��Z<Y����<H�����p�ږ=�m={�<��켈#�����;@{E=�&=
e�<KP��z;��	�w�ۺ��<k�j��%��T����U=E�=�A ��j
<�[ӼL�B�Qʳ<*��<�<��=@&�<^�W�q�;�[�;6�0={k���a�ׂ��!���3����Mv����;��aἥ�����.��;_<�?=o64�g�=��<��z��rZ=�^D��=/��D=�R<��X=|@�<R� 6:I-�=)�=%S=H�,=F�!�=</y=^G=*���ߺ<��=Fdu�X�A=كU�8b�49O=X�&�z�D{�����<�����<���;�k�:��e=ոH�e�T=�����C���ż�G��*c�<VL���|<��=t;;T�1<S�';�� =�s��vO=�j{=n��<��٦���2�<�k(���=���/=�<ok=h�󻀐[=ҏ�<�� ��N�<|�<l�A���_��E<�	���tM=C4��?m��!3=��h�H<֭ۻf�¼�&k=#��<a��<yLO�k�m�^JC=�N=��<I�Q�p[�;�\�;�s#��/k=�EV=tO=��6U=߯T=��<��c��jϺ�	�+��<��=Jh��r'7���<��<�)�<h�<K�:�:=_��<aN=��P�i�g���?=p_<䕅��� ��F���I<V&���L�No=	u���j���1=��<���=�S�w�w=?CP=J���i�<�oD�сq�=�C=g��y>;�*N<�6��h�4<��o<��=����z
<�����C�Ԑ�;�D�}���=�B�4�<%�<��l�Q����<}���z�<�?g�<=�=36W�?�<wp<�X=���������{���<C=%%6=�7�<I�3=�[�Lm�D���D=%x5=����6�<����j�:�F�!�o{��V��$Ƽ��=�	��J0<��<�P=����i`���=G�����<�e%�����J�=�@�;����;<�I�7=�vP<�w�R��;2��<�:����K���ܼ�n��2��;jR=>�<J
�<��
<p���6L����޼=�1���߼�9<5���a%=^�=<�<��D�U��2�<��~=�m*=H�B<X�4��2w��3�<'a��L�<��0=0��<�:�y/�Q�t<H
:�7�������ўӻ����6<���X�H:�[&����:���<?�;]8�<h��<�Ί���E=0T�����<�3��G;;d<j�N;��r<�0=��O= �@�px��7ǋ<��*��<�<B�N<�9�<*ٗ��Q��c =�~�\�<�w��W&�<�<����4Q=:�u�f�=��/�@���wo�<z;;=|�G�Us��ؽ����菶<�:�����:ͼ�'S��<[c� �<�<���r��}�@�N�W��<%��<�R^�G��H="�?���q�(y�:���<�)ջ[�(��gI��=�`��x����=�t�<g� ;+��h$;�4 �������`=�*H�F̼�ټ'7=��;j3a�#|��(�W��<��=�����C=���<9C=7�j=�G�<K�=�=H�@���	�z��:�=�O��L�='"1=]-=|:=���:㴼!a*:����s<�G=ti#��[�"���f�<��X���</C�<����'�<­�<,��=�&�����fк��H=cyϺ
M��(�<�2�<��o=%����pp<Oc�<6D&�ψK�L
@�
9�;�ֽ<=(��<JH���A�<���dK�<��f�g؃�F�J:D=�)��"�<ێ*���=a4�<\o�<w�=Kv>�h9,=��;S��<��<�
=CZ:��=�Ɓ=`��<8�<�7��]]=�f��W�;ɘ�<��9]��>����<�����k߻Y�~=a�;�-+��`��A=��4�L��<4޲�p�ּ4mX<�I��9!=�b��,̼���;�=F<7�|7�<���8X=Q]|<�K4=����];i8\��d�8V<]�=�=-l�;�O�U�<C�<	P�<Dp��&7�=B�9�9=�j:=AB=�����=el_���+=�$=��]=o(v=%� ���4=�LX=!j�'����X��=���F='��7̼U|z<|5�=��L<7�H;��<���*����>�ި��T+=��������"j<��Y�`�O=��Ҽ]'U=�&D=�e���(7=�p<�,�:�	/=F�4=�<����PU���?=��<��s�MF=(k��i�=���	h<�oK��^\<:��;�| =KK$�Ǭb���Ѽl�%=�kh�"�,�]�G���ټ��=F���v��1����D=._<��:=
#=���<�%'���Ǽu �<t�<�=���<$"@�������������
��Cp=���<w��<w�A�\��;��\���:<��=6U5��[����t�C$�U�?=֫����|e�:"2�T�X=e��:U��j"�)�c=��<x;`�4ۼM=��G;�� �}�3=�k=A�<���C=e���]����&���=g�!=r��<��̻���`�<��Z��"0��2W=+���&=)N(���X=�b���>,���7��P�q<L?4�Z��d$����}:{�ݻ�Gl���=mμ��^��ռ�և=}$�<Y��<̂<�x'�-ƚ�k+<��L�,�E�2�;�Fݻ��F<�T=�s��C:=~�S���l�g��E]��"����*Q��T=[Pu=컻���=��1=��J=}�[=y�=U�<[��&�p�<YPI�����'�Ӻ�缀Q��G�<I�;]L�H�!����<'N���k=��<�����2�c=��`==�S<xؼ���2�2�qR�<Q�q<�L��=�!��h=��G=}[��I�<,;?>���7��);��8=tr�V�]=�7.=�?���#>=H�$=X9=����������=��<�=9;�<��\�?�nH=q��������ͼ]������<T�<{F#�hy�<n�e=���d�m�.=�v�%^���=��=�6�<�;=�9�<����B3<ͫ�<�.�<	+���?���*����<kyJ<o�e�~�;�K�^=}�=�i=�a��F�;��<�Gɼ͇�h���~
D;�0K;ޠ��n�<���� E���2����<ߩ=mC5=����h�$�>=ތ�����7=Tj.���<%yf=3!�;���.z=�c=��C��9�<����⸼90=O�=Q��;��p�$���� ���%���O���C<Ī���Z<�T=���b~���p=����f<���;j�=Y���׊��eI�=�D=����ߒ����U�v�=ƅ�M�����<N>'����<�Lмz(�:��%==�ټ��e=��B=^�ٻa=o!=h���L��Fμ�Ϝ��8f�ԙ�����<��5<�Fa��OZ=�۴<@X:�ۛ3�hc�<�3(���W= �u�Q߼yv��Ԛ<NB�<�t!�������|�LeE=�=4=1N<�Ǎ<x��<��;^4C��Y����U<Ӧ�<��4=�L�<-�Y=a�ߺMS6��w��R�]�Q!�<��<:��<�,�<��=t�@=�e���i ��/B=���+\=�-�<��׼qP<��7�2?�'%�od�$��=<�y<� =(�:� B�
��.�<w��|T ��m1=Ͻ3���1=�'��c����I�Bq1=R�;(U8�吋<f"���T�&�xvc��?�<�@k��dz��;y�2���;�q
����<ՉS<���;d��%:����8<o+�<�<���2���%=$�:��<%��<�#�\�=_qW��=���/��j��(
��̼�|=�T<��c�t�T��jA<� )=T���e�<��=��¼�����}=�z��S!����tC<��<�.G��f�B-*=�޼�L��J^a�񆾻�����F<�2��}��;��==�6=�Ȁ=��J��7�<��T<��<z"�����5JK��< <��P�,O��"�L���b�R��@F=���X�	=,Ͷ<�B=mŖ=dk=�S$=� {= �<w�5�*=iS=���<��]�-E� �Ǻ02��wK�h"�<�f�L�!=t�G<�y�<��B=��%��W�2��<8��E֪< �ּ9P�<�5=�=�"m=� 7�?=h�NE���0�h�f<�=��Q�s�=:x<���b��cS��q0�z��<�S}=del�����}����I��WՂ�ő׼`a�;����(�>:`f��Ӑ��K���m=���l�;��m��<�iH=�5$�K܀��O=j0.<��y�{��V��<�B</by�Pw�<-���c��ED=!O;�f>�+K����G=AѪ�8Ձ����L#Ƽ�t�'*=t8M= ]a=ޛ2=�9x:�i��zq���`M=�k!=�.�m�Y<b�.�A=������:sb�<Ȇ�m~F��v�<�{���=���b:=�<�<_<�(%<'<�)�f���KEQ�~=�{�<|v%=�����6="���w�=�Ώ<Ҿ2�Ck1�:���S��Vûr[���ȯ�n��ȼ���;�b鼨��<���=�6=��r� �7=��˼�dG��m�<_�Ӽ\��<#�Q=åA��0�����u綻4�L=��J�ZQ�<��<�ˎ���(=	|�;ZM�&5�<x��<S9=�"<�%=g25=��p�u=�<B;==�<>[��c=���<�=J�g���;jL�<K��[��i�=���W� *=!jK<A��<��;�H!=���<�����/�$R%=��I=��@�~s]��,���8��J1�E7��H;���<�"��������I��;�^=��<+�:=�k�R�G=eױ�e�==��7�=�R�=;A�T�z@��=��+�9����K���~�lc��s�=ޘ�<�a�<x�b�y��<�ԝ<Ӄ�<����N�Ð�[�<hd.8������D�}p#=0=�q%=�?A=[id=(�<ϡ'��J=Rg�<�t/�6�q�b�;6�B=m/%<�D@=�U���?=���;t_�����v��������պf=�n+�k�L��8�T�O�dp��Xg�>����~�L0=(鼬�１=#=��<Mp=�)@=�TL�P�*��(Ѽ�n"=�u�r~������1>1�6�E� ��=�b=�7<�Qj��LG=׸������%=��M;�=���<�{��f <�4u���'=\_��T����#:@���H��h9<|�_��4���":��=%�o�'���'9=ٚp<�f��^ ���:=�<G�Q�`����</]=e���=�=@=*.=o[=����;=i{�5�<����
=��6���G= <����j&��i"=:�=K,/=��;r�һ�d�������<BR���8g���y<�`=1%���<�l�#V�<'�s=n�Y��m�E5=1s��%�=6���
=�0��ʇ;j? ;@��<�=a�1�V�y=|+������ݻ�0�3�P=8�4=�C	��炽�黍!6=hc��&�3���=h�������/=������<�KK�s�&�=_�;8Y�:ؿ<_"�=�zl�
_=��J=��9=�l����7=֑���w_=�<=^��<i~�<R�C���<�D��,hռQf�<Z�%��GB�~;��<��[=?�R�^�<w�_=�Ԩ:�R�;4wS=$�;Up��}c����*=��̼��f=����^�<~���G��i��<�w���OX=y�>="�j<F�+=,2<�v=8���/ �t�-<�C=qI��_�ґ��-=7�<v==�(=�d��#��<��!���
=R��v�$�]��<)=�<�<��ԼS�#���.�c)�<ЙE�����+��Z�<_��G��+`�g�������<r�<r�>�)��� ��<�����	�YJs���C��=����=���b�@�6i�<a?<��_�wm<i~9=�I7�I=N�S<��d=	h��F%=�*�����&�<=�V=u�F<GF��U�#��{h=u�.�Ѳ!=�a�Qo:���< �����g��<��X=�|�<:����H�<�����Ն��&)�.�]�/�3��;#<Z砼~Rf��8����A;wE<�m.=��
��/
��ּiV�<�HͻD��<��t<�Hd<���<�z ���E=ٺM�Ѳ;�~���u�7���L�F�8_�<�f==7E�ae�<����C�ݼ��g�~Ͱ�.I[��M��2 .����;��x6����A�M�~�=�k�<~2<0�<�h_�� �<�r����ļP:=��<3�����m=9�<��
��g
��z<�O=ɷ�^�;��=R6=�1v=LIZ�'{s�k=s?�<:+^��Qͻ�)�<�	S=��8<��0=k"5��7˼�!F=��!��6�=����=�9=�촼�U<��3�@i!<-��<��2�v�F���Ҽ�,�"?5��V�����;`�U�w�<�=NlX�&�H=�I:�Z=�-=�hx;��[��uz<`�B=?�T=��$��H=�ژ�j����ҷ;�Ɍ<�;�V�<l�Vi�<��:�<��<(L=�� �`�8�-�~��;�6�si�<{�a=�kU=��7����U����5<V)�<����>+�<�����-��!�<�l��:=d�<�9���� �<�MA��d4�g'��*�<iH�<Y'�<?9�Л =I�P��h!<�ߓ��.=��t�IZ2=5���'AT�'�%�b�	<�=���;�FK<��{=� >=-���%=Y�����<aN=7���}���8򴻯���FT��'�.#l=�R=���oκ�`��6������!�<==U!=OA��)�<�O=�	̺�o=��b�PQC= 
'=]'|=>B�<��D�p-�<��< @/=��Y=�a�<�<�꼔nZ=m���oO��Z=hS�UE=aļxm�0�S��#�E~���=T�p=�7;�����ݼt(=���u��;i���K�;k�=�:-=t`Z=�����x�<VDl=�;\��Wa��m@�J�<��B��7�<O� �p�mfs=�[o=�rG=�>�<г>��Z�<p[���A���p=-RT=�5(��J<��y�j��s���9�L�Ip�<85�f{8�m^=Q:�<�Ǝ<m�ļ�)6��X¼�G<ռ�#������;Ԓi�|B=7U�9Y"���W�;��R���3���D��CP=6v"�^9M=N�=��f���X=�<��N=@���<��<�3=	�"�
h�#
H��;�WC=�o=&� =�b���غ�����U�μ��?=��f<���[��:Λ)�g� �|m?���;=��=�,=Vw��L��%&��2<��)=�k[���(�Ҷ|<a)=oe=�oD=B�<��/�mЃ��~<�j=<j =-,Y�GH<"���P�|:E���W�݇˼N=��<����E�8�`Ѫ����&$=N�1��vm��I]�;�==��<|�R�]ʼD_����n|���<L<�<-~���}/�x6<q>��3J=Z�żr��<}<�oh;&qڻ�Q�<��=�3[=6���6=&G=B8?����;���<�<n=�{�<���<%6=��H�)jٻ55G�>6�<S�p��b^�Y��<NH��2>�<؍?=�tc��Y���6=��M�տI�2.�� k=��e=� L�ރ"= s&�'$��	e=xh=Lj�;S��I{���F=�M�8=��-�6=̾:=	=kj�5EL<p�=�n��}�Z�	����0�<�����c��d��<|��;!h<�Ɖ<�	�<�~�ӴG�$њ�ܫ�;NA=�9�u�)���=(- �)��;{$���<��?�<�9=t�Q��90��y=����R�B���%���o=�a��˼]��P$��0<3�=�2�=�i�RiJ=E�u�\=>���/Q��]H��kP��Q<l��<��+=��=dn�=;�ż�aa�%s=��5<�Y=��q;[�<\S�<ߢ��딈=۷2=�j�<Q"伧b�<���<M�X��w$���<��<9;q��'�<��?=��;�xN�$N%=��<2J7���=Ij<��:>^=�-��;p=��=�) =]��<�m.��
g=}�m<mC�Y"��{�^>-:���*y�!��n=c=K��	1͹�5���d�z�����z�<%�����<�99�b
���ȼK=$��W��X���<�����	�9:�Eڵ<�u`����m���<mey�����<I=�Z?��G�r�<�F�=�7���,=��Ώ���1�4G;�zJ��W�x�H���=���,��9׎��w��#� 0����=KA"�_� =B�5��_<��I��ч;��%<oI�<+�W����<�,Q�<��mנ�yl0��>:M�	���{���)<<����7�*�nb��\�<��%�w=���<�%=Ūf���H=��6=���
0h;��T;6F@�4�$�+*�<7�<��V����ca=U;x=y뇻�S=�^=w �-氼��[�b���4�%o¼����q���_W���O)P���[��(i�͈B=C=8����v�i_:��	=|\=g���2���Y<&�=�3�<���;T<jG=���Y�=/����<�M<�u���<��<�ҟ;�7=�6������?�<�����jJ<_�%��qf�H���\g�4���u=����j��Z�<�L�6���?=[�����Q=5bc�G��D����W��<�X�<��~<۞�;<R��L�{���E���8<�GO</�;�A�;��=�W<a9!��G�;v�=�|��0��D�7=�\��d�ڻ@K(��w��P<�om��:=�<�Ȱ<�~p=�6*<.K<D�S�/�<�*����{�;=K,�3�ڼ+��+�Q=v| =�(��h��D����{�ԎG�E~2�6�ټ�譻��2=��%����<(��<�Nq��+j=�?^�L��뎈�/F=�75���C=��<���<D{����<�un����<�2����;:rN=�\���=�Y��V=�@6�,4ڼ��ɻ�rۼ��r=�wD=Lad=��g;��O=MBl�O��;���<P.)<��F�e:�<b�(�%:������<YG�<î�����o�<=�:T���<��)=2N��n.�O�����<Mu�{�V=�T(=m�-=,��&��<c���=�ۤ��)"��CL=�ҹ9Թ�;�z:=�D0=i�R��|<����@2=��r<��V��K�� $<�{��:n8��J�;��<�����;�A9=��B��<�eb=Hw��<h��0k�<�� M;��=�at���6;m�ѻ���y�P;%=`2<�{Q�������<h��d4
��0��1O=���7����7�-y�<8�=�Y���;=@?.<����yI=8D��U ��> ��<��u���<���B��μ��<k=���L?=�����>'�U/=�=7����M߼D��"��=��4��3>�¼�<?EN=���<�t=��4=�t=dl<�:=���<�I;{?�=D"�E�ͼ(�=�b��Xu/<�S=�s3�E�;H޷��h��z��D��K�n<��B�Xcw:s)��e<WJA=g+=�2W���i���[=�Ҽ��T=��=P��<׌���G<|Y=W�>="^�<(D=1R<����*=�ǽ<�/�� �<D�7%�6��<��АA�n<���~���;=�=?=JR��Q�:�hx=Cz���u�<*�ۺ�a;=x�u<�q�q�S�������,=�����-;/�}�lp#��ez�/��<@���@O�Ur�;�BL=5�����@;�
l����<�:<�~^9�;,=�l�Z���!<�I������F=�;w���7|ٻL	=�;�)�|�1�9�D�=P�;p�A�!�6<e�:'=٣>�=�;�A=�j=�<�s����;�`<�Ӄ<0�B�ZcD���=�)��u#=/<܍Y=�WV=?[�;ჼ=7E<�~9:a��D����}J�<�q<�e�/�bE�;�V�<<�W<
��;d��<9%ƹ�;4V�3�Y�$C=Z-�;ZwS�U��<�BT��he=Pj�;�Ʌ�i����B�{�<�� =����ז�<b�"<�BD<�p�<B��:<�M�i���*;m?�j��=~�C��/��fl����ڼ�=��ϼ?�O�V�Y=�|E�&9=QU=�1�<�F���;�w,�;@h׼�Wμ1����<e���mr%�;�v;���<�=	�;=�u=6�\=$h=��<��8=d?=��W=�逽ء�<��=@36�e�X�;���&�=rA=E�<�چ���;�W�z#:���<5�=�G=��-�7�GU^���<=خO��28<d�<�..<g��r�Z��[@�u\_<��I�c\)=���<���<5UX=[��<g
��^)���\B�c=vrj=}�<��<���<�8=�Y5=�O�{��<w���E�SZ�=�؅<C�u<�&;ٟ<���<��=i�U<u&��'nU����P��V��<�4��S�=�Wݼ�U���=�/b�<��������7�����	=�4k�9��<pܕ<&<:<�n= �H�&�x<Ӽ���Z+���8=W�
��O¼ڼj��Be=_���"6=��ȼL���!=�D�<	'=.��O��I/ <�5v�U++�6�<�r�!�ּ��>=C���l�f�J���M8B���{�)����I��	B��Z���Լ������'�^�`=0�*�0�!=�N�a<�MP���;�~�t��)�<���U?=�6�<���:�&��W����)F=ź�<`���i��U�=[����N��n0<Ѡɼ�IC�ާ<{�&<��<�V+���B=9�<Z[ <(���yN���n��Z =N;�<ã�:QdI=��e���h<f� ;���	i�k/R<$�M!=*Q�<F�/��C
=����Z�;�@���S��=��ۼS7���6=ΩU���<�(��`T�� �.B[=�	q=u#:�|��<G��:2)P=��3��5�<�S4<q�-=s�9��M�l�=	-�H�H=:;��Z;M��)*�,�4<4cy=MN��=�sD��? �6g��
���	�SA��դ<�D�;p5 =�o�<C����J�|��<i��<��7�c�=� WJ=��6��j�=� �<_����3�G��;�]j=�a�HLM=��+�o�����<�x��\=�*��w�3=��t���_;r�;�c�$==��>=�!�<l&��)q���4�Ͱ<3N{��r�O�<'��<���;�R%=2���Tf=#J��o�)f���E=��3=�=�4˺��=��f�;"�:�B�;��I=��S=��<��;�<%3�<B�����sa;6=ֵ|<�L=�@;fG=x���.�T�rT=�d7=�.;�oH=��=^��<��v=����g늼^`==��;Pd>�¢:��2=Eg�<>�V=��B<����E�=8Aj=�e1=1>�<��E�W8�=�y�<���<��I=`=��7�k��:�����Y<�)=�F�z�+Zv:Y[~��P
����<#������U�<q��+��<6_�<]AF�m�N=����y���C�͟�����6\<�r��а�<�ř<��2棼�i<�1v���A�T"�:��缧����+�<�EI�uMt���Ҽ��<X�3=��T=��=�_=K�?�M��-bM=��Ȼ)'�/Y=�^=�x,=�!&�(�= %��A2q<����<��3������㻊+M�����h=Ft}��Q=��0�rּV닻!R	=#:=�S��,��i߄�CF�<�Rp�\j�<�FO�����6H=��m=G�`���)�`A,={��d�SB�;��k<���F�����<��^=\.�<�|Z��-��ڜ�<u^�;:�K<$����a=���<��9=\��;yj�:����\�;�P2=��=m��<�==����c�]���Q��g3=D<ٕ�:��={;��I��E�� m�<�oW=�`=�r5�.��h60=��"��*4y=�$�kh��_$*����%�I��������Z��:(�<��;&'�<�<=�d��F+=��A���e�%�24�<�(�a*�/J�<���۔=ӆ�<����L=�x=bat=�&����w5@�I/= 9�㙾��'D��N
��(*=������J�-�#�ؼ��+=�T=G��#<bt;��?�/蓽�'��=pG=H�>=���s�<�=ډ��6�J6
=/0���8���>�<H�}<��J�V�<L*��6��̇�ws;	��<̓
<v�9�j[��F�0�B��LKr<����R��T�s�I^1������}s=qO=�V�� j�ϥ��@��꘻�]^�Ѭ��Ԭ�������a��;f��y���2ἪA=�<���
�:<��R�8C���'��8�"=��:6�d<p8=�d̻��&=�6�<�}��NpU��M�<ӽ"=+.L�;�
�g�0�*�
�r�;�!�c ���<
]?=��	=5����W=l�N�rn��$F>� �W��Ƴ�4C7=�Nd�w�f;���]�F�Q�׺�!<}��sD<��V��:���6=��Ƽ�l���G��mO�Pn�a��9.��8�;2�<A�Ż-l�;%���S¼{�4<�������u׻	��;@�0\漤3:�AɺP�� C��<=��껅�Q�q�	=H}�ا =k,;u�:�
nT��֮;Ӧc<�h�;2끻�<zZ<���=�ͱ;��=���٦,�d���Bء<��;>�߼L@=G�,:5N=�?=V����[=�)z<9�i<�ڼ=!0=�!=�����I=�==�ސ<�܍�h�%��Z
=�|�<��9��J=g�S<�H�<���!m���"���,=θ������I�=�F<	�j;��P�N�=���Z(;)����{=�=؈C;)�ܻmW�{�K=u�0���0!C���@��qu���8��Fj����;8V<�Xn=�� =r�
���%���d=��#=f�I���;�*;`^=-��<+��&�<+9��p&�p�!=�<a'�����4���j���b�=�h=��<̞��O�2��U'=ɍ�<��;�����:=A������ ���Ak<2#d�����r|9=��<��p�<�H�����9�p:�@,Ӽ'nF�U��z�Ƽ�<DZx��J�<o������j���<�1�����<S�<ӻ�<�$<=O�x<<�T=p�G=��]=`~�<�TP��=�<�y�k�ֻ�л�;�"=O{�R��T/�;�8�;������E=��*�ם:=���<|3�<c��;��j�t���LI���W�1EJ=l�E��0���1�·{��{�<%�<�i���5=�l;�6<��&����< <X�=͸)��Ҽ�]4�f�!��m=?�*;��$�<�/�;h=�٤;�<v���g<���R�bfԼ�����޼L֒;�~/�n�g�D��<I�B��u�=�F�<��!;Ӥ;���Y����0=ܼ3�)���Լ�)T��Z���/=[�>�8���9=*�<%|(� ֹ�T)��@<�ﲼ6WL=ަ2<��=p6��)=�R=ʹ��{����i=�	~=�5L�KD�<I�%<&=���Wc���L=��]=w���y=��=��D�y��!c�<��w=�o��[��@���C�4KS���n]-��c)��-W<H���ļ0ԻHqX�2l~��<U�-�u���=�A=��=��w<C���>�5��*�D6�<-��������W�{�y=QPS�4��<�g%��w,=�&Q<�X��3&����5=���<b���*=��<��C���,谼��Η���Э� 6�!%=l%D=+�"��U��K�=Af2<-�s��
�<DX��>骼�輺Ry=���<#�� ̼�23�}�#�{��<�f��>�\�.�p:W���偼�,�̷Y��<=�ج<�ܖ<�4�:䝬����<�k�<��o�%1;=�_<��G��7�<ΐ�J��= **�L�;2�-�vx���<���;��t<��
��& <y/w=Ad1��^A�s
0=��C<�d�<g�7j5���߼�| ��i�x׿<��n����)�}��<�a�<GR=M�Ӽ���;A3�<<�=�#R��}=�j�<G��<#=�������c<=a���0gǼZ<=&�:=Z�<s0<�ֈ���=�g̼��<�}�<���;N><��<�У<VU���j�Yr�sZ =t=N�<��3� �8��'=���;ZR�:�Ҽ�E��Gt���=���<���B�j=��Q=���9���;�Lؼ�r;�<A=�{��"8;,�=��%=���9 ��8<&4��<�<�N�h�W=g\����4B=��G<~y��ka �>�"=D�8=!�M�V0<,G1���ܼ^Q<C`=}�����,J̼U������d����Ǽ�o.=y	�ᾴ<�o�tƼ�Q!<'�3;!r&=�.�<$ʉ=�)=SC����;m*<[�!���<���<jg��%?=e.⼹P�<衈���v�j�����<�/c=��9�|_=�a=��<Y2ؼh]�F���c��b�<��>=��j�����;8�p��&���}i����;���u�b��a=Ŭ<j[�;�燽P-=.����s=�$=��;���=tZ��K��<��J=V�a���B��9�<���:��NP=%�Q=��=��;�Ċ;�"�;��<���� �<t '=U���0.�<�YT=����Ӝ<K3��;�;nm ����<��5�,�]�_��<���<���;T�A���ؼoS4<��<�`���==:�R�]���}����=y��<]�<��H���<��&=~����<|=$�-�$�-�0e:��E	=)�=�t~�������2<���:�I���1d=�I
�7� =W�ڻ�F��@���������K��<�k4=���W�K:�\��ļ� =��`��}[=��i=���=v�<��&rG=("T��&�<�|ɼ3�w<"�J�$nx=�R<<5ܚ<��A<�Z�<y����q�X�$=��8<���<:	���U�X Ѽ&���nּ�v།i��y��4��]z��@"�;!0{=��l�AO�;�7T��=�:=l����B=DgT=V���q���q�<�P��7=��;lC>=�8@=�'�<�]�<�,�=$'��7?�Dd�[Ỽl��<����ɼ61���b=�A=�.��~�Һ����#��:�BR�`ȁ�v�<Z<��Zo=��X��/=m���؜���@����(� =j�\���ʺ�}\��&��OND= �'=�dt=+��;emE=���< ���u��VI=*R���ä<[��A��9=��;���z�<���<~<�;�<h��:B��Y�< '=�����u���{�<� ;<�}�;�Q�����߅�=� ��Nӻ�����~ ={1%���9< ��<o�-=�nZ='?9m�=H=�ǝ��i'<�=�c�:S�N<k,(=t��#�<؈��h�<���;Hm��K�|1d=mͳ<�J㼍�&�w�=ث／}���<�A=��r= ���9=�:��S;���<��ݼ�j&�?�a=b0);�C
=ꍰ<5��=�_�ྷ<�Q��o$��sq�Z"-=y�<���.���G�Q=V4�:m开"�� �<V0b<���0��<f3<��.=��Y�2��2=*{W�U��="$�OoT�^c<g�)=��0=�Ũ����<4�ټl�V��^�=�q���k�<j��@����}�����^>^=N��r��:��Y�����<��=��<��9�Ԥ�y�i:�2&=��; �=M7=¯�<'8=j�=;υv����]$����[=�=��ƼJﯼ��C8vB��5�!��bM�fm��o/@�%9C�ü ��=��;=�ގ=�m$=Ũ#��5=�kM�n9;�?V=8�=�W�=��<�)���L=��b�G>U�"�.+	�g*=\���G�X�K�[�p�6$����V��h8��u[���	�P
V��Ѹ��Y1=P�_=;d;<�A=C<i_�<Hy�<�r
=~��������=�Zu=�c�9�筼��x�Z�=%�O=˩�<�I���S=:	��zu�	���uW�<Gv�:٧P<w�<��=��W�#rx<��=I��<����Ƶ��~g=������m��	⊻t<��-�o ���=��0��]T��o�o%�����]ü5��ޥ�#��<�"�� ���<E8p<z���X^<�ل�5�y=�ݼ+�a�W��=����g[�ޤ=ڨL<�O�<����8Պ��+�Bٷ<A�<o]=|H <�W6=��<��=U!�hJ�r�Z=� %=B�j�t˼`F%<���;�>A��^o;��P��I-�
��L�n��;-ch<�}O=z�<��<�*=���<���<K�z��Z���l=C���7�<���;��=��7=�����
�=�}��.��8#�]=�$��G�F�|�X�H�O���^<�==ΰ8=�c���I=h�!=�b=����+�:�ּmI�<�7�<1�#���Qv^=b�&=0����=p$Y�+KB<��L<A7�<]T<��!��c_=��������<�q���.=��*=8t�;��;@O^�)������<�Q=�/�<]��;]}K�3�=��<&���%^=�y��a���T�ԉ�3�+= 9=f�����<MP�-k�;�ڲ�bh'=H�=��'�m�#=��<m��<��=�ƺ;1(��CH��#�<֞�?�*���MQ=�<�=�e*=c`��&�<���:tZ�#�=��a<G���f<=a����eD�^�1�~����o6;��K�$G!=̌�|N�<½߻����:��O�M!�;s�X=�2p�O)�<����b=x�r=���<Im�;(m<m���'�e<��q�k�T�x��֙�<*��<�.X�����}<�Pk���<�/]<��L=�S��1\м3�!������<8�2�{�q��Z5=�焽ς#��UV��
=�c»U��B;�_����¼�Dg�2��<�ҧ�r�p<w:/<�Y���_(=�=�<b=5��3o=���+�=��	���|�����"���e=*[;37�;�e/��.�<��b=�?W�*뼨�x�b�<Bi�N�9�4=����.=$$x=�=ޓ=Qځ���
=���_��P"<�=���c�:;�%�9b��`���]��R=�e`=��$<�O$<wEJ�_=l<��=��<~@G��%=�>n��S<}Kֻ��̺U=	��<f=�M�	F=g|�1*4��@=�G�<[�h�G���On�<X�^=��<���EOK��.?=��<����G=�ܼ��=�)?�ʕ�yFټ��Y=���<�H�:��[<��m���漵�%�I{�u;�L����A�<���	9�;Y� �k�=��=��X�B�<�0D=q�2����<��＝���<X'��"���@<�H=�y�\1��>�=��9��pP=�l+�QT��d`=x ����+eF��7m=�*�<Ob�<j �߉E=����7���<�qx��8&����<S~�5;��G=w-мY�^=�4=�r��m��<��\���k��<�KL�a�$<�ú�5�<3���;NFf�<��<saV��&�:ñf=DÎ��q�<�Z*=�
�+��mf-<(`=�j�:�W�<W[�<�!���!=��b=�3��tu<+���5�=����G�<�������f��;n���Rl����0�.�7=!�P=U���X=�8(<��<Ldɼl䁻k�=b�<TH�w�<_���6ļ��g�y��<t�⼗�<���<� =L�	=�sh���=Gp=���<oc#<ˉ\==�R�<e,'=yp/=B/<1�<���<#=A��O=���<�&<��C=҃��U�&�(�<��3���=i�~<f�u��w�<v�n= w�]ź���<Z��;��:$)=��%�aO<;�_����\8[������)�a6�<����Q�����	�g�+�ؼaZS=�Y>�)m�<�l=E݃�ҳ���/y��UN<)ݼ�a=�:t�?�G;��͸F=h�;���<b��<�t=Hz<Ri�<I^�5i<;�=�J��?�`��.�<�L
�s��<Ф��C�<x���/�<�=!��<�v���#=l�c�r+��?&���l=re<U�8=M?»��i��3�;��=�F=�Y�<�n��
=�"Z=�	=n�+�CL�<&m�a���ys�4�<�V��?�4|��[�&!S��!^=�?���\�.*/��@5=g�:/O���D=�h	�%��=��<��%��0�<eGd���뼿-򻭻;�����=kP�JÜ=y��,����h�<��U�q�i�5H=uF���Xj�<�����W뼥;*;��<���<a_�<�=p�s=FC=�ND��x�.:Y�R�;�D=���<�we<��D='_�<��¼M�=�j<�;#�=�`'� ����?�N�]=��;�]=��s<�<AIh;~�.��,�;c�����<�}<�y:=$Z�<��b=I��U�<2�����-=͛1<<�O=¢�<گ�<�j0���B=�@>=��"�>�=q���L6=� =���&�������<
Sf��R'=�a��_��L=(�<�g5=Dǳ<՗���s=��=����^8��ˈ�'�=�X��%P�m� =^���+ڼ�Ⱥ?\;�����M�w��<Fz�0Qj;��;:0<��a�a�=�'a<--=�8
=�_H�U-:���&=8�=2~S=@ϒ���Q��w;=��Y�«��";��<��:=�e�4�Ɏ!<Ϋ6��:�<�_#=yH�4p9���Ű^���˼��{=Q7�_pY�D �)�E�
��ܤļ|�����<���<��<��=�	^<��<FrP=i�p=sRB��н����<�Z=��
=��=�=1+�p�G=���3x<=�N�����G,=��<���W=P3G��&����,���;(�-��	=�a�������<�$��;��#|R�I�<r@�<6)��:	���;��-��O�<��<�Sؼ*��<O<@<��;���<��l�쬳�H>J=���<" ���<��7=2c=��1=�N�<.K(�6���+��E~ؼ�־�Tߝ�5�g��s=I�м�<[E��=L�(����\=��;���b�<��W<x9Z���������~�b�<߱�i���k0=2p��j��<�E����c��Q�4���=hB[�W8<=�n����I=G�=KY4�9\G=:u��>�('��/���=�:��<��=K�!�*z\=C����\���<�<D��S�{��{/=J��<�Ny�.�+�B�Ҽڲ��eB���5��!=½��<�E=�(r=��=AE=�Kx�<f=�pؼ[i-��Sc�Y�-�:T��k^�[|p�a��<���wC=/N=��g<��Z=k��v6<�=m�����X�<�u��V�J<�E���8;ç�<��F�p>f���=^dW=�>�o�4�q+=�?�<t��;��C�{"�>/_=�[�<C���7�="|�;�;q=��;\�T�~����O=0�L�?�d�z0<�0��</朻��ºa8��A�X?=�`�6M�<
�=n+O��7��P\��m=�,<=�Z0=�퐽�΂={�O=��J=9���w����_�A������<��3�a���ƥ%�G�P=nx�R�]=%Y�=U�<�&��H�<g�W���м��<��<_$�>�n=������==��L<�=��(�J�$��<A����:���<��<����=	�f ��{<G��G�h��W�:p��I�<@�[�afq���c�L�ۼp�=�7�(��0V �cb��Qx�U��L�Ҟ�<�E=Ɉ&��)=/�q�5(��A�9=6��<��]=�g�pAc<A:\=��;�I��P��Q,��3=��<��=�� =�`8=�Dż/�<�u<w"�uU[=ɵc���=v|=AN�����}_�;a�=>�A=����R$=k!�<��S=�R=�A��:J�ȠV��GS<+>�vk��-� 4��ID<�/��D:�<�K�<^6+=�-;�x��9R	<�-<fG��s�;�ȼ�%���<рQ=9^={�����Z<I[=�7=���tȫ��p��IJD��8�;�9ۻJ��;z:�	��F�b�3=
#��R`<��k����9(���żz�=�t�<"��gh<�1q=�3=]�Z���G�,�M=�&Z����<j3�:���<�f��<6�o=2Y,�g�@��^<Ip�<r�:��S=��A<N��ʭ�<�@v��T0=��=�T��p<�a�=�u�^ �<�D<���ɺ�yX���"<e��:�/��_�9��0A�4�������M=Lr4���[�_&-�u�b�	μx�=i�<��򆆽d�+���F�����	�w����G<F>��$_=�F;��}=�-O��+漬�={�K=�ӷ�:U=ॺ<<@u<eU����9$Հ;�Q�?Y=~��\i���l�;`�=A��<L�N�@w�<���<z! ��/=i�<y�T=ށ=�ȉ����������<�����F(��k<�1� ��W*�z�;���!'�;b�S=G�1=��<�	�<z�<C�<|�l���<���[�]~����<'�����f;�&=��?F���<*m+�%�(�>��<� S<������a=F!�YU�����<ZH9�BP�x�,=������<�+M���<�kӼN�X=fH=q�==���J���b�a��!�X�����VƼC\=b�?=\~�=�[$��E�NIB<F��Ls����l�1ꤹ~�#=��<*<=*|?<e#n���F=Z�<��:=uV&�}�r�O�v=�d5�eK=��>��h���<��F�������<��5;��;h���9�<��;�*=�:q�aH�A�q�j<e���BJ����<Qf�<Z0����|��8������|_=���[��@=�^5��$-=�Hn��#�<)O=�s�kKV���X�� !�
v��#�<�����$�&�=�c;�B��g[��n����C�<�M�<��b���;;�Wg=~J=&��!���<� 8=0��<�?=�<�3#=�"��=�:)=�_S=4<�=�V����D�[!1�8��;mPӼo�ݻ;� ���T=�ބ<�E��^=�ڲ��L!=
T(=L0(=�	�"���W<6<�����=PW9�t�Ļ7�=�iS;?������1�*æ�q����<-������<�5<Ϥ���pżQ,[�`\�Ƴ�<��=s�=�G<el�<H)���W=���v�����*�
�}���<y\^=ִ6=g?��*��J=��	7�1C}��߰<�5�<E|=�ڼu�P���#�nbA��y)=�?z=�j�:���:�\?<�{�9𼛄%��>:�����~pn���Q�4[%=m��<Z�)=&�< +=C�ɺ���<�u߼w��;=-���V��ئ��.Ku;J=��f�υZ<��<R6��r�����L̻1�=��6��|���༙�$=#��<�E=1m�匏<�n4=z��DP�<s�<�M=�A��v�G�������M�"��<���<{,k<�S~=>R=�~�=/2�0������� ;���<ѐ��6��=E='�<��]<���<�}e=jQ���w��b��iQ=��T=�6�+Az���V�����6=����S끼^���1���\a=6>���;Xoa=_2�<��x��������:�I�:�;B=y!J;�E/��H��/�ü�R <7׼n;=�G���d�cf뼅mA<�=|BC=�g�<���rW����7[�;�)ļt��yD�:Y��l�û#'��=���(F�:.<=�9�
s�!��Ɖ��B���DF����=�����;YM'=@H���e=�*�<��P==E=n a�.��cU=E<�24=J'G��Jk=/��<�_���;�-�]�4���U��ٚ�<�P���v�Gǥ��{=5�];%�e=�{=�%��~��<�K�;7��;$��J�g�>�M��!������<Xn=�%^=i�k��<V�����<Ԛ�<�7	�G'�<�����X=�;=�#��,*�̟:/d���o�D��vE<bQ��G�G��p���a=�T�}����;L+���(<�to=����j��^�n��3=e���ψ=д"<𠼸�9��o=lL ��J�v���Df��\��#�ʺ��;4�^=���<Q�</��Z0�<�����;��%��-<q+ ��\=��'мH��k"=��<��ż<��-�*=L?J�*'#=�I�W��a~H�Uk@�����n1�;Y�����:����Bգ<c:=/�U�@�'=�	�����<��:��=J�=�)=G�;���9Y�R<�]���n��M�<�=[81<�-�<N?��g���>=וd<N+l���;�D<���<���0u4=:p$��7@=i�n�lʦ:�yN=K伢�"=��=\	!��d�f��<e7N=��8=�����<�g�R=���<�,=E� ����g�;��=��<�lH�@�-d<Ҝ9�a�<�)O==�L��=��J=;�b<�
̼�<���<u�z=���<�%�w}=j��ra<'���mu=�P�<�V\�>�R�0G�/Z�<ֽD=�9<�HM�j�h=� ��p=ÿ}=��A��<C<e`��'ۺ�<�
D="5�A�=��</f(<��2�{�|���-=e*=�����=��)��������<����c�;.�[��m=�j��˯e���� �X�[�W=�Z/�+ܹ�e�=�|�SA&��D���<��
=$9o=C��8�{�G��\�{�W��;�l�<P�<Օ���67=õ=}F=�6j��M@��eP��c�*oE<}rX=rv�<����<��</Y缽d1<�/4=��7��^�|�&��S<LԒ<؎#��<���<�Y��cI=VԼ�x.�q��q��:
���@F������$���<;<N�-\&=�=�{���=v =�ܼ�����:��[;.����� ��h����R�Z=�,\�G�U��-.<��8=�!]=��>�F�4�ě<T��<N%;=��1��	¼:�<��9=�μ�`;=6P�/J=	���9Һ�̜��=�p�<q�@�<uw<�C=�$k=�h<�ي���<D�<�@~�M���q�μ�ܼj�>=��: ���h(a=
��=we-=\�x���=.]=;�G�<��3��x&����M����Y3�xp.=��&���>=M�ü�(��#���;)-9=򡙼V�����=�)=2�T��W�<�p��������<#�a��<e���n�漻��� +<|�
��U��m����<��=�!�<=Y�P��t=�Z��2R2=�{�<�;���;�P������P=�iʻ�'�׼/�7�r��<]�.=7A�ײA��qD=Tc=��=n�3=6��<�$ <�I,��~��߼Y�һ?8F=�!��T=D+�.e'���I�U�ǥM=s��<LFW��䄺��\�V=ڊ�;xqz;+��<�2<�Qzx=��l=��r^*=U��;(��<I��<�P=�����O��$)�D;�9<U��c=��0�2��=D�g����:_p𼺘=�r[�T�v;���<����)�;�9=eS)=0`D=̆=I�J��"μgJ_�]�=F�9<��s���I�>d�<K3�;+���/<�3�$v0=m��`��;�'�;YPY=�^�<zx�<�>��΋l��o`=	��2�;�0�>��<�����E
��2����;�{<��	<5�>�X =�ἅ�8=K*<HԼ��!=	z���)��yn���Ѹ���
=�
;��=L��9�e�����;��C=�W`��\�<z����L=��d�pH�<|ܬ�����������:_�=4�W����<~�=F�=����<�����w�=�Q�14�<G�2��'U����<��P��o����,=\�=Ó&=��=6�90=�Q=
;=����]�<�-H=w<e��<	�<Gm=�<h�d=7Q���<����Q#;&��ͣ<ZϹ�?ǲ<�����S�Q��@Y�F/�<¼�M�B���=;k�QTh��8@��O���]=Y�_=��F���w=ky/�i�eOA����<�G:�0�g�'�;�ۜ��J=df=�0=w׃=&ѼNn˼G�����<n�����;��O��!��F|Q<��:=��V�W@�$�/<G�8�a�<�����~����;���tЉ<p�]���O���[]J�Ϥ-=�{=� �<�h캾}��E�=�d����-��c�<С��8$��_J�<����<� ���F=�J%=�����N���8=��i��$v�u��:�aۻ}�༚7@�wdk=��
ͭ�]�9�>=�#�ۢR=���M�;�����Y/���=�LZ=L<���IR/=���<$���o��<�>#<�T�<�f�<Y����$�_�w=��V=/�w=���<������|< �w�Cv<�6伦C�<ߤ=�0��TK=�3=b?5��uS���;:W4���_D�JL�<�=<O�_<��.<kU!�Ǐ]<SpE�̈��-ĝ��)��p��[W;7ID�J��v�E��
�{�;;,a=��p�<�<e�A�<����B�=k��<��<��W=��<	hi=?�-=U�-�	��=k����!�;������;�i4=y��S��'�B��;S>�<ݳ��
p�2:G=�GO<˖3=T�=��M<A����T�1��	V��A&��^��d"Ȼ,8=lL��m�<<��[3=��<VVX� �m�+��<�E= '`��ؼ|8 =��/�W����=qR�:@��\����<���<���<��<�#V=1d�8���<bW,=<��AB� �T=��<�"O<�Ā=��� 7����<K-&���#=����[��<^)���;� ���M%=��g=E�U���<=��I��E4< � ��W�<ބU��� ���n=�~�$��jY<�5�d���p����{>�o�y�H@��������<�N�')t=��<P�<�[!@��d<�=m���=H�#=t�z=��=ڶ漁N,<��<���`2�{
Ƽ��=�^��<ő��'�<��=ȶ<�U����������+9i�E`�D��<�ii=զ.;׸O=K���F=�c޻<b!�<���;��M�d��<Lp*�5�T�����Nx<��A�X"e��Pټ7=Q�<�G�� �&�
oͼx�#=�u2�B�	���3<��=iʀ�-H���L=WY&�<Un<x�?�~�)�I���'.�[)�;�������<��5=��<�;62,�����a�&��
<7B{=�5G=��<>F�<W��<�=j�=�s�W���ۼ�Y�<��o�jZ�<��=��I<����ڎ<���2�ڛ<��%=��=2K8:9�8����<$m)��Z=��U�7F=��<�;ϻ�]��*�<��<=�0�<�զ���C=�z���Y�>�{;ۗ=��B�ݽ�< Y޼��<#v,<�F�=�I�=pg��9
��q��9f�
i<(8V=H�<�K7��G׻�݆<;���f��;�p�;F�B=/�1�=�E�<<H��S���|H[��Ή<y%=����o�� �:�(=�V�<�ȗ�V�<��^=��==��i=������6;X?Y=��]=����ŝ<7C ����������=q��<_Zp��[�B��!�e9�̄�� ;�O̼�\=YE
=%
�<l�"�UO=ͨR���(=���^u�<�
漢F���:1�^����<��*�B��dN=/��<x=��y;�+<a��%^�@�@�v�ؼM����μ��L���<�1�R����4<U�Q=n�6=���=ƃ�����b� =�bj=����9=���Z)�<@� =?�><��<��;��x���=�K��<���ȡ<f�}<�A�<
6�<��v���s<����%���$<�d��:==Ɛ:=A[�<���?=�����z�=H�#���|<	@r<���<�(�C-*=�ǆ��?�<��<��b�<��</��<���)<YШ��R>��};�������<�G3�6$1��J�����<���<�6꼛M�;|�~��
����(MA����{l=�Y�<��<�T�<jA�<�jv�Z-���"=��FL��=r;��]=��K��m�a`�Lμ ��<#�
=�;���N=ý�<�5�6�=�1�<f��;��K��O=V�N=~�H<�7���A�<=[^��h<�V��23=�T¼�8"���==��'=��%=c=���;�(=̟I=��<��Y=�t+�1�6=f�;=]b�}��;�=P�*��љ���������:��<*ZP�<]<=G<�j3<���<+�һx�b���<3�r�Rފ<����(e<څ����8�<!f���绺V_��0�B�v=�1�:Ġs<@5<w�;w�#<T<.=��w=b�=*�<1�=��<na�<	tS=�6�	���E/�iiz;[�p=�fL=�n�Y)�z�J���p� �:�)={���N �+�=2��Y�T=#=}I�d�=Q��:���e�=�;���;���<Pϼ�B�<x̼IM<����C=DV�M��<8�<��9x+��8�<��=��ͼ�(:�5;�\�ۼB}Y���J����<I =� ������U�=]����B�K�<ۢ�<cI�6gm=��f<��=�&1=P�O=g��<��g����aq<7|9��WN��o���gʼ�u=��.�i\=�ߚ��Q=���qo=��;�1=��6<���sy8��a��9�!=�,=�z<P-8=�mH<��0=�|:=5�:=뷐<b�}�M
5=�,�t�мܮ�����sȻ*	$��ܕ:i=_����Y=ɍA�;$�H8Q=\+=A��X�����6S�;OQ�;f�P�\��~�u� �Eu+��P��Ya<P�<�?=\-���<�ļ5��;1�����;R�<�?�n�h�va���Q.�W�<л�;U�l=T�Y�D1�<I`�<�&,<�p���N����'��,�)=�Q����<U1=��C��AF=r�7=D6�<y����!=��;���<�]�.��<M�@<��:���@O ��#����J��;��<�i;�&�:jQ��a��à9<ycQ=�����<�}D�כY�&=�M�<NA=!�<�7��K������g=c����˼U��;����yL�,�b=sܻ�=/*;x�m����<Y�3=������D߼}�;]�;�D�<��Z�m�G�J���p�sV�@�<{u =%V=��: �<��_;H�<~᜼�E��	M�;��<�/�<I
�H�<��N=�6=�䝼p���8�"=7�&��|V���<�*�eM<fH}���N<G$L�r�<�&H��i�;���J˅�3$�^�o�4b�7Nh<�z�<�-���c�d����=<	�:���<�ĩ<m�=�'=t$ռzU���3=i(�:m��C�w=t���וS��Z�=�Z+��6��Z�,��(��<c�&=��<p�����<������7=e|P�u2��WŻ10�=I�g�~�D= �ػ��c;t�*=�	<RO�U8Ǽ�k=�Z�<�$���׼4hk�Q��z�
�!�B{��G���0k���<b9=t⹼��*=C:2�� �;Q�/<S"�;;n=������*=)!�|��<3��t6��=t{��詼�u�[,<���<:s������+=KC�<Z��<�*)<��.��g���.���<$���ӑ�{�x���7<�s=Ik =�*<�T���;���<�~^�-?�<dh���M<4��<-T9=?��<����y5�O�]=ZC̻�\K=�8A�
���H��<6��{�.=�+��}G���=�(.<d
D�L���if�k�b�����z~=3�ջg�<�	�<F1'��I�-�	����/�<��)=n�F,=׹D�'ݼ�,k�&���#J�� [�Q�<���<Xs/=#��<�+ü�j7�"Ы<���� �@����D���<�w7��x.=�}�=��h��߮��*м�J$��l��.���r��� ���-�����)H�<3K�;��}=igN��f��@�	�e+�;[��<Nx8=ܹ��`&�M�E��'��Q�;�����<*^A=V�`�!*�=��>���v=R!�C�<	d�<6���P<�0k=�����Y=�8><ȼgϢ��k
;��<q	C=qI�<d�ػ�9=W;
=%o`;:�8=K��<��=V֏��Ǽ��<],;X�2�T=x�<��<ژ����:���<��:���j=a1�<?jF�I�<���A�/<U-h���������P����C=�o�B�<.VE<�p=M��<�VH�[��k ���<yՂ=NV���%����|;)��ﺺ�7=\<�2'=ī^�����=xV:=/�����&��+�;�G=< R�w�=��g�<����]����Mj^�����d���ʯE=_#=��� >Q���T=
\:��j8�ρe<���a�=����x���-f=�x�;��'^=8���Ue=G)N�� '�hY<��<%�S컼�Ձ=+I(�_�R<�/;<rmb=ɵ�<$��k`=�k��<2� +=�O�a3����� ��;$=�O-�Az�;V3�<вY��f=�����`������{)����<qk=��<<�{�9L0=T2l����<����Xe�^������X���-=�o�<�_�m�=��;���M�<(�$={�@=��r��Q0=7�E=�i�X��r�h���=�H<ĸ"���2�X��4�Z��`R=0J;_T=��=�V=WP)�u��;�H=%�C��'����:y 	��o�����\�U���������a�AL��.����r]~���=FS=#f༳���<oa���#���M=|G=X�<m�<��9M�q9N8�<���,7Z<t{=<dG;H��<P�<��q�_{>��2%�eWr=ŃX<�J�:Жz=�,L=�!8=����?K=͵%=��>�Yο��� =�<=5V=�C=��	'��F=�^=��! ���=|0x�Zv��Ƥ,�;��;"�=�Q[���?=�=�<	TK=C�L��0;��<�I��,���]�ی���X�W��<��;�� =md�<�Sp��"�vy7����;n��?=�T$�{5�~*ݼ=�|�[�j=5���t�<�ƫ<��=�|溣��<�.=8��<[�e�<{�<��\=T;<%�X=k�>=dd�ļ�f��Ć�E@�7*����K=�����c;�%/<�'=Ə =����Ȳ�k��<D)���=�=r��)�������=FW�=T�ͼ2$�;�7�<y"9;-d��=�g=j�V=��9=m���m�0=��Q��W�:�:=y� �S�c�f<�
%�5�:���u�W'�L*W;��=�@=yyf�Gn@��߼U���+�'_������q<�U=����s�<-�C='�.��� <W<(=I�2=N'�y�����<�{����p�V�˺+;q/W<l��<7^��ѡ=�3����-�./��8l=��7=�?���ڼ
gF��'l��M*���p���=�=R�<��=��a=��8l�X��<��g��8i<�6�;�������Ǽ��<=N�$<���b��<[�F��<�g$=`�=�����=��=mE=���<uI=~H��ë=H7=�` ��c�;/�=jZ�	L���1�N�2�-���?�{0�<��O�m]�i��M���r޻]w�<�M�<A�����=_Vi=�"+=����^Ἂ�c�Oك�`5P�u�߼�J���/=�Է<IH��m㼾E;��������<�B<j��KuD=�0Z��ৼ�Wz�R��<���= ���I@=�-���E	=	�Q����7y[��۾���=r$U:�Z=.�<(I\�����Y{J��5���9=Q��%]d��.}�)�ȼE5*�C�M=N��<d���)Ȼ�b=�w�<3����6K�ÂK�xcS�����9KQ����X5=q��u����G�v��:3�2�[|<�-��!7=TDR���E���%<*[�^M��!��<��
=69����<zJR�]k-=�Z�<ZP#=5�K=�R|;��=�YI<�g<�^T���]4;�G���'c<1R=ttB�7�K�I�=]Pc=|��<>;gK)��A�5�2�'�6=9�	�=g/d=�r�L���f����<$X�'G�<PEm;e�@=ݡT=�М<�=¼hr=�J;=�t��;���_<�-=~��<h�"�|�k<wS����<��m�-�= (=�G=τ~�6���}nV<�9�<m��1u���5�PP/�k�<���ߍ��L��;��<��<�%N:o!���=6�<k�:bP��,�<`��;�r;�5>=���KE�qO��Q2=&�4����*��<�4Ӽ�2�<��S�R��<f��9���<ijZ���=<d������6�<�ϱ�p��r�=m�/��i�<��)=��<�j��8J=-� ��8���5�=�5�<K���g�w=GfH=r����1<��T���2�D�l�t��<]�9��g`=�7?��5㼱��<�Ԩ����;1q=�P�:F~=һ#�6�J����|)����9�r���4��M="*�<�W:�T%�8I˼å#�Vw�<���:`a= ⅼz��T�
�p�3=]��;O�k��;Z.=��A�DG<$�=sL=v��"%J=�=�u���.<1=ӻ�<R���������<Z�0�\�3=��g=lѓ;�nټ@��϶�;�FĻ6�4=r��<�<
꼌����Zf=�Fi��:�<�E�;�5�Q?j=ЪԼk�X=�~=kP�<m�5�5��=��N<[�U:-=n�%�bFS�K���^$=�c�o{������<��w<e9��[�F�Z>n�,ؓ��h���?��=���;�Q��i"�6/v�A�
=�@�<��D�k���dB<8>��T�N5 ��=�W9<�N���+�q�+���ػW����a-�<��C��'�<�=l\==Rz�{Ω<�|�9�e;z�<=+ƼX������=\*��e:�n���4���Y4;oͼ�=��{=Y$���<��C<�	8=�(�<��A�(=��%��<��Ƽb>=��<�t����cG��� =&\�/p=� 6=S5�<���;��T�ՓǼ�~�����Q/�;[,=�9��e=Xe�m�P=�\�<+�+�y3�o\{�׊=�=xμ�<�2z�����ی���Z=�����}i��ּpʣ�Z��f�=:�<�\��b�˼��1<�H��hH<L�R<��q���:�f~��.��<��<$�W���$=z�6��z^=�E��j�K��_;O�<���V�=�儽>�9;��~<� <.}C��]�<�S,�*̇�8�8=�=�<e1����$=�E�:�7��s�<ݦ#�z12=�B�< �<	�ݼ�m��2� =�$r�7
p�	b(��\��!B<2�:b�<���=~������:��<������<L׮��7�;�:E�u��<6��<��l89�%<��(��Y��RA�<��+�A]��loD=�K�<�u=�wM�3��<ۆB=y0ּ�gH=�_=ԛ��@���лoP��{S<<5<�q=�#=C��<�,=po='�<;m�:w.<�C�W�=�U��=C-"=��j�_�G��$w=+��#��#>�<��N��*��a� �^%8=v�]���1�ܙ�<e����ջ�?�<&rJ��U:��:hv���;n<Y�.=B�"�L�ͼZe��5='�-=���<�^���k=���;=p�k5=��� i����<u��<и�<Re�<m.9=o�6<b�<!���(퉽�S-=�m`<�LH�
���A�;��]�=�v;�U<��-=��u��]�I���t�"=x&��<�^<Ӡ��[�x=v��׺G�n�C���b��B<\u�=�=�7�;H�=<}�ͼ8&C�U�<OjD��R�HͻU��;p�<��#=߬�<�\= ]v=��$��"=�"�<B鼈=�iɻ����>=An<���wp=�����Z���=;F��b��ڑ�`�E���=�EQ��=�+�<!
7��o�͕U=��h��d��f��`=uW<�� ����;�d==4b<��T=0P=V�!=[}<_t�<1!�����	=�!Լ�i=�I����w=���<O�3��W:�r�<ũ���<-��
6<#�;u]��{l=3�*����<�;�m�<��<U+��C�3��?�<��a��|�|落�_�<<�j�k�h��20=:��<r��p-=�<s��$"B��F=�10=�z|�A��G���;o���� <�ƹ��9�'>�;�7�<��<*��<6)�<��0=�.��.�<��<��F�u1�;���<��;�(�����$��k�h�.��R����X��o=��<��Y=� =�-|:�f;��g�<(�=6�;�J�!�<==�UF=�2��m<�<��#ü��<όb�()b�z����=�s��@0�E.I�-����T�<A��;�+<��]�i�=Qִ�9��<�I/�I�=E�=�0̑<�*�{�<�b:���a�<�a�<����t
��/���;4=I��;�%@���)�O�W	6���<���)�<:+�5�i�r� =�Y�$����<H�<A�y��q<�:c����Cq=�>�֖�N�<G�U;e=t�b��_ü�d�;���8>=�uH<�d޼���$G<��<e惽�2c<u�5� �ӻ2q7<Wߧ�p�<�x=��^=0�R��� ���E���˺t�<���&���:��ɻk�>���c<��W=�W�<MG�6� ;�n�</�;Q�=&%=��w<���o�b<d�<쏔<��<�F<����:�<3�f=ѕ;�3N�<�=�>!�r7?=68-=��{=�u���O���(��J;�L==�Y������:=!{!����$$�<�9�,Q<��D=8��;!A�7�D���'=>P��W4=�>��n������-=��r<9�C<�nA=����@9�T3=�3���A��l���=Β��$s�soL=�?�;R�hb=�5�����<��<�93��t<����\0-��� =�A<��/��4ݻ��<Z�^�jDX<�T=��<�G˼�XF<�jG=f��=g=�]�������]���=�F/<��;J|ܼ�d*�d�]<��=݆?=�*���{�:=t`���:��27�4ot<�Ҹ9=�=�Ǝ<�ͥ��d��u�~<��*=$�P�*�S=Z���[=}H;�ׁ=挻%�-�k"�<�+��A��<A���
=j*E=��	,�2ȹ��\����<:R}��qL<�]X��tA<�c���<�Z0�<�:=�
;��F=.�4X<��ȼ'<b�����$��<����o	��)��V(�3L<<.���E,�~�=m�<�Dj;d�=�6�$�	�O3���1:=�Y)�ड���:=��37��Od=x�,=�NI�e���N=O�"=2�Q�e6Ȼ⹇<C26���pִ<��=Dʀ�9kͼ�7`�N=��;~�����=�<��;�[V�;�k�;�����h<��t<���<�~���=1��<�ټ5�S���QDM=ɩ�Q�}<c�c<�|�<c� ���<�#=��k��/0=}\=��I=;x=Id3��F�;�S�E?E<*�<�'�=!?@��@����{���Լ�M�bjͼ4�s<ˁ��_6�أn;�-<y��mf��˭��:�:k�=}�0<#�<�񾼼18��M=i�|<��<�c���i�+�Ի���<�;%�̤�:Z �<�@���e�;�W%=Q�ܼ/�r={j�����;��<��C�������7��\r����<�'��=��eλ^��V���<Vk�Nϝ�Z�����!��F�1�n`��/���"<	�=� �;$ě�V�i�|�?��B��Ϭ�<��x=�@!��l�;� ;+�ּ���=���!-��~��6�<�Ҁ�Ƣ�;�N<��[�
ju���=�9�;C{<���iF�<z���/�	=��=b���Ҽ��k���Z=�;==&�{=x�h�^=
=�(=�K�Prr="$u�Gӏ���<�X��=�м�.T=��"��G�t\}=�5���g���C*;D� =_�o<կ=xY��׎<葁�����V�;綮<�A��M0<}�z�t{�U��;��<�I<r ��;K<e缭Uȼ�K��T:<�f<����Q��W�C��<���<T�#;ms=N�:��J�P ����`� �<M�<�L*=��< �<L��<#�<��������0�ř���7��u�=P(9�(���M=�[��kK=��X��}l��L=s�<Wn��T����}����<��U<�r�<L/���"����{'Y=~2 �6�?V <V���+�G��=�i����?�>�=E	�L��<ɯ�<'Uf=���<	P��œ��A[<�Ɲ����/u	=�<�1�d<j:=H��O9,=�8&<���<灼ٌ=�|�� 33=�=̽ �kp��4q;�6��=IA�<�z<��<E}�����:T���!e<`2�����;r=�D[=4Y��?�)<�U�<7V�8=�m5;ea�=�A��b�;cKS<�]<�xa=$=��/�~/�.�c���<��=�Rƶ*_;�g=�P���0�L0��D<[�VGI=���3<�7�<�oV���c��!���i<���ڞ����Cl[�.��i�<>,�<���=�K<��*=T�1=� =< ����;��2=�5�7`�;A�=cFq=��<��[��S;]��<�[�</�Ի3v�;������!�rU'��h=� G� �����<�$m�ɺ��O=��wME=q�<�V����;��I���M=!۲���$=J����Ѽ��a)=��K=eG0<���<�h�_���l����a<ex�<ē��_�7<�o����=���<��%�8�<�*�<kS��U\4=����
=wT*=����p�|E=��E=,���ź�7�s�`լ�XZS�ի=�����<�(	��g<��)=���<��;p�=j�.=1��<��|���1��]�Џ��=��(���u=���<�I�=���)3%;R8h<�rμ+	�<��L<�}-�T�M�)�A<��������ɼ#�r<hb���q�iѼ�i��Am�����<1�Ƽ��k=,=�\�����cDM=�G=\B�<f���j��<o*$=�=}��`|�<+�߼}�W= :=��H�$V�
�=�;�B�� <7�=g#H<w��ѕD�&�<ǃ�<T� ��NA=��m=Z+=rn�<�/0=����|�Z=-`����=��<?a��Gӻ�r�<��h�fX=8֞;-�=�;�<RU=�����ν�[Q=�&;<줪<�g@�y�����[s�j�+�p�@T=�̼������u�<j�J�h}�:��<Ѝ��Ә=��=6s�<DB�<�&�����G�P=>�(�s�����<�X�>=�A>�BiQ=���Q�<-x
=;/����2&�{{=�w�<��*<N>=%�<�ż�r
;���<�<=�>=�3=Z��,��;o�N=\�Z=Z̙<��8�+ʂ�0�e�_(=^L�A�}=,��<�;�<�`m���,��Һ�[=9D�q���a<`�J��F��pn<��<�j<3U�JO*=��4=��n;+:�M�@=
�?�}H=N�<��V�<��$=�G�7nD���!���%W�<�3W���_�<}1���<����M?�b<�L�<�Y���X�;�=9\�*o�S#���z=���_�=��!����Iϼ_�g=����0�ypn��� =��]��ܼ�����+��X�=���$[=B�T=�e=�=�05=Si�<n$s=$g$�7+=~���K=��<���r�i��`�a�\��Wv=jv!��΍=��(<��<G�#=�Yʼf�-�����	�<Z�������<xm�v3+=l�-<��Ӽ��ü�)�;Ɉ	=-1@�uN];(����y=��ݻ�z�=r����Y�?m��B<�G��� H=�!+�{1k��.6<B�)�����,���`+��"���ڹ�;�#�Ԡ��3�<��;��s�1�p��;.��'R��r݊<�K�L?<�cb����ܓ}=^�4<7jἇ��1��;�:�<�TT=����%\:��7=�/�<��-��ܶ�o��<�;�x�;���<R���<�K=�,=�M��P���=yڂ�[ե<�|�<��= �z<��r=b=�=�} ��>�; ;h=��0��S�<�3��	��v�x<�T; �=�@�C�0=��ʻ�B&�馨�h�^<V;��Q���<m�p<���{K��@^��S_=U��0=�FW���������;�W{=!^�<s�< ����{���K��R=��<=�i�<��"����յ<�O�!�Q4<vD��a�;�lK=C��<%�$=�e��\�(=��O=����I�<8�u=jW=!��;Sz3=�c1=8����<��a<�=9="ږ���<3�9�0����w�<�V�=r]�;
=P�3� =
s-=��Z<l����ۻ[�<��-���<���<r�_<D,8=��E��t����л�6��==�b�ʫ�;7�r:`�	�O&�<-�=��#�м{���:��)���1=� 
�"��<l��Ӟ�<�:=�$=D?=��m�~�G���Ѽ��#�����k��I�=�	1�tB;=N��=T<y��@�@=�Q=*�7=.�<�g�<��}�r���=�Z���U=�x �9�G�*�{�;{T¼Ώ�=�~<;�	<u�<T��<L�=��<'�S; �+L���R<;�gu������>;T�T�9�g�u(=����d[��m�9�-[=�G<=��L=g���7�;���A;1���<����I���J=.�b=���;�̓;�#o<7<���?2���>��k=[�W<W:@<�7�ex7������C<�ޜ�-���&|=gK#�y`����?<vJ���@j������8=_qz��x<=�r;��*=��(<L�7=��(<;Fd�~��<���n���Lk"=%d���<�G0=N����a��Oq=<n���h��Z�<*Nؼ;�<�/��7�+�j�`�χ��T=��l��)=�k1=u�<��=��=�%���@�bM�<+gc=k���Nt=�F;Z1;�A�8�iN�<F���3l��$m><�<?�O�Ӽ�b:�RE�<	^�<5�<�����=za;�2��;)<������ =�d���/<��k�Ƚ>�͏3��h���I�<W��<j��<��<5cD�Ф��\v9=<Es�V�׻}���bd[��?����}mw������¼��<L�H<�+=��9H�P=#�7��$�<��<�ʙ<��<���;�#i������v=~ �:�='%�O�.�mgk�Æ=f��<7O�<�F <C�;�1�� XܺU���V
=&����#���K��\J�>	8=���<7�7�X��;���������&�3M=@���r�5����ʤ<�d���9��6"��cX��>=�A��:�;�s2=�>&���e���;C��<
܅=�\G=��8�G�=�W+=�v-����<9(�<����7�<����30�����?Ѽ!w=0��<M��<K���8=�s�i���3=Q�=�\l;����k��;:��;�m���=X�_<e����=�:<�=��(<�<� =�Żx�==cw��=�Y;	�� }�;�;@��!K=��TM0�H��Od����<�<����<�	=-$�����<��;��)ڼf@=|J�;�;�S7=m�f��<Z=��<��L<�E�<�-���%=��q�H��r���9��*�;u�<�ި�"��<ѡ_�s1�>i�� ��!���.=J�p=M=G����5�<�\�����]�<�=5���3=n�=s�J��)=��c�;�]��,T=|Q���o����;v��G�����;t�e;o�	=�g�:�^=�$�y<2=<!=�mv�4W��N=�=����ȝ=8�=ڡ9<�F����=Ў<�=s��<�X黨V=0n3=��w<WԚ�|+{�|�=�+����gP�g<��G��釜<v|%=�	,���<'�r=YQ9=�FQ=is<s��<k�꼺A	=C�5���<�.7=�П;�nk�ïh��|�L�/=i��"a�;5eR=�;]�:��2���g=��&�<<F=�E=g�	�����<6���%m=Z�,=������3��w�<p�ռ�}d�b���yS=��<��v�O:[;;j?�p�O�s�;"h�����n���-=jrr<����&���к�+X��;pH��Su=>�<��t=�=�=�:$N�&�>�?�<N���>�;q�O���<���<�-��a>���<����]7:=����L�<�߻��<Ƨ��)l3����F�x�����,7��+{���廙��<6�3��4��Y	��>=�{z�5v�j��<��=t�/���H��/�<�U��$C���(�M<�����;>"<�G;.�-=h�#=�����ת<�"=6C����=C�=��C��� =�]7=�r�<h������`���e����8<�kK���-�QDܼ�k><2�{�^ =��/;�;?(d=�.7�^��L�ϼy`���=��d��y���5=J�<�73;�U�<+���,N=,T=�;�'�{=�Oą<j�V=U�{=5e�C~��/�)=�$?���U�&�c�$5�<�����C}���T=��=_Q�\�;P^(=h�{����wi���S�{|:=R��<�C�o{�; ��<�v�<q�������
��=P1V=x�z����<Ba|=���Jp	=�� =2Ҹ;<V�{�o<M=�Z���v)=���ڎA=�|$=�s:��P�0�;���ټT�=iK=Z��<zx]=��1=�"M;�D���,=��(=�����'^=1�5��u���=�綼93�<��<xR�������{���j;�ż�ݨ�WE#;�mT�N�r=\�R<�X$��i��H�<"��3Q�Y׍<�&M���
<YF����5�o�F=���[a�<�q㼺 ��#z,=����<�F=�q�'� �]ޮ<5K�<��l=�LO=X`��譊����;�;�oQ�ذ"��A�;�S�f��9 =5�<�����(��$t�<�ļ��=`i<���o<�
��a]=F�i��f����=x�Y��0=��\=�'2���߼�EʼӾ��=���<�ʃ�<�%�/V:�j���i���l=:{=�
��}]��~5n<������=/Y򼓪�=�����<�,�눖�����H=K�Q���}-=�����7�2��<���;�=�\��"�@<W3?����<_K=_$�`�@=�h�L5�̤c<<kn=j���<�=Yfϼ�AG�����ۀ�:�żpU=GH=>Ҩ��4��m�Ȼ@��<�cG���<1�*=^��;c�=�!�<�S�;���o6Ѽ?M���9W<��;+�&=����4=!���ջ���=�K="�<�D=��Y=�Cj=̊Լ+
(��Y��=�lмJ�g�E /��E�<����&mż�
���ڼϕ=��Q<{ ><,8?����<�-<�[=��/��_k�V�v�:@��E�¼W�:=qI���k���#=��I�C\�<z�)=����]���r�ׁ|=��M�^z��B�P�¸6ɞ������$=��:=AP�;*�;LL��%;"���*�;7�I=8`�=��]�4"����ü�(6=WG�;3���0 =�x�%԰�*���&=�E�E��Hw�����~<�=�{�=0G�H����Ӄ�LA�<Ԥ��W=x�o�xS���zW���M=�U�=�"I�(Z�;9)U:Z�2�D^)=@����"�Z�=��<�wk�bF�:y8)=-B���a<2bN=МP=} R�> ��n��G�$���:k&���]=��<	��$�i=�@����ȼd?�<F���	=��"=��6��_!<��P=�$�<i�2A(��:ϻ�D�<�����pƼ,��<��	=X[�<�V-=�E|�q7=}{N�\�;����6=9��<��d=��<��J�I<
�໎U=��-:��A�0����$=�_	����<j^�S�<�l���d=4�L���4�㿿<I%=�>3=vDy��HM��P/=.��<P@H����:f�@=�ֽ�>x]=|/=.�	��ރ����Ə5��;P�3%J=_`=��K=�o	�
�~;!�?<e�b�?��<T�2���<��>=~�K������];7�(=籁���<�b�q&`���0=^�_=Vÿ���C=��=0k=�����I��0U�8b��I�Z�H���;.C�OIټ�L�;�H;A�����U=gD<-]�< �!�懅�?A<u����`V<��2�Q�X=��-=���mf�.~3=�1��<��<{�H�<	F<��<���;�?����\��K �K�$=-N�v�=��!=��n�tM'�,C��yf=d����F=���;�i7�CZ=�',���1=W��<1d�<PE}=�H�=ƕ�;

���8=���<��*�ʼ�L)<��':C@8�Mh�r=�ɩ;�#=�ny���l=�}D�ϭ"�Y�����ELh��޼�N�<{8�<��#<2�^Ҽ�S,�R|i;���<���<�<�T�45�<�����<��V�I�O<���<�`��ҏk�s&ü�$��%3<p��d=LH=�L�/M�:��� �ݼ0��<׬�<�n�<�F=�ż�E��+b����p<>�#�Xj ����<CU�<�=�;�����>�<��=t�(���<��=�ס����<[~�<Vn=��O�P��@lY��?���.U,=�+k�b��DF���;����< ��1k=���;��X=��X�H�0<&2Y���)Ab=��>��<=}�<��u�oW���:���t=:�2<ه"��T�<ϲ�:�A�3F�<��P=RL7�n�һ��)�%� ��ϼs��<M�&��(/�)�N�#A��8<qG=��߼��a�Ϲ��\�;C�<��%=j�<�d=~n7�d;��[�1=�<�j@=�j����@`���m�b�X����|�P=���<�_=�ů�����;�6�S�� =e�?�{4=h��E=��׼>�=��	=������<>>���򼯆���y��w�F�<ϔU:�4����=�M<��0��&�~�4=�|/�}��p2<=;�=�M�<hª�P �<Cw�<ku =�芼O���s$R=;s=�,�V+��y0��3�<��Ƽw�;�;��Oc=�/=u�_=��� ��<�W��r��:�)1<�A�,G�����؎���=%nb=,���y?q=u(=>\k�X.=tt=��༿oH��\3=D��ۼ��=c)�;�(3��\���<4W�_V�<0�q�S��,���&=�b=�0|��@���# =a�����5=]�=y��O�S=Ӓ��r"<T�=
�E�]+
:c_=R	=�y�\��G )��6Լ�~���n%�6w������4b<��g<�)]��:=y�?���;���<d$�<�pL��><�����<<��:=Ng�;:נ:��C=y�%=��X<�2=i�p=\eH=�h���4<�Q�H�<�@�<�\-��7=��l��e�la�=��gE3�z�/=n=�?�r&�=�sA���D=ݱ��6��Ziw<�~=��D<αp���R=����+=P.=wb��%���-¼Z��J==�F�;{�<�� <Y"��ܵ<ӏ<�4�<K#�~�p�@=�d,�5]Z�*==%׼�������Gs<"�&��7<[5��1=1I�=�%�]E/=�J7=Rb��ߍ�<�m��kK<�t=��t�eHb�����O�<-�R�\�S=Ǒ�����<.V�< �=έǼ��=�j�<w�_�ad=������1�۟8=����u��X�K=������<;�;|n���a�<x�p��s#=\M�;P���G 0����<�w�;��Z=1L��5`-<y9'���j�D4ػ;^ɼ��<seq�z����O�"=��*�&��<β�6?u<���<�/s=�ߚ�P}�<�������Y�_=Q{�<�=Z���S�<��_=<���G�<n>�<[���̕��^�=�5
=/Y+=@H!�4��;�;=��-�����p�<�7,;���eܡ���ռ�s��=��<:$O=,��<�q,=�����+��UN=u�h�>]�<Xnj=7�һ��<�0��q�<�����k�nI:�տ"���y��>��ǵ��p����<1�=�	W<�2#<�)2<-�!�Ý�:�kP��ju= C��q��g|"�\�2�u��<w M��s����m%�^��!���gW��G�=��+�$�=��!��%=.�/<N�=��=����7��Y��(��8=9��L���A�¼q�b=@N_=��k����蜽q��=0��<��~��c6=�_���_����<:�=b�Ǽ�|=��i���Ѽ�U:�Oq=J�=T:��R��9i=��H���
=|���~/��{<?������W�h�_��<:y<_B2<�l��c31��_l�Ιc��Fu;nP��z+��F�<�!T��W�8�󼏪U=ϓG<�I��6JL<�Fn<������<䛞��vD�S;�=�V���<�J�<��V<��.��?=�c���O"��C�B齼�⸼Z�<$����||=���;�o�Qt<!B}<��	��HI<p'=\x��i���ʇ�6�I�6�Ѽ�[<�;�=9"U���̼�,�z���|��ļe_<;�3=�>P�8���E�����'+���ڼu���|"�<��Q� ��<0�'=�-�<]=/ϐ:������<�g=�r{��{W=��$���=�N���C�<6Zy�jb<�m7=k��<�*��l߹œ	���7���=ͻ =�~<�.��U�=��S=�0�<�P�<�>������.��ꊼ���=�!
<{,^��/=K%e�r�|�Xͼ*F���C�<�-<ǩB<�O;�`=r���Mbd�*o=C��#�M= w�<O�<��<7�:�sgX��G��[�<H&=�h�<	=QF�U��9)<"}�;8�l�8w <��8=Jmٺu��;�*�:Jxt=&ۀ=��t�[�E=�]����d���=)�S;F�(=�+Y=�.���$����,<<�ҼE�B=�6�;-�Ϻ�p=�L�<��Y���J��#�<���<x0?=vG=n
n�M=V0?��/=|��ے�k�"��U<�����<Ni���+=�q=R�P=�J|�?�I=	&�t�5��&<h�;A꾼�<�5o<�X^����<�j�ws*<�
�X�!�G�-�n�E= �9�=�{��#i<���;���l&�;ʾ`:����@��:�?��=J}-���f=$0=�=�=��'=�D=�k��
?=����n�;>�=#T="6�F+�hn鼟��<����=��=�C���>�����>���{=3-/�k��<_�Q�P׺���<�d�<傪<�J޺;��sNe�	lV=�g��� ;��==��?=4�k=#n=�*=�_=@h<�����A��Z�RcH�{��=�L<�yE��@=�꯼za =��A��<ތ�Z��<ǋ����|7=Bq<e�=P=�wf<:�h�ӽ�<X�=�/<�o~=�Y=yS<��v��G߼(�^���;��)�ء�;e�=Ԟg=JU�<&=o��<�%=4^C<���;���̄�n�*=
0r��0m
�i��</=�z@���@=S�ʻT=ɰo���P�)pJ=6IZ��3�<���D4���P_N��<���	��ȿ<�^�A���"�!�zG"���8�� �<�N�r�<�R��;�������(z�<zen<��9ۻ3{�<	��<�=c�n��)S< �R�6��<c�;��j�;���<o�Q=u����＞���ռ?7A=�	ټ{���I=���<<�Q<�Kür]~<܊���N �(p%=�:�<����B��AS=�$�<�&�<F4�!�B��7f�^Ur<�^	�<�<锋<WIܼ*�Y=�7��X�Z<Dw�+����么��3;��<�7g=p����0=5��;;S=t�<G��<=P'��=h�{��5��mc��=w�?���#��(1��z���f�V��Y�8'C<�"���a�</ =a#7<1�T=t�J��p�CJ#����<"��^M=����G�g�O��<�h7���;(^޻:�;�U��)�6=�!`=��a;d�-<���<�)���3�D
�j�Z=���S�;���|�<��[;BO�<�=��<�g=���=j�`=�T�s�ż>ȼ�U<�`I=F��� �`��)`�n�B=�-�[�̼%�һz��<!o��nt=3b��g�W]�A�N=e�#=�I�|��0�N�~ȼK�@����d�j=���<�.����< �<$}=BR����e�&ib�e�꼭��;�C�</�2<~Z=���<&yL�9�<	]9��%-����<$�&�r_Ǽϔ;�M�<=%��M��<���<���<l��<&g<�uJ
=eG=d�2�'�Be�<P�z� �2�X9L<�ɔ�5�[=����j��+��xy�ዺ;^)m=$7=��4=et�<jo��?�0�
c���gͼ�n�<��<߇:���6=BFt=�A^��}Ѽ��{=f��l�������S<�^=s�'=��m���A;��I=�gN=�
�ww��<>�G�>=!u�<��0�r��퇇<ː}��mD==�<m�M=�_d=]���;=�.�<���1㼣o�J��<���4O��k^���Ws��'�<��=��������:�6��1��<�F�����Mj=ŴU=�:�i�ż�AB=�~���b�r�*��=�L=�pO�:ܻv�kj�<���&���<n�������M�
;�=�2��
}�:�C<<}�;�� �?�;ݭ;=���;º�X]=PĂ��u�S�I��<��q��+=�=E=�(5�{��<���:�d�<[�E=�"�<qi=��<k>$�9U��X��;��2,Q��/<�U�n��<	>;<��4=ƙY<�=m:=S�w��ru����<�E==�T���Ǩ�eˊ�߁;	sn<j=�W,�	�1���˼l�W�9K�v<���;�<�9����W�Ƥ���@߼ئּ��;7�8=Y;��`1����sՙ<S�ֻ�u��CA˼�^�<Ճi��Ƶ�u�R��5=VpG�������DZ�5����K;�������=�2����û��w�&n��s�;�c�<��Y�
F�=�
��6M�Ư2�ڛV�3_��8=�6d��葺xa�<�=B�+�4���0=�e��<�#����<���;�m:=��E<��l������?�->*=<���:����+Q<#/޼Qw%��$�<ǵ<�O�]��;�	¼q-�<$��۸<��_=`������¾Ӻq�=YV=�v�|{(���a�����=���=LA��s�<$�P=iR=�?=e@0�3���`\=��=�H����~=ڮR=W��<ӤD�m��H��<R�j�ÀK<�fj=�m ��J��M=򛋼^z �E@=�3��?uN=e�м]%=��?�Gɼ�tT=,���Gڼ�n�O��<�Q0=��=�\<�l�Y���h���3=t �DRr=�F+=��H=��0=
�W�O<�R�<��:��������D�<��D� �6<n�２�<�yZ?=�<L����=-4'�Ƕռ%!F=�^'=a��<�,��G 0=��a�&Y=�m��o=(w�"��o2���*���7���-=��[����<ѿ��4����<�U��:�;�Zh��^��~D���� �z�D=�˦;n/�Ѣ��1g<�&=�R�<�>=^��;��'<�\
=U8"�Z�:��*=C�ɻ	Ar<qF(=�87=�j=f-=�+f�٥��ݼ��>��F���L�G\=`J=n�<e�"���<Ͳ;=�T�5�E=be��9����[Q�;�Z-=�2���<AD=���<�!��K&��!A=�=���^�<q��<8�%�e�<����E=t�=e�"=;=�׻u@=�"�;��z�c�X���y��K<�59=O�;�c&�6<�pD=�=(�H��<pO�<��=�x =��ծ�����<��[�w��z��DF�Δ=�;N�:�x=���<2?<=y�d=��=�eI=Nmݼ�l�7�T������@���1=S�O��pb�;�a�%�3=��N<�F#=l=9�������jr�=����8;=/��Oj�@ǹ;��
=Е�<e��<1]=�[��H/=�5=�e�<*Yd�0Ỽ�xB=�<���}Ĥ<5�a=|�F���q<��m�e�C�N=�'#=c���y�J�/�M=�v��)
U��D!=1��<��"���Ǽ�=B����N1��6�ud=H���@=T�󼉋���S�۵a=0��<RYL=��B=$��=�f=��!=�Y���Ƽ~}�On<��p�AK= �@=��Ƽq\=�n=�q[=Cz7�ԑ��&˼��<��U���{=��
=�/m��y{��
��f��=Lg��}<D�׼�	N��hx����)c=xp���b;���<�G=-t���5�c�<���k�=�Y��e�/�Ue7�:���P=��;��i-=��u���ȼ���y�=X�Ӽ87�G��U��d�w=Se'=J�� ΁�Z%2�w�;=�p*=9P?���B�l*<`��=l.ϻ����w~=�0<�4w<�DX�`�=Ws=P�5=Y��<�W-=����օ=Lh>��jɼ�Am�0��<`X�V�<�h*����:��<B!<'b��] ���<k����;/鰼gS;=]+Ƽ��>�O�F={�ʼ'���Ͽλq��p�<--I��CQ�#��<��+=�S:�}:�<a�|����<a�k=�׼\p�<JO��v�	=��=wY�DL�X;�����9��=�VR=<VJ;�����eW=F[�9�*=�B �0W=� v��M=�;�<��v�#2z=���<xyO=�@<�'μ���$�;�c=�������<�x=�r=�^6=��<79<����:I.i=Z�F<!�_��+4��7k�Zb�<#=��j��cW���!=�ʆ<+G���0%=
9Y<����<a�<Y���k=}��<�U<c1=և<+��ܢ��\+�����("��WR=!��uЍ9	TM;O=�<�D;�.=�QF<e=ܫ2���U�r��
p��=���h��ռ���ްY=��:o��<�N޼eI	�����b����<,f���p�<��<��!=�k�<Nh�~�G�;4�<4��<ې=��U=|�*��״<Cµ���<'Y-�� ���#='��;C���T�n#o��`!�Q���VR�rɅ<��ƻ�;&�oi=�e
<
�;�e=6=J�8=��:�W=�?��B��|h=��o=U6���4�<[��<����Z=ιG��s�t9����g�<�ֈ�c�=6�>���0=�J�G1��.�C����<u��<���<�μ��7��ņ<s�C��G =�N=��&���K=��<&qG='���/"���=���=A#�t�ӹ�H=�����<�+�<c�/=\�<Ӱ=;5JT=��<�@�W���K(��us�Ћ(<�J����<ڭ�;��z�A�<80�<�7�<���;�����a={{�U�����<ѯ)���
�g��Bi�<��ļ�	7=��4���M�@���=y���)�	wͼ^	^��������I����:��'ߺ� =�>M�r4!<5�Ѽ
r���=B��H����������<��=��/�t,�;e�1=3�>��=ƼCb�<uP=��;?=�}�;��<��(=�V�����ϼ�]ús�P=�E�[���`�ü��=��j�S��+=��;)�#����<�Zr=��9��{d=&�@=�\�;��\=��\=ձ�<��<�'<BO:��oA<�:�CE��Gb���J<�=�Ue�\����h<��v�_���+3%�QQ=��S��#�ۖ <� ���m�	l��V�s=2�Q����3�F�NLv=�;�:���<:)g��x.=���:�a��| =TW_;�<�<~?�<�m"=C���߮`=�*�%I�J��;��x<Z�!��<���;m�л?E=�w#���v��k<-�J��f:�R�=�J�<���;��s�|=2lX�[�=H�N��!9�봦:^Di=���FH|�=\�<%C=G;=�wм$
�&�=N�[��k�m8<�M=`c=+�1������nL�-��:�F;<)#�~����?1�F�Ｓ�;�L���I=1*�������t<���-���L�m=Kq=�������S��G�J�;+:�05.�$�}=&��;�r#=�N7��X�<���;�!�i9W�Y�<s�l��a]=��@��G�@�=Ϝ�<l������锼�4=��=+!��j���/MW��DƼ�=<l�<ܱ�<EC<��W��<���ȼ |d=+઼b��<t����<�j�p
�g綼-=�m���E�����>Aa�v=������-���<�Nݻ��������=Y���2����軗*c=�T�<�
e�_bA���,:��(=��K�{�c�΢ػ�)�=���<]^����<?|P��=Xp��/:�9��X���<Q�`���;��=�񤼒=9���,?:��>�pc6<��K�T�<� $=�Ӽ�<k=",3����<Zm�<p�=P`���^��LǼ���; ��<C ���e�ҧ�����)�;D-!�k�q<{�L<"�s=���zp��ɁC��	����<$f����K=�=�7k<����Z=�F=��<Z��<������\<ÌB=�{��e�]���r<s�<5�;C� =d�
���h�<Ed��^�K=��8=g�<&=]m;=����S=R� <#--='>.=�¼�K����Y=}ca=Hx�;����5�»�"����<�E1=ąټI�C<P�<�+=��=�Z�[^ ������Sn�&O=' =Q���L���9��O���)=}�&�qT=	ռJ�a��ЂX;If��Qd=�a׻�&�l^"=���<�"<I恽�)���;�0&��O?���C�W��<&6���?=t���5�N��;ЊB=j�|�Ƹ�<_���M]���;�X�o����:��+ߧ��dͼ�|�;�M���4�x�*���c�<�=E��?�����L�gؼ5+�4�=��:�a�;�H�<�d=�/��6�{�=�E����<������n<��<8N|��wP�Z�����U��;=�>="�[=q�)=���zW9��)���y���<Z�1��=�C=��<.ns���������O=�2�<JQ�<eݼ����F;��;�_=l<<������>��$a<a��<� )��;=����q��<�����!�'��/��\�V�f�Ɗ�<�r����3�V�d�;�Q�<��=>h=��j�����#��r���?�<����+>=��;H=�=Xa�;i.<�l�<��<�L�<V��<�����u�ӛ
=��6;[��<E��!Z=s��X�;�6G<���<��j=���<{�y=Hl=v5=�q\<.\�<�=��<�G5�#��<�V8=;f=s�-���_=a6�<A!��W'�X��<&?b����<נ*<�eG=2�5���<b韽��g=�!�E�ݻ�)=d
2����	~Q���+�sB=ƻ�:���<zA:T=��;̊>����<��:3��<AR=	*=]�]�	���َ���f=²�<a"��!�:�Do�I|����<���<�`<PЊ�)�<5N'=So=1dh<�>&=9�V��G�����<��5�).<����yV=i�<U=�H�U��<WJ;�cj�B��;��W�d�S���u=�_e=^7� P�<[S1<��6�Oz�2�)=Hk-;_x	=��1�0<�82�@�-=�L�6�X� �i�@�n;x��_���z�<�[�<Bn�����2��}=Y�¼��D;FB�:-�K=C�a�$#V����<S"���,=�16�uJ���Bʼ(�P=�T�<�D2�ax	�@$�o�	N��"��e��<����˓:,i��|<<�=�|=@�B;r�e<T�O<	J꼜mT�>��J����&�W=egX�
h/�2�<�V�<<��;gu�:?�ü�LD=���N�|��$��������== 7�<�hݼt{]=�H��L�;8qh=3�4�ǟ�̼��D]��t}�Ҡ��?��B����Fm���	���=���<�>1;�$��1;��rr@���;���	 ��(g�j �c	��=Q+J<��0�������:��cc=v^=�zѼ�1=�w��0�L=*�&�2$x�X�@�,7���}<7�)N8=�v��O&=������|&=�RD�E�]��)�d��n�B=��5�LZ<�z<8;�=붴<$���p
r��mX<EgO;����5w=,;
�#_<�X-=��ٺ_���a���S1�NK =8�B��W���&h��64=l�<�/��9F�[�<y��<�|�5�,��}�h����u<oh�*d�AQ��,;?��=�0-��H&�&dE=
W���2�Q��<3k��$���6=��^;�ZS=�
�<a'�F�N=)c�	K���׼2���#�]��</O��GZ��t~<�6=�(<��:����k���ؼez]=�NU����ɼ{6�<�ӼeGC;��ܼ��w=i��ؼ������
0���H=:��<�Ѻ�贄=�!1='�ż/�"��ea�`�O=+D=�E�"= r=�=.݀��z�<ђ<=Rl��=���m�Ƽ6�Ӽ�=��o�b F=��;u����=k=xB�2���~�/=��<���;B���(<b<��9<�����h��7=��n����<(�=\�����=	1���c���S�I7==�R�X�&��Ҥ�&Ｐi=<�(R=�6ȼ�e=��*=�O��q�5�DcF=��A�EjĻ���<!>;<� l��k���<�B����<�_N� ��#"Q=(S�uA6=@��;�T�*�\�\��<y��<����9��ۏ����3��ּ��k��xU����: �=���<�[�<a��L�JSY<�U<N^X�N�]�<O�.�x<A�G�H����p8<�7A<�X���=����h�V=4�=�h��t(��[E:�����o=+	�k��/�V=�Y^<��Լ��'~=�BZ=�����q�8�<��E=.�=�Eļ�ȼa��.��oX=7�3|!����;��M<r�'�D�K�>��;2_=�~K���e��p ����l�N�!U~�:�N�z�$<�<�V&�2E7��r�<�6�0{ <4�@<I�=�5W�l-=�(G�K��r;=ɜ��O�2��a��6�b���`�;�s<��<��s;3�@�2�b�#P�XF<�kϼ_;J<|8���
='�]���<�JҼ��4�PE=%Y�%���<�#P<e� =&��6�����=~�O��<N �9;\�a �c�0�ݻ���<��K=�pA=�[=E>=��U=�"=�%���U=�6=l��5A;=�Bs�.��g�K=Q�;=r_d<W,������G4�<����<�-��:��<�
��˨�<cuh�@��<���;�h=ة���:=���#,�p��@x���.�;�b_�����-�{q㼎�3=)r��{�P=4:��ܣG;�4��<:&"������b\J�]p����H=7�<'� ='��г�;��=<+�(=z'������'={LԼ��=�b<Z�'�؀���<u�B��p�ڳ�<��ݩ=�A�ټi9L�[f]��X���&<��{��A1�u�_��
���|=�ߺH#�<��9��@=c�l�=y0=O�<�ra==U���:��<�oX=��:� �r�)�+0G�m�=�KS���;q/�G��[���N�<��5=2OѼ4[�c�M�Ө�<P7�Ű��8A�;r3,�����D�l�b=:�!�C���<D<�>p�2&-��y�
v �T1j=ʡ�:;0��O�=����B���S=�?&��z =�B��X�<�G�~:�;PN��C��ޔ)�|�=û;3�&=�4=�9�&����R=QHx�'�%����:<��=���<�O0� {̻�!����=Q2K�%oc<�J���1�8q&�"hn�ʟ:=#�a��,��n�!���`�C�6=RҼu�;s��1I5����<&
�; ,<�%T��3��C�>�μ�������@�<xu��̦�<7a�;p�;�I<v�+��\E<�b�L�
��9��#j���3<��A<T<���=���<E�==�����
ɼ4?<9n�w���Q���*Z=F�=D�'�����e�-/s; �M�j�,l�=����=Sc<���)��#l��=��<���ǧ-=}��;���;o�<�+�=+���P��<�<eK=��O=����0B���M��}@�p��;�vS<��=*}v<���;��&<-=aC,�ˠ�<m{?���T=7��<�)=��߼��Q<U7�<��k��32=�7��ȼ=�=X���k=|.�;���Gм�P=�W�|�.=]�X=;T��?�<�2�<���;�R���<��=o#=���:M�<��D=_`�<l�߼��C��=��C�*m
�s"<���i=�]|�<���g�ܼ��1���P�ظ4�=D��-��0�� �C�o�`=���;�D{<��A=�O=%�C<����G�<�!��beo=i��=A�W��`d��Q��_��L�a=�y�<N�d��7:����h.�<!����C���<r�=��=>�:=y��<�G��:@;�`�<S�Z<0̊���X<e[.�F]�������<�<�Gv�\�|����;uч��j</�ͼ��M�s�=?�ϼ�H�)!z:1��<)�n���H=|��<VB�;_*�Tg<ii=&��R��<��<%Bs=��<)�K����;r����<a>e�m�}�*%�<ŏL=�Ȼ_�߼��⼡ߢ<A&�G�ü(��<A�S���8�y�_��X$>��休�{�=h���o*�;�(���E�C,(� ������;؉�<��=CKe=W�ٻ&��i�==�$�&�:6=,	f=�wZ���2=
G3=x���U�<?�<��d�I<����O=ޜ�<��O=��N<.�W�M�2���<݂��T��<Z6r������t��F��cN=�] ���z��(�<c��cH�<��8=y���3,S:��z���=�|B<�_���9M=ɽ+�v7E=F�=��ƈ<�ϒ���'�ݼ�^�~�(�q7w<�I�<�Y.���j�$�<�[=_��<��@=C;O<���Y:���)=�M�<��[=���A�~��ҵ�Y���E�=�V=��ټ�L��1���m{�L���!��~e<�/��,����(��qP��ZV��8+=�l�p�R� <�L</��:)0=�v��9�;�;&(<�ܞ<�[=�}*�х0;F�`=뺄<�;=�QS=�-�� ڼ��G��� <\��<�L3<٦�<�&U�!aG��R�W�W�\�<O?��*a�<�5��_��}����HI={�<�s�;��1�Yn_���<�_`=g� �(��=R(<�F=��O���<_W�J&���p=��<f�,=�m�<���M ������<O�"�+3�=;�Z=��O=-s�L�m���/���[��J�<b9��F�b�g��.v�,4=��<���;Ԗ<�Ҍ��Hc���<3O=��P��G�MH\�u���3�;W�<��6<�"=��O��;���_&w��K绶7-=®�<�ڠ;�M)�fX��z����̼�ہ�1&�h/w��-=tA�<`M��z�<T��<V�9�|���{e���;�H=��;�����-m<2{e=�\@�?�x<�pE;9�T=��ݼ��B=#�#��J�;L4	���<��#<o\<��d=�C�<"�O=-�h=3wP��B���r���L=���=)\�<�=ϼGO�*����M/�))t�9�ۼ;�����<�����g=Nk�<ݻĻ������<�ũ�NV-=�m�Cj�=����<=�3��`=6�?=�4=m��󤇼Ȫ*=��ݼ����T＋�N�g��;K�ͻ"v<=t�+=���ZO��$�;{
=���`B���B;Z�W=��;����ǧ<���L!<���<��=�����:|�˻0��΅u��6:={<�c<�1��<������<#?=��<���<��=<�^�ivO�|��F	�]���G�E<ψ=�!+=�`m�R���Wg;W�i���:��&��"�<a�M��*�;:=8�=u!=@^-����<
Vj=��Y���7�r�<5L�=�Km�̣����A�Q��U>��X��� �bj����G��s.�ֲռ���g<�м|I���=�2^������;��!� |A=��C�y�˼�r=�Q=�k��'ƻ��ּ�Z������m"N=���N��<
��z.<�)=5#��*.����E��l�<��;E�<�t#���$2�����<��W:�
X��4��x�U=�g=����滆�/�S�i=�(=��Z�m"I=�Ɂ<f��<��I<�1c=��;�=%ü1�y��쒼,��;���&�Z�ݧ<��;�
l���:��0�䉼�Z<8t�>��;6�=��L�I�ۼE�#<�;���<=�wZ�<6�2=�D\<ߝ<mN=ȑϼ\�<�b=А��p	=~S�<���<�]f��9<F�u=g9�VR���r=��<f�뼢3(=a�8�p�R���S;-Ĉ=�(����k@=Gl ��|!=��7��VG=��; �¼(!�vF��i�=�+�<4K� -*<
�O=��b��q=ҡ$<�m'=��n����<]˛��%�<��<p�He�;�s=�/�8�4=';�<ĕ =��'=`�X�P�#=�Rl=��Ҽ��!��/-='�<B-=�ɉ=�`<=V(Z�@n<�ǡ<*t�f4<d(<q����)�;�=�<-���vd�<�V=����y�h<�վ��xG��=�Q�$=`F�r��ɧ$�
湼�=ÄK={4(�T�<�<]�U�;6t���ȼ?	Z=�,(����<&�	��B�;�q=����a>���=�L=���H��<s_[����<����=��\���Y������(=�<���=9|P������;����;?�^���>�ā=�7�E�?�ȏ;>�X�[�^='XF=S�A=��<(TT�̯�^%��]�H�<�WZ=��ڼ-�<�"�<u�8�%���ȵ�<�\l�=��;�-�<��<`=���<�]=�x �$7#9p�c��x�ڶ<��&����;�	Z�rS�;����<Kټ-�����;��<�5"=�Y���;�<��ݼ~�=[��<�]=��|<��.=y=�t�;M�<�"�;��7=�� ���f=�z���=���RY�V���a�<�6M<ȍ�;I�S=�Z��{�;�Ֆ�����,�%Y<���'��<����A.=��=�g=���o2���D����e�)=�X����ۙ;q�=࠶<����T���<़l�E=}�=Ɛ=�;�Q��t�z=��P���;�@u;�!�<��E=�?�}�ͼ~��<;�<���<DJ�<��5=����F�;�A����<h��<C�;�����p���� <��R=��F=d�D�5(d��v=�"`�u=�*C� �`�#ֶ<Y�7<�߻��<��<��v�l���<�<=��<88>�9=D�;D��<?^��0yƼ�<eq=�1u���n=�����:�h�%v =VMX���>w	;Cq�<Ԙ;;�쟹o�z=$�=۾��6����$��6ػV�����<W�6����9�1P�]����[�\)���CC��{k<4$a���'=c;>=ޒS=��<�xS� s�;�=UJY���㼉��<�p==��F�~���;�=�~�;G\�����V��TF=��	=�"���v<�������P�<L�S�l�<k(��"zI��������0�.�#=��0@=�S~�^<�<��*��a��L=,��<��T��<=�z�_���<E6��(h=�=8c*=/�Ѽ��	=P�5���g��{���4��v<yZ���z�;��><ڑo=ė=��n<���<3+F��I=���N�A=x-<�<X�<]�=W��<�e,�e6=�� <Z`P;V3
��<�!������<��7�H-`�ޣ�<u���4�B=��5=�ߎ��[9=¥,����і<�R5=�X�;!�4�=pV=v1��j.<�D���W:=9J\;I��roԼ)P�A���/(=�Ĭ<-�O=˦s���:�����'`�藀��H�Ъ�;4�<&;<<�u�<����S=���Uټi�ۻ���>;��pA���*=�Y-���Լ�M�<����/Լc��s{��$F=��%<6B�G�.����<���;!%	<��<�����p<�"��c
�(��Q�l<��u;�N�<�Z)�]j�<��;�F�<�<�<�c����.�]������=��d=6�"���J��<�������/C��Dp�k�g��Ξ<��9�܈�<��i=�`<!�W��@;e���x
���(=L�<�k]=���<��`��;�3胼w倽G�8��r:xx�3��i=V'8=h"=?0�;	��<�+=�X���<���<�=��#nE�<��&Ծ��и<>K��~rn�������;�2=�uZ=�9q�I�˼�9��C)��9��Z�<�"�<	*�;9����!=E|���G���L�=8�g=����P�<�
= �X=��T��;'���;{=e�*������W=�"g=K�_=��O��p��ܷ�;�98=��R=��(�Đ;�O�<�*o=%,/��s�<�<�?����-:=�}	�:�<@7$=+=�O�;�5=��V�� a=A���b����G�w��<�<��<ص8�a�ڼF�����<� =.�&��o ���g�<�H=,	n���2���z�C��U�&=��8�~2'=_��<wIݼԉ����t��[=�ĸ�Uf9��n,���;�	6*����<��A��ɼ�l�{qJ=��k�7�.�ޤ�g��iJ�*��Bf=:�Թ-�?�c����^T�R�=�k�<$�<K�r��^y=�ƅ���<�$�	J'��aS=a�<`�6=�p�<,|=�~L=��)=��<��<?�=`�R��� ={���[��Z�ԫ#�}�<��<}&e�b�a�P��5�мM�&����]�]����<pfa=�	���Ӽ��\�eOB���==�~�;�kI��[g=��<��P���(<�3�<!�����;�G�,��; �=��6=F���Ka;�ad��ۼmH1�?�@�Y�;U��?�= ������==[�<�v�<����D�-�U=%2����D"��^7�&m�h�<p�l��@�g�<�&�r��<�E=3��(,b���9<(�h�TF��f�%�R�U*���<�g�L�i�)Y���@ջ.��<�ۼ< ?��w>=��T��=V+ռ���w�{�$�W�<������+B=�i���/��Ke�f,�<�_5=��e=�l-�͚�j��:�9���;�<��</���";��et���=>H�����<�0�<���<��� L�<L���R�<� =�P<����;^H=ƢB�(𷼑32�	m�qa(=�=�H@=�Nc;z���l(_��F=A%=�F2<8Q��b�s��� �⟝<Gp<l�U�:Ѥ8�  �<U�=��
=��<����u��<X����:����:=�v=A#<}c��t����˻��k������,#�d�=������%=ay.<R�=㱣<i=��\=$��f]=w�u�R��+����Д�Mn�����<V�<q=E���U<=�ј��۝<��K=��d<_^H���<��C=s�B�G��;@���[ l����<D�<��f�N,�;�9���<�U=~�����4��N�eo=e�����8=�L���=|{`�k����=��=�4���Ǽ���V�<L��<��<��<�\�5��<nz�,�:=�RK���;���[N=F��z)<u>��Rf<�}`=͚�WiU�A�'=���<KJ7=���<�5<g,�=q�;�X�uT.;���?=���<(y�<=�}=w��H8�<�` �8�ۼ^�:=G�ɼ�=��<-�=�=h�<�9��-J�j�Q;d��G*�<Ҫ;���<�j^=&	�ܰ�=pqn�Z�[=Y��}S�<��W�"o�<ݏ�ƮC��^�<A��<*+=�=�(�<vi=W�z=K�7<����А=B��XzJ=DC=�3�<==7�p,=�u�<y����.��+=�Q3�(z==~��U�&E����C�v�P��e><��(6=������]��	�+D(�S��Z5$�2Uz�WYr<w�<$C<�wI�`�ü@=�ם<aĀ;�yw��8�:�Q�ǝ����<�D�<�o�, =y=\<3�=p�]t<?2�<�3���R�_�<Sq;�}]=ll&���(�F�#=k�2<���<��<<[�~�:�j��;��=|9R=\��hE�I>�Ǜ�<��;��f����&=��T;"ڡ�!��P�	;� �<bh�x�A=�ʼ�Wc��8���R����;G�J�q���k<ޅ<��R<�nJ=fg5�o>��x�D�I��K����:W"=����2=U�<��E�����l7���r���D�^V�,!7=����@��#=1Xm�T�����=R@=^�R�T�
=�b�|=���xo�;�9=����,I���d=��=/�)=X^H�������w<��>�� <�r�<wY¼#=\��c�k�M*�R��<�QY�R*E��D;|�ɼdj���X�<�Ǽۋ<�I`;ZN���7=�:�C�=��8�kڼ����<�;�
=7�����=:X��!�=6-����_���@���=�Wd<���0�e<��I<��o<�tż�����<*�D=�����<�$h�<a�S=\5{���-���&���T�'!�<7�N=�'<�m�=��Q;��O���"�z�H�5ũ���tj��B�<y%G=D!ɻk&�z����砼9�<��<֩�x��;��c=��[=j�o=�@=��+=Xdּ�4�7P�RY='i_<��D�<��<�I=����-�lnd�+����=�X�;Kq,=��S��$]=_���U�<�0����P��;�t�4-��[�-=�z8=e���L����<�3?��I��[�;#~�d��Uq.�V�H=����wiʻrl��{A��"�<�I�����]�;��ļx2����y����u{��V�"�>=�G�_K��a� =�^���4Z=�XZ��=�y~= ��< ,��l9�<E����s�<��� �<\I�2:�;޽]�&ǚ�Ը��*�<�M=�ϲ;̫�<kT4=k�J=tr�4���+=�U�7ZP�%=��7=�*��j'=��=�������˗����<=;���O������;kP���2=*G=Ҝ�K�A��p<�C�;�˼A7�D�C�R':/�+��w�ՕƼ�U:�}"��q�Б����żE�	�"��|J��hǼ�-F:ih��zP=��
=�z�=�2��P>��?=|�.� V.�������Ҽ��C;R����u�=�?�<,a���%=��U�%������-�;R�ǹ��ؼ���;��<-�; �;zw׼�����:$�#<�^=,*a=�[K=���_���&=O^�<���<k_����}���m����;�-�;��ټO=��缅V;=i�<{�w=t%�d�E<���6}�<(�;?͌:���sZ�=�5l<\��j�&=BT��֛<#A/�����4���7��d��<E�y���=�7�j�"�u	_;�m�<κE��X=Β�<48��?=�nQ��ZH=L�!�����TP���)�{4Ǽ�8D��v�;���<<��<$����3���<��<�:;q[b�Zy�<��<�3��G��+h<�-?��B<��ݻ�o���R�<��˼�@����
s�<&e=j </3�;�����}��U;���<��4;]��<�n���<�i.�����#r�|I=~�?=`�=ۻ�N��u��<���7�&�&R��󲼚x�<�(���U<�^Y;J�?=	D�<)����;�8�<\,O��i=ݝn���N<=2=��D=[} ��ܵ� �$=O0=y^��!=�9=��b<�D6���_=�R�pȼg��;�/��<�)�
[=p�<�㟻>�<m����#�:�ϑ��˼�<�<�t���=.�%�d�=�XQ<q~軁�b<��)�͒Ƽb=l��<���<�
 =���l&Ի��+�;�P1�Q:�<���<9�S<�<μ*��<p٣��o%=�J�_�=�7��x<Ua̼W[:��t=0F�<��x���*�a��������%<v⳼\ƃ�q𻜓};.Ǆ<��6;�7q�+<a<����م<�-b�ٛ/�)"=��<5-g�\ U=��=<w =bgh���ϼ5�T�f0/���[���d��u�B���=� =���	.��$V�ɉ.=���R8<�=��-�:籼��������`�%���={�8=�_��� ;�$����~
=e�%��i��&O�B�;�V�MQ�8�=RX/���׼�q�<�@?<ޕc�Yp��S��<���<o�=�z=�|<��=x댼��c��[~=��;S�.�N�=W J�_�<�a=�x����<O�=�����h�����:���<�n�<D��<'8*��}���!=ڭ<7!�r`�(�Ѽ�$9���T=�$�<����1?�<��E�S�E=
����t�?SԼ���;�,1=���;�<XA=͘=��)��tL��y�<ţ<<��<���]�<s���n�h;�L;F`.����<����J=�����w�O%A<D��;� .�RyN�?%�=�L�=IUO=�&]�Z=%��w1b<������Ҽ0#�</�ӼjY�<��@���4�T����<���ےO���p�m�#=zZ��e�<�q�;<H	���H�<e�=<��o=N<�3�<��9巼?<��m=����Ӊa�kY�:���<7�����g9=���<w�=�4��FM;�����=��k��	.������<�aT<pU*=��p=���#7C<b�l<�n=�0��=�<͚�<�6�<W,<=������Z=ӈ`=���:s�<�^l��7Y�]w��w@��c�:�V\=;7k<��':���r�,=�����<��󜼽r�G�;ȑ[���N=lv����λ&�<��u��������IXF<�����<���;Ы0�(&;��¼"'G<2���i#;��;�@�=7��;��-���]=R���ƙ{��7:�ړ+���>=C�7���߼j��Q~��29=�yn=S¼y|7=%o=#�⼋�=��;lx���z=��G�����e�9=��k�n�9����4�!=��<G�W�EN�;�Sl;�&�<&B��
=^��<$����=��Ŷ�J�@<yN���\�:�g���4e:�lr��vK��4k���_�d�e<�K�<�⃻"�
=��\��J<-�	Y=��j���v�>��<͌=$|�-G�;��6=�JN���n�h(�<1W=x%��4#��:4v�������}Q�xľ<!C5���D�c�Y=�Z<o"��Z���=��Ff�e	��`�<!?=f�a:b^3==1�e�8=�0=��<Vk�� =nEɼ�=�x=B�ۼ�Ȥ:k==cY�����p�;d�<O|B��e���ϼ��!�́��Hx�	�f�W�X�vѼ��n=pI9=��m���<�G���R=sPR=^���D�߼��<�	��=��>�����V"�7?���;HL=�=�ң<�_��Y=��.���=�cκn��L�<���<\�<���;�/��{�:(�;�$�:��R����<��<c==?�V=�"=�E¼ח3=���m�<itl<[ab=4d1=�/=P�����<v\<�ϼ���<e�=Si�<Uo��L[��l ���<Z�"<Zf=L�ӻ(�=Ru`=kud��|)=ߍ<�AǼÏA���Ƽ��Y7�Mh@<���G����7�9�5=↾<�G���t���X=N�<���<U'�r�4=��<j��<,����mf��;nf�B���{=��+=��:���=��J��⼉��_�Z�o�<S6c���μ"���xc=D���b�>jV��c-=�\�mwѼֹ��VɈ=v�7�mP��(�d}:�QSd=�6,=������m=�W��>�;�2=���=qʁ�GH=�@y�L�;S+8<�UB�i�u���=�#��';�K�<-eݼUd��MI$��0�3�B��i"=T2�8ݵ<ܻ<y�	=!����<<E�;ue��=��8��i�7=�����;=-=�̼j�<�	=g>Y=�gs=��q���S�̺�/@�:@��<ǐ<��^�}�ɼ�@u���<P����?�����<�T�;Da�F5G�9:%�?,c��p=�ɘ
=��|<>�N�o<�AB=9���Rx�<)��o�>=j�1=ɸ^�����!�;!8��'.��ρ=X�u;+�@��!W<f/9���G��;�[=!d��])D�4i���%==i�<�i^���*�D2b=_S3;�s=���X�K=�CZ�G�
��������d0����<a5�9�{9�r�T�Z�������ȼ��:�eC=|f��n�<��O�k;$Z鼱�K=zϋ�����T��=�Ua=��u;]��<�����DW��P��P�-Jc��� �
D&=cN�X=;� �)�ǹv��<�5�<U��X��$=n)=*׼�uϼv�'=
� <��A�J��E�;{s:��@=��:�#.=�*U=�4T��-�����wa��� =�Ɔ;����S�<�;��{�6=S�<�e;J�t<x�H�?����7UG���<��L����+��߳C=�6���r�<���͟C��%�;��$=���W,=L/;���Z�<_�e��VQ=�����:�[�<�C2=�7�;�+�<^�9M4U��$X�@�/=�RG=	e��ƻ�u�kH<��r=�?L<̴��*�;kcw:�m<����\��I׻w}E��eu=�,E�[��<��a��;�����<�����<��ȼ @=uP1=oLL�RBh��� =�QF�?�'=]��=�b=�"m=��4<�AX=A�"#�$�=�L�����������<�Y=�a���`��K�<�G=��ü/mo=��J�_��Utz������=��M��/=��?R3�К�<�˻z�#�i�ȼ�8�1q�<F����+='�=�}]�����&Pi=v��;�i=~ M��]=��w=�����7�t=��U;���;���k�< �<��=��ټ�\p==���_Q�pn�pR"��gL���=ĥH=4Q���X��	P��v�=��w=�Lf<�g�� �K�>�Q�%�:ˠ]���ܫ3<�"�4�^��������N$=���q��=|��: <�ꪺ����
s%�I=ܢ'��F�<sjo�Kb<|��<�4W=N��UN7���X�E���T6&�͛f�V~t��O%��p�<�I�<��<�`=�J ���<ϿF�N��<=��_=���<�jB��]��� R=�<�NL=OrT<G��<�M�<�J=1�O=f�<��o��I;��yۼES�<�����@��+��W�SH*�٬��r�ϻ�JO�l,��	�<I�ͻ�s;�K��J����w��U��< �h�)�n�/b;=�ښ;9���eE=��A<�e=�����0�$�<$pp�A�<5E;����<{�=�����Y��Z=l6�<�Ӑ�6��<с�<�
=d-�<ȴźP�<�؊<np=�oE�M[�D 5=;�<�4��'=U�<����"=�cѼo�,�1P)=��{�l�=�|^;�(5�s��p�2�3Ez���<�}����#�W%�<�BZ<k�"���=uw<oۻv��<�u9=�c�#�Ѽ�}�9�8�=��6���{�ͤ=}��fX/�{��������)0=\��<j�]=jU2�wM�ldo<��	:��3=<z�<3�<J��<�z=�#"<:��|��:@��<��g�<H��<
�:=�B=�L=cļ�9�<��<��.=�~��a}~�u��*�<z�U�|�d�r�5�� �;<v=��¼=>3�Zi�<�EC<��J��%Y=��t=���<��Q=��s���r=��K��"���V:;��'=�d<>W=!g�q�\=���<���E
��[ʼo��<D�ƼLoQ�g2�</��<�w?=�<v�Լ+�=��l��,�������`��Oh����y<hY�o��<8��.��;�Br�M1=D�,; $A=:�=g�,�E�l=8/Ӽ��=~=��o����ϓ�<�
���nL=�	,=�������<[�üg_�<���9������<��ͼK�ۼ�C�<�uf�ڴּ#��<�ݢ;�����$�<jB�<�	M=s�1E��"���P<Y��<���|)=�c���2�<��I=���<�^�<�x�=�k�~���<�)���?=��=���3�=��=�N����qs���f=������=3�c=��<Ä�瓤<��=��� =P�u<��<)��;(�E86����<o.K��=L5�@�<t�H<�q�1
�ANA="�(=�b��c�����< �L�<�61��4s�0;�@4˼��=��l�, ��l�p=���<Y��;�]X=�q
�����#������v��=)�]��C�׼N8��7��<��K��WF=�.=?���Q=h[�<]�K=]�K�F�V<ʚ�:|{����;��)�V>��{�׼� 2<w"<�V$=֟�<z�a�v}�v��<S�<S�o�s�ڼ����<-^=�1�< L�<Va�}W�<��<�6���:.=�(�;c��"���a���Q�oF��T�<PVD�M�f=�����H]���=#�V=Ǵ=͓�_�=b�Q<�����=�S���6'���@=Gͼ��<�����<��<���;���;$b��y���9�m<��=`�<#En=&�c=��廟�=��<�P/=��-�C'+=��<�?@�|��<�`��FQ=�rI��V��e� =
5z��Y�L=�<X=~�,�f=����G��<2%��[�;�ۻ92�:��1�<0��	2�a����i�qw6=�TO=������;�	;�;	w5=^�F�m�3�wt4���7�~t3�KI=��e�h<*�������<�`��2����4���̼~�<�	�{
�<!*�<��<�O�s�����Uܼc�O=!s�<���<�����Q=�	=g��w���noj��ܵ<H�;��/����<��<�=B��:m�7<i��<b.�<"TF<�M�<v�_�0N=\uO:��=J�F�a�:���1�ޜD=�z�<o��^����6��=V���n�9��H�f�<�'���v;�"_;�&=Z�Ѽ��<k�q;=	�鐽>$[=Ô��Ov=�*=ǔ�<@R��"��=��
�ԳP=��w<��R���q��>=1;R=h���\�<��=mv��߀���=&�S<��:��\����<�r=�^V=�$�w"V��<�^��3�3̉=Z��9��8�<q�����<"�<V<�K�zP���=�W]�G�6='
]�� ������a�=x�n=�7���K�<����@�Z���X=.h�<߾6�����c�="��n���()��<�=V��<oH8=�58�S�+�6\�<�i-=�5�;h�\=��ػ�R�:��=�;#<x����A�;�&;=��I�Z�p�[�	8H��<���<D�=�o�,��<�2=&�=��j���)2:�t@=_�����Ƽ���; �=�qk<���������<z6��kA
=��:�ȊԼ�q�A<BE߼�_�<;� � <�,�<�=�]�"Ig=�cJ�sͼliż둩��#��
N�ښ:=��ȼ=��<r�;'�H��e=R� �p�#�C_t�QϚ<)<Ż �;��q=S=_=���#ռI�;g��;�` =t{�<(�<̓�G[J=����J�[T�;\�:%��L�(=8=�<?u���>;��t��"�[=�v�7�<F�=\B;4�<�==aR�;�L9=%x�b�<(e��-(X=�8$<K��:�ZW��T�ޤ�޼٪�; �<=�Ff<�$��~��S~�<u�ݼ�l=� ������r���\]�2����������q��`�?��'*�n|=�L�����7u
�y6�v�Ἥ�n�Y��<��*=��L䂼S2��(� =��=-<�R`=,��;jļ�Ug��d=a�F�_�=� 6�s�5��Ti�%=ـR<��m=��)�1,s���л�iW�`Z!��0�1��<�-��+t<�����5��4s`=����΃:y@v����ךb=����(=�a;����A=�H�w�<��_����<q�<t��f��W�p5W<W�=�=�Lh:�_��<��,=@���3��<X��<t�\���<���@7�<��м �g=ef=��<v˥<�(==�;��k�=��Ti?��a'<â@�oq�<��;HB��xK��'�<�Q�:>]�N<�<��<��=�Ѽ�y=9�?=F�,��x��0��� =h��K�6�(t3��I��'��=6P`��>��s:͏��A�;�R9< �6<���<y�R���u�s���Q=:be:�PM�[�K�w�0�8���O=k�1������9=y�����.=��-�*�����;�.<��=]��f�=�>{<�yo=<5C<�E<0'=�??�<4=$-����=���<�Pz<d�*�y�:p��!�\<J,==�ݻ}�Լ��;��=�ĳ<��������<x2[�*���ጔ���ɼڑH��=��=:{ �L{+�fJݻ�K<jJ�;?�=����}n��qH��G=���o��<$G����<���:�п:�𼼔���:�;�2�Af==,s�r�M=Mټ�ݦ<�q�/5Y=���;')�9�=�l��F�<WDb��l=�[?=8��<
k�@��<�<z=�n��?m����:�k��Vu�<6FA���k=:PK�������l=<bxh�:��<��m<��i��
�:��ּ��c�`��f$=�`��74��Ǹ�3�}=(�O=G�=��b<���1L=����<ʤi=>��<�F1=�p<]��<n��<�m@=�<�"�SI��#M<g�;]P =N�x<��i=q�`����Yy=���<@D�n�= Qp=�g��)�;?����� ��A3<��=��=z��r�<2�4=����d�<xB=:]<I==�ׇ<�q=�%�:�}:�ہ�q��<d�a;cQ��8k���g�=CK ���
�l���+�F<%�Y����<�D�<�v�<>�j��4w=���8=�t=V=<(�=�B�
��<��ļ�H==�[~;�����C�P��%�M=G=�,�<�S��!;����ƝV���C��'���s/�n�����:/��<����Z����4�aw�<��<�U��=	�.��a]�����4<�=
��Z弳c:���$��Y=�g��Aἆ��<a=�$�p�<��h�;�j=
��7�<^�\=h��l̺�h-=#:�<�M����EԴ�ک�����<z�L���<���;�#^��=�P=��W=��Y���<I�=o���4i�<%�<��<�S�<�u�;'�)�eV:=6ĳ<�����n-=�WS=��'�����9���}�4����}c=M9��w=.R��B`����<�8���&=GTL�!f���z=�����;_�@�`v6���@=�Լm�*�倀=�[j���BT=�Gr=�O���,=���z9���?<2�4�E�ټZ
0��R�<f
K<�܄<g�]=���<��<���;��ּS�T��x=�żwS�<�7=�w��!<=/�F<�=pz��Cψ���=�9`=5����?�x%<�`꼄�<��7�Y��<a �����Y=N}��ZR|<���<bJ=�iI= =~b<s{U��d<u�1=#��)eH�����&��;Iю=ܳ
��'%��y7<Df���F1<Ob��=yD�	�k���<���R���<�)6=��ϼ)d�<�t=���<���N|(=/l^=׌=���<�wG��k�<�[��_8<4Ǽ�9��<<���fW={{�:��H�p!ȼZB�KI=���<i@A<�:��u���Y����d"<]O<�>g=3~a��ݸ�c>=�}C�/�л�~I�{2�"Z�<Wl�<��c��R=�O�<�6໾)c=�Ê�fϑ���7�J��<�)&=��<j�����<�j���0�l�:�*\G���F=��W�]	=��j=���nH<�V"���6��=&�K��:=����梕<������ռ&2w�����	*���4���4=�/�=��p����������E=W?���$=&t���>B=0\K=Lڂ;�t輅ʊ����@ɼ<7<���6?��q*=
}�<%s=�S9���=�hl<L�;v��<C�[���<��f=��=�A�<�eZ����\<�>��<�%���<��;�f!����e��;[J����� ��A�7;�U���S�=�i��a�l=O@Q=%*�<$�
<��=a�j<��<��߫��ĸ���>B=��'<F�%�R}�<v<���;���;�<��=,�=e����E=]���q9��l=e�Q�?:
=���;7뱼�NL��H�!f"�i<#��;�b9<U
�;��=A<̼�¼�f?��8;+�<5� ���ļ]���KA<��<�j=}�5=@��<p�Q�uO��V=�;=U)��R�;U�<g\T<ޕ=���Q�(�{�
�ϻ̵����=��?�`�;��G�3����<`E����;<�9�����=s�	=_><��<A�<�3��&=z���g�I��! ��$�a�(��$�2z�<&ܸ������0��6��Rr=��S!=*�=9{�;�x�<�?�<F�f=��/�D�<��'����g��L�<�T(=x����=WS(��E3�F}λ�S����<�4�i���
�0����(��,*ʼ'`����A=}�9=��s<j-�:�z;I���7k� l�;�e�;�E��n�]�<L�ټ�q;���<6+��au=
�/=�NX�0�#������MN�m�N�h	$�4	���2���r�7z9��=�;h=8�`;� =�-��\!�� �<*<i��k���K[�S�=�V��W/7��=�D�<�6x<��u�q��v�9�<N=r8�:���<�%�<��=��<�3=��|��0��b8����n�Mn:����<g��<�;=ڟR=kQ=ߋ�;|�4�+��-���R�%����\��c��=�|%={�@<�1=��e<�v<�U�&oq=�,=�ȇ;1��<��<;g&�:��<�~�<�\M<�I�<��y;{A��'W=�J��KJF=��<�1�'�E��L���i�0u?=��y�g�w<�8��h�r�\���M=� '�ml��`�@�,] ������m�z��9�(Z=��R=*�,�y<�פ<'���iʄ�K�=���<a�R=�&Q=��3��������;o�D=�*�<<~���+=�/Z=�D��O�1�Sk�<�=;<z���_������L��=�Q��Hn�~�c��_ɼw�޼u����K�L=���=ϟK���D<���ł�0�9��<={�&�O�<�S�<�C;C��1j�3�Y��Fm�6�����w��J-=���<c��sG����Z�=<Ō=����J�}JE=�PO���<��4��=M�i��<N��!sx=@�Լ4��<"o#���<�k?��C =����?������[���R��*hR=�+�<V�e=�4|<�M7=��{����<u�<=(���!�=��v�*�e?u����< =�5N<{}3��;<&4P=���<�V=�L�<�/�;72t���T��K�M�:=��<�d�<��t=�
�<��>=>�߼��9�"=q�3=�dy=���<��<0��W�<�R�<>^;��������ӽ1=�|v���!�}���?R=((=8JK�2��)�$=d�V=��S;w��mf=�n�<�%=`�0��<�ļ�]f=�5F���'�E�j� ;�΁��w��#2����ǼZ�<��m;�rk=�ڡ;_�=q��;�<=!bT=9@"<It�<�2y<3�;�Iv��@�<���T�x<p�1=-	<i���`=�G�� >���u�<_V�<���8���E"<��c= +����<j�'<ɈN=s�޼Z< =����.��o���;=<����}<rJ	�̒/��_[�]%�(�<�3H��pY=�=>�3�_��h�?{�{J���ü8a���s=p���)=)ٕ<,�=��<��=9���$���.�@�="���j=?O�;M��!�:v9� ۃ=4�<=$9�<��1=&�<��<?�����;N�;z�3�����G��9(Q�]8�h>�6�j<�v=,�;��1�{ ��==PK$=	C=�=L�����=�b=lL��AP=��N�8Ğ<��0=hޛ=�P���H�=C���봎;�}��7�H'8�B�<�� ���<�QJ<�y<MZ���f='=09={�k����%;TGB�bg(����<�̻�h:��=�ߓ��t�<U@�=��I<�=���<Z^'<�َ��<+�<ʫ]��kI������_�~�l���.=&[<46��S<���<�\=�l:	� ='b�<,?=�
=� ��6�R�ƤO��D/=q�:�F��u�'=u6D����<ac��<�4��sx<��?�,�=]Z-<�G�*���[�<)(=��9=�Tx��2=��=S"=���V��;kH`=�nk=r����9H%@��3�"�W=%_�;�e<�@1<`wS���λ@��<�{�<�~U=�,!='��e��ފ;d�	��:�,<�݃���H<�6*=���r]<�!�Cx�GE�g��o��.?N=��:="`�:n��N����6��3=���;޺;�sּ��y�����Fa�����l�<b�==����:�e����<J�X<~-�<��q���==2�2=��<�ü^�<��<��<+#M=�O����<�S-��zG=�b���<9 	�J�1�x_�<�g��uļu��<��"�)<�zF�0c':���<�i�)�i=z
]=#� �E�;�A��G(]=�@Ӽ��]���S��$
�r�����|�q�B��q�<��<q~�����
��YU=����Y<�K�����;�u�=��h�7>=8=��,�����b��9�;��ȼ?�<��s@�w��;��=$�<M�=<գ�<3��<�z<.a����1o=�����|0�s�D�.��\6�;��B���X��#l�\/���j�<�N��~�=�E(��c\�O=�����:0<|Ԫ���3�e��;3��<�~,=��ջf�Q<�S<�3=��:��2=���q��E�
�<Uu;�7=�����9����2=���-N=�V�K2��Ȉ��"M=@�_�.�5�D��<X��9I=��~�*��D=�X;X���7���J��q����=`�P�A��;�o�<�Q��$w�����*	��"=H�ּ�K?<��.=�p<�_=-��<��<�t��cr=DL=/�=Qv�<�~<�H��j$��Pw��E1�T/J�m9��S��̚?=�OJ=��:�{k��=V��h��<��9�4�=<�<4:7q���=�u�J��<+X��~�"���5=܎=	�o=��Z=|k.�#߷�d��$C</�V=2�N�a��<"%���Q�;��<y?<���<҃��^rX=ޡ=]8ǼoC=�ͼ��&��"b���+�N=�\=�� ��S(���L���4�������]S='�=K%<ډ��|i<�?�:6���GȻ��n�u=�)����ǻ��5�c}�<v)���^�<��*<�&�9ϣ=p$�#�Ƽ%!=�=(f����<�,G�V�)�}��������<�̭:�7��n�<��/<�g=���z���E=�����==oB�������x�p�<�t���_"�y��<�JR<���1��S�/<J!=��<�I;���a='iY�6��;>�@��5�(��=
�E�$<'���}P=	���<^�=�1J=`Ӏ�P�m=<����I�p�p=I�7=䔼<������j+y<.�B=�Q�<��λJڼ<��"=~�"=d�G=AD�0p&��V��1=z��;ư�;��e=�t|=��B��a��o"E=QS3��,���/2�����B�a�J���A=��<*=�~<�ꧻ��`<�:@<��ug;�(=�~���˼�֕���r=�׻]��4�ϼ��j��wt�J�]=$��<Xw=X&���x<��ݼ��<�@X���ʼy��;Ҵ=͏=BW��Q��6��G�4�k=��z���<��=0�5��l��6X=RW=/�=?�<�_�t!���=��*�RAD=)�t�������kQ�<�i7���<�#=�mb�M�1�R�"=�a59 y�c"�:���<4�-�d�<�= ���=k�<
�i��^�<!^3��j=�R��4��;8�=�L�<;2V��-k;�����<�Ql=U[!��+I<�/��� �<eu�=�<��M�U�;�;�^����;4ȟ<s˼�Q ;v�,�	C<�$=ΖԼ�4;��(ݼ���,*�<x��_H�<�lB��о�^5�4�Z�c=���1��q�=�qE=�pd<1F�<ܨ��&=lw'�R�ڼf?<��I���ټ�8���R��[��<Ȧ��%�C=�U��{~(��NE<��<g\����7��cͻ� ���"�`�:=)�6:`�<�5"<�ݮ<�B*=���<�e��(�j���y�,7>=G�O�o�b=Ygռ���)��<�)μߐP�X����V�e�6��N�뼈D�<�P=��<��r��<�fͼ�-��:)[�m
@=�4�<P��<-n-=w��@;��A=��u<�!=Js7�ۚ���܍<�b��?J�~�<*�޼3n=�&�<E�J��X�<�"{�%=n޼�\��K=����='���m9�ت<�yX=7g�;X2{=C\=<W=S����=�!=O��=ӻ[�LH/�(7���:uZ<�k�<n�ܼ��N��v7��G=G&ƺl�&<A���3u,��Y1�J�;�{����ɇ<�=ip�<1(��j�B��<��8;�+=���8N�=C�L<��Ѽ�� =NN��M��뺖u�<��"���A=�=��<%��<��<N��-F��&oM��82=x�;��E�a,�����:R=�o�;LFm��M�:.V=J��<@S�e룻�(%�Y�e�����=bü���\/a=\Q�:��L=�6�<�7@=;:���t�г���:b�B���Y-=,R<m�Ѽ�5��p����<�bM<�eS;�w=�&X��6��(;�>����Q<*�R=FC=�4<N�\=g���%=��g=����Ҽ�솼n�&<|T=�<�r-��~��Sg����<Q=�һ��G=`"j=�%�mL3�Y{�<��$�Y��D�<Ⱥ����=�G��Լ�Bf=C�W=�U{��(Y�tuP=x�!�I&/=���(� =}?J<��%=/�!��ߚ��M'<s�h=	�W=��<�僽Ԉ�v�U�+E���R��6��b�:U�w����<�N=��<����*�;у�<I�"�����o��<��=e��<�yK=�XE<�UɼV[���/�Tf�#zR�@��K_��a=�G<=s��<����N���{�˼/m����Y��Dh�J��:ZA)�y��1�<($_�K�Q=�!F��N�<��N��̐�7&��<��<���<�o=�<5��*����E���&=�=��a��N�r�� �:s�<�	����K<mȻ~�G�_�=���Tg��
��:�-><#М<�Ҟ<ݭ>=�
��{=���<���~�e���Ӽ^���>�/��<n<#�8>=w����;��<pF �	m
=�wU=9w�<{
�A�=#z�<`#�����d_�mKh;ɲo���f<��=PPR=Y�!=�=R:��D;<�P���=�9�/S:��D=Cʶ<�c�<�L=�OL��(y=�^C�F�Q���켏�̼�'2�K:�=$��<�$N=�չ<�d�<̳H��I�<�͇��X�_�=̀�<�'�;�������RF���.=��9�c��3��)��;��t<���;iX.=�fn��u5;r�t����<Y�T�?F�<����ӻQ�Y<��m��ռ���>8���
/=_�<2�B='EV��<�ù;&�<���B,�����9�Ѽ!ȸ;7f�}��;�k
=�ɥ;(�=�I=B�%=s���u��XU=Σ`�V�,=����N��<'�T=oᮺ0e{��/Z���T=s]���ٻyW�}Dμr<�<�>%=�7@=ÙB�f <<�'O=�����+�<��޼|&=y͕�,�2=�G��:O����<��=���#�6<�����r-���T��˵:���<\�m�f���D=�b�<�<���v(=ZX/��<�6Y=ӫr<N�=�����=q��=�e�;��={�K�Q���K�<XlT:0^�=���� ����s��,6�jm68LU���B<��#���:=�=�X�<"���Ҽ��=��]���}*1=\�g=?2= �K�d��I:[�Ov^==��;��<V�>=Wtm����<�T���:�1��ߔ���ʼtӷ<ܶ<;%�<�B/=;E��x��J�<ಽ�^��TG0�XV�M�:���;>�(��U2���&=�mD=�%$=��򼡚��suD=�3A�T*�<@Ԍ���<JU:P⭼5��.�<�=m�n�?s�<�'?=p�J� 6,�ƭE���z=A"��7�=���<⛹<�{=/L�<��T�}��<@$�4��<�4=c��b];@�$���4:�Iļ�1d=m�
=�}�;�9=���: ��<��;<_�<�����ַ<�ɜ�P�$�;�9�V;�A/�p{?=���<1�>=���<֝S=1�=5I;K��<�"(����]�����F�6=,X�<��6��@%�S���G��
P=�L<�a2=DE<�"<빌���b=�'�9^� *E=��s<�.��dā���8=)Ҽ4
�<�NY�W�%=��Z<�7�&�V�r���ڕ����<駧��μ�d*=tN=�f��jmq�YZt=J,�Br�b��;�.���^��T���d=�!L���j���:<�p�{�5��Yr��� =��]��Ν<3,��t�����<��<��I=��;㊦<�3o<pR��7��E�;ꕐ<gл�w3<X͌�xIV�?4,�{�λ��R�V�	=P���c�<���u��;�E�;�fi=	�G=?K<�2=���Ec��z���_<]�D<1�=>P\=p��P=6�<�u�L�_����	��;�{+�}F=ר/���&=W�C�6S�`{_����{켲>�04��6-W�^�P��N]=ެ�9pλ�܅<n䃼?7,=�p���cP=��<gu;E�<<���b�N���7<��?<���;Y�;8�,��tT� kҼ�\c=��Llһ�9l=��y=}o�:�š<j�g=7{&<�=(�N�2�Q4M�9')=���H{ �������Sn��x��a�_<�nN=���<0v<���h��N3��O�<���5[�J�<4�j������<Y�<^��<����N�2=��3�J�8�*i���� ������{=/�J��BF<�Mͻ��������5sV=�#s:3y6=���@�;�%<R�3=�J��Uh_=/��w������<��T<ܜ��qN<���Ii�+�O�(P¼�u��td?=���U�$��D=��@=�V��= ���~V=�v.�ݬ=Ā2�x ��F�;< ����;TM;;9��[�J:�3�<���J��;�	�<+�	���ͼ���F��<�
�&�a=�<��<��:�C��Dz<��V=1�i=<=?(��D=~Pm<�L=S+=��'��E����L��x+=w�H:�G�E==#=3�˼��?@�<}��?�z�=h�<�L�<�5==6�<,w<SIּ��<E�-=��m�a���7�;�C�f�T���<=��C<@R<�M<�↼��{��=��X=dAu�*]�;]�M=�M,�U��;�͕�6�$��y�1ct=��5=p�3<\�W�5M�<����&㼯�����<)��<ڝ�<y����;p�=GY<���:��E����h=�
=���:� �D|o��?�<Y�E=���5��<I	�<���8�tQݼ�&=X�@����i<|L`���7=.�|��,"=��;	O)=(���͂�D���;�sB�D�v����<)�<Fu��U�==?�2�3=���<��@�'n�p[G<��^<e�P��?1<N6\�Z��<�F��'ܼ��S�x���aϔ�@-=�Z=+/=����"F���s=�	�.=������)�?��m=V��<6�L�]�_1�<s)�"�U�/��<�c#�!=�<�@;=j�<��;ͼ	����<7�j�]b=��9i�-�<$�[=پ���t<�bܼf�u���V	�<���|1�`c=_�� ��t|B�*CT��g	�uZ=^v�����m�;>]���Ob=LK=&f<�$���Z��}�3=m�?�E��<h���B=���PX꼣���s�:=�m��_=��'�&<�ͥ;� ='>��;���P=�zx<���<45q����.�N=>H�;�-�<t�<���#='����w�=��;W|=��n���U=e8 =��,<�̻<�τ�%@F=�<�W�<�P��8��<�oa�_U��Ǜ�J����e=O�
���g��{������0<G���p�*ݼ򺓼=�.���bT<a��~RR���i��?�e��<��ݼ;��;
�?=��w<�v=�BZ=>һt<�=M�<��޼�C��!�;��=��=p�:=���;�A�<�7`��hx=��8=D��<P�?;"�ӻ��=OT=�%2��=T��<�p5�X%�u���,������<)kؼ�G
=��y����;z�1=�K<¼:ݖ,��i�	�:�mƺh!����8X�<�K=WH�<��S=�펼�ˁ�7x�3�z��$=4i%<[PF<+��: �˼�1=�μ��w�+�1�A��<06꼓Bۼ64�����:Ord<I�<D =����U��q�H=A~ʻM��<_n
��M=6�p:��ۼ}޻�o��<=Am =�0�<P]7��6=>�t���*��4�<��<1�u�6���=�͛;�����{t����,Q�< �<�(�,�ἉNr��^�;��O=˕\=�}h=�#/�������<-k=����\�<���;��n=��(�L<�,=�Ђ���Y��1$��B�Vp�<�qU=��:=��Y=毆=��<�#;ן2<0��<߈�<�G+�� ��&G���;<_(�<���;��%<�gs=�4h�ޗq�ށ�<Eh=N1��<=�h���ۼ�j<fG�<?�,�rɡ<��<���=u�I=�u9	_=���<����X��<�^�<19i�����*.<�� �Z�����˭Z=����=d�V���g��̼e�-�n�1�Xj �޸I���b���(�ϋ�<���<��v���;������'=�޼$Zj=��<W�]����;H-�<�e�:���<� O�0�=0�k=���<��<�T�<�8e��b@�'��!%��-m=�@�'������Oy=�Zw��P�=��N�Z�L���_��N�<�'�d�`���;�U)���!�	�;�%�<)żD���̖�5���h��R��<=|/�m-�!���<��H=�fѻ��S������.�!"�1��%�<@�9���C<���%���W��*(��ە�<	E0=i�0=�Ǹ;���;u<X�q=��M��f��μE�Q=���}�<RO���C<9 0<@�&�o���U\=*�=�P4��H�<�a=!h<;�;��(����3�(���]��%�<P
==�		� 'J=0	=jM��pg =�-"=ɮB�|M=0="D�<y|��+OQ�A$<�/U=ӛX=����-<K�B����=E ��(�<Qv�vu����_<�	�<��X��	ɼ�/=Yߏ<�m���s���'��MC=��:�Ҹ< �`�<d�*=��C�,r-=œF<�b,��H?=�.�	"V=�=6am<	�u=\���K@=��μ��;F� < y�<m�G��in=gھ��^�=�����<B6|=Lk��+��T%&=1�<y��<pd����FO=|�����������\Q�����������̼_ˏ�?�<��ڼp�o=X��<�x=����{|S<Л��f��X!=��=�4K�AuE�<��TQ�oO5�NGg=�ld=�[���=�[�����j�<j>�J���6�<1�J<=�g��%=gR����4=-��<�,�<�f2=�ʺJ�=\f*<��\=��}=�?�3<l"5<Q���cd��*>�RW�<xaT�(�<P�_={�<W8��m�R����<�<6=�xU�O������P;t��&�<!�=�}�<,�r��<���;k��<+����`=��<��5��<<{Q�����@xO��Nļ[5{<]Jd�!Ӟ<Ɉz:����I� �n<�=T�*��wټ���<�G�>wu���\�� ^�L� =��<�����}<��.<�@'=H&X=�T8=�]�<��K=�C3=oE������c���(=w���q��<�c<K퐽@�d����;5�
=�6�<"ND=�x��U�<���-/"=�I�k����}M=O� =c�<����<;)�<���Pd4=:� ��{�	J�<�я<�<M�J����9�;=�E�0�M�ud�<V��=�X=n/M�+BC��E&=NtQ;��r<�O<��=~�<P= ��"���8^���R��zm��lɼW����;b =�P7<z�d;���<�������p�<�ȵ�$��<+�%�������Kڗ��l��RV<�^=�7�<����
n<���1KX��:���M\�q=��:��H;��<!Y<=ʓ��<��������e�� 0�&2	=�v?��A<���<�#�����;�Ҩ<%E�=�)D=�L���h=�Pû:y�<�!���,��$_���=F
�;�9=H�j�]#�q� �=���e����9Ժ�/;�9=��<}%�;�"=,�2��ּg�:<�1=�2=� O����<u5X;�=!_&=�i~=�1���k�G�����<���<)l=A/n=���JǼ5ai��b?;1�^��wȸ����Q�t��9r�n;�*=x�o=
^�:Z�?�_�=��T�K��๦ż@�Bg=�y��<��P�޲�<��<`�X=ӆ�<����[=5��<��A=��<Bq�;<!=�v2=[�*M��U���6z=n�s<>,��"�<��p��Mc���Z$��c@9@A�ȑ;}9=t(O���;�h��~z�/�z�aQ ��0@�Ԁ='|i<_�>�㼎
��'�c�NxƼ�R2:����~�<Otv<�>)=q$���;���<�]&=x.�� �<�1=jWm��F=?G=��K=*�T<t���ɻ��
=:v]�2gF��X��>�Z�� �|��<�B�<�y2���H=�u =֓q���=-]]<�; =��D����<iW�;�}ͻ�C=�&X=�E�	���c�<�)C���#�x�E=��E=$c=�j=�e=<h�5;P�K�� 2��[<qc>=��_=^�!=�Ļ��<	�̻�u�aZ�<`w���=#&�T��S�}<�Ρ<��Z���k�Z�,��E ���޼��=�=q�G=|[=>N�;QV�;D?y=Z�ǻ}
��1�Z�2=�m���(�=�5=��^=�����<aF_<S�b��P�<�
!<��V=9C;t��<h��<@�^�
��i�L��u��W�:�8<�����<���<�C>�x��5`9�8-=i5��؀=6b=٨�<�����J�<�$`��Q��-=9d)��;��� �#��z3q<:�=x�J���$=sF=E^���
��=�<��r=e!Z�<��% ��j�<��P��6=�ᕻ��8<A?�4����U=J�P�-���	=N���a�ռݼݍ�;
�ۼ�=/� �������;VǼh�=�<J=	�<��+=�V�<SN_=�6h�y�"=��<i�W���Ǽ�Z�<��+<�W�<��f=]`�W;�R4�J�=��G��b=�(=d_�sT'��]1=jD�<G��-�_;8�C��
g�3�ƻ�/=J�n<��<H!a<�]1=C���fA=Y~��;#��&�<�'�<���;�.����<_�<f�C=F��'&�6+���}z< ̎��p`��r����}�=�<U�=?�=��"��0a� ���n�A=.����<J�ڼSHA��x����f=@ڛ;�P=���k������J=ZU+�@y_=�6K<i�=�J���Ʊ�l���e=�Ac=�'��^�'=?=.��<������M=��H�<<�<t��:@B����<�0<v26<#����=��;b��<V�������</|�Q��\=|c�;����<��^��;-�w��G�<ܾ�<݋���p�˻�jX�<{�4=��d��"ͺ���<RA�<e�����=3�<��=�58<E��v���乼1��~��<��,��"�܊��[ 1=��,:���)s�<fI̼��==�꫼��<޻-�̆<W=��T3�=�k�#9��m�Ì`;��M��qG=_�Q=S�18F��<�H<?l��:�<l����l<�}+����<>}��J
I<�v.���9<��=�&����
=ZS��<g2��:�<���;���c����1(�
@x<v��9���<��<��<Db����<M�W;Xȋ;�E�G=�9�<��<
�=vj�n�;����9�<ۍ���Q=U��;J�E攼��.�#�<�A�`�����<�y�t��<�!�ܔ2�[�;�t%��o	�/E��o���1=��]=���<3¼��==�%m���2�54ȼ�IǼ��+=��F���<��<�^���%M�؇;��0=9�={b��bW��-<Y�S�\U����;ʝv��=��<=#��:=^���<'�
=1"��>5=|X1��sE��ڻ<�����];��]�?P��b�<�D=�F=ԋZ=��{;�Z=�<�x򼚤�^�;<NU;==�l�B C:��<���<�~��Ѽ��3=,�d<��<�2ͼ��P�0);��<'Uw�u��==�2=j뿻�At�J7�=�	)�n�-���;�b���y=�� �y8n^�;��<-�]�4/��fi=�UG=��k�����L�<P,"��n.=�-�<��;f��g����_�;7�R�j4-��oݼgh<�KO=z^���伟�9�N��d�K=�.(<z�7���=H�h:��K�!3O<�(�R�y<\��<��ʼ�8缱d�<Z�=�q�<}b$<R�;[E������:º*|)��Y�_�n=��<mM1��	�KY<E��<�(=5��;�Ġ��a-<�Bi�ߦI���4=:����I���پ:z,�<����r�<�b�C=��+�=�zbq�F��<�E���b8=4cW�P��<�Oļ����&i <�[=1)�o�==j�9���<=��<��<?\��Rc��@��z=Qp=�2S=��-�)�����=;�J������쀻@zK���<�X���Ϳ<����1�޼I[<LD0=�����AE=V�J;�ax==�Q=��|�]�s=�>=jе��F༿��l���=�x���5U=�/=�;K���@X��=`FӼat�<���<D��;��<?C<�_�<G1O=)�I���������1�@V=W��<P�д����/<�Ӽ�4:=��<�#����<����h9��.)=fO(=�@ ��`��N/=�[���<zkx<��)����<�S=d�=���<7'�?W��;9=�䅼K`=s^<g�1<9f\<�6�<�����<�n�<�	&<f഼�<=�w=R�J<u���g�%��)�4���E=���� <rS���Ѽ
Q���Z=F�>��{���H={2�9�:��'6=Md��A"=PIr������.=�C4�WB;9�<Y�0=�����=otP�kd���K�p޻��7��c;C���^������=.�z<52�<�KC��/�<�O�<��P�ZX���h��͇v<8/�<�m���W���Gέ�#�o�����7];ph��8�e�m�\=�X=^n}�8����ʼH=x��Z={�9�1M�Q�e�S�м	R=4zp=�9λ(K2�0c*���V<�/t���>���V;��;W����ؗ�X{ż�Q=W�<��<aSZ�T�<�q��`c='�7�ao+��7�<5����0�<����J�@m�;�1�< X�<W=-=���<6E�<�aO�I�U=60����<�U����<�� �<=E�9�/ϼ�m	<Ne=��Y�n��<��='��<bv�M�r=������=��;��ռq��<��<�;�y�g<�h�ӝX=��<�j=�=O����"��>Z���#=5��<z1�<�Fz=�@s�t ɼ���`��nj�<z�}��� =�p��q��<PdY=�=,*6=��!=�G,=UFL=�kp�3��<�H�rI�h�=ɳ=�n�;����D%�Q���8\=��<ռsV6=�e��D缩e�<n���R��H�����<�$=P�=��=��;X�+����s��<FO=�;�<��;=И���A=$?=i�ڼ�t=ʱZ;���'�x����d��T���^5�~#�^���<,�1(w=s؈�j0)=��<�J=�3=]����N>=�pϼ���<��<`H(��!:����*/��*=NrW�"ڼ�L�|�T=\�'=S���΂��N�	J=[3�<!i���G�<n�B<�8<�U=#=�<"#��`{=ӄF={V=}�h$<�5O;�r=��I<��9=B=��<0�����9��a鼌�I=�I���<t�0�"<��4:�����9���f��qּ�I\=G_ϼ��Ti���<��B���:<�C��
�;�S=�ݽ�Q�<0.X<]b���6���o��]ٔ;�+=X�<�����:yň���<?8�<�N�s�ܼ��=���<��P�"c
�$q�<B��B��a�<4�[<?Q�<���<ӊ���Y[�qN=�O��	����K���μ3�5�c찼�]<��	=�j"=�w#���=��3�@L�+0g�K��<��H��9�=e�U��=��=b<~��'<A=7��;�ٶ<��<`Ц<�缻&~=iu�9�8r�6��F�=zR=�\<��.=��=�O]��	�<xGW=�7K=>��<��K���<�%��k�a<k@	={f��Pie��W'<+��>w7=��;fT���Y ���T���0;Y(�;m�<��l=V�6�����_=��4<:�ѻ��Z����=S'��
���<�M�<9d=�J�ꕈ�������g�<R1���<:=jb���H2�gʢ8���m������S�J�'���=B;b�>��"�����6Yc:ȂP��Q���x����0<�a�+��"ڑ<��=����`=� =�ܼ��k=c1��^U�;\rh=ze.=��x��6���ۼ}*:��^%<	�H�^j�<f_�;��#��^�<�t�<�W�#1˻�Ee<��c=�Ow���;��<1���n�<��ؼ.%=��9=��A�h�%��=)
G��o8=<%Z=�t=�jA�,�I:'�۸Py�;=�W;�u]���aҼw�&<aE=]�P=�<�� =gG?;�:a<���qF=�̻c��;H]�]7�@箼2���ki;'*;:�ܼ�m��(�<^7\�̡<��ڼ������=�~ͼ�;�^���i�=0�f=�a���*��v�<��G��8l��W��;��<;[���x���=�U=����S�6= +�";=�^�ڧ�<gc=8ZR���H��)��g<=KX=4�⼨`�<�BG���켰T~<�m��Q��DsA��$C��#�;�&2;#F�~���Km���-�E��<W&^��<��eM�;H��<}�6�$�"=�2D<�'����:�l�=��fD��G����h�'�Q��S�UL���&��h ��v>��Lɼ��	�r뱼��м_28��E=|X��OQ=Pe�4����<�iT=��;nk
���v�'�<�4<��~;Q���[�N9g�<�y�<�A �R�<�_0=r =�S=py�|v�<:ȼٯ=��u<�=<\P=ӱ�<-��@��<��<��;�u��6����+����c���@��2�
�2�=S��#��W��.�N.n��n(��<�<�o<x^�9M=�<½!=V�4<M>���sni� ��?;e��2�< �F=-:��ln<�`t=�K����R��z!�=(S=��<h�����TL=%d�x/S=�����<������c�s�o�r<+�}�%X�����<��`=�U+=��=��<�<�|>=��+=e(\=�Y�<Z�^��!p=�.A�$
����K=s5�<�<x<Q�;<�.�<ͥ9���C��B���&�D=�֏�����
�=����1���UQ=`Ҭ�7cf=|U,<̍�IB�)�~��/�<W>�<7�A������5T�S�����2���]J��rC=/��"�%=�$�(�;�B��O<�ul5���=I=�8��h<	�<=e���E�z2��������<̺U����n!X�7�b����lA1�$�;<����YP�(&��Vf���bJ=Q$��9��]E�#�=���<E'�<�T���8�m�<�4���5��]�<�[:�7_=�I�\��<�e9v|�;�l*�U;���r.=��<\@�<����==3p<T<�|�<���<$߭<�?�;[j��8�<�<6+M=�5 ��9;���<c	 ;����D�G��Y;lc�<4�B=?c=���;\ļ�����)<7�<��?�<m�<?GJ��-�<D�<���R��16�F�Ҽ��q��<�>J�p�W��μ�e$��.�;��_��]�<���;�|���V=��`=W;�<ځZ;���<��=��:��μ�P9=��I�������Y=��={��G$̼|=<��[��]G�׻�@�=O��<;��<A*S<�>��VG�)V����O=\%���fT='<�電1����>T=/m���9���(:&�9��:�=*�]�5R�;��<9�<f�Y= �
=	�=٫�<'�1�S�W��<[Y=�'E����i�ݻI�<�#�s����輶�}��RԻ{�L�ll����<��B�bX�X�d���;v����`�=8g=��;vb���<g��[�ʼ`������J�aȼ�iD�>΃��U=��ۼ� ��ϋ���g=�`<�gr<��߻��H=��
���)�s9�<����5=e��#�d�K�Q��[�!�lNG=���`;����t�<R8�:
�����[����<�R�D�\����Ѐ����;��K��<m=��m�A��=�AQ���ϻa�*=�`0=��H�Od;h��<��~=*Z=��Ѽ݀�S;'=��x<u��jռ������8=L'��B����=C�j���M��e�0P����<��üc�Ǽ?���漵�_� v8���A���v��%=�7�܅�=Z$6�<�Լ��;��;�	<	��<"e=`E=~f(�b:=w�B�7\���-/=�ٻܞ�}�-��)=)��<���<:O�<SW;<�/�<�ȥ�65��\1������9<�C�<e�<��A=���݂���E�p��<<�K=�};A�'=m3��3K<o�i�-�&=�z�<	�|<�Be<���a�t=��<̓�W���	b�f�D�F^�<hм����к1⣼�D�N�m���K=��"=�^缋�<a\)�xD1�n
��\=�
��.=p�=ɯ<n(<8<|��X�;�8�;��<aA�< ��;2|��Ư<$�_����6���6;��<[׮�q�\��I�&�<}
=ut�4�<+��>����<X~���ۼ��#��-�0��:r�!=G���g�<����(L=(L�<��W<N!I=� 
=u�ǼM�&�;_��Q����h�<�c�q{
� 6=���;u�?=�n"=���ֱJ=��
=��]=�,=0��@�<:�ah���
��,-=��!�Z��8����q��缇@�<�'���d�a=.jg=���2�s3h<��������\_޻�O=� H��?F�85<�cG�o�<�Sj�c>�pL�<|�_w=������4����<�������&5=��Ӽ����n�`�=��<aa
=t��jS=�}=�c�<6��tY��Y���P�F��''��s'<�<qO=��L=�>��/��:pզ�HV0=��R��{=n��;2�<���=c�ټh�
�d��;��3�����D���f=��=�7��|�<�A���=���X=3l���?�����<�V�< ]9�|G=��S��:�=3�d�'�k��< @K=2����5<�i����<����<�m��
��nR�~�<�J=�R=�Vd�m��<���<3SC=�4����(�����=BB<��<ĆO�=jE�j�,�'��� �<��k���6=�R�<��C�J4�<-~�M�P}�s��<�Q�=�E[=D�9����<r{<�!=i2�<�Nv=TnT= Kp=p�1�s0�<�)=pF�J+=��e��o��$��&=���<�Y���"��s$=��N�"T=4�C<X(=�;S^=M��>��:�;źt����?�ƶ@:pč�A����Z=*<J=z������X�6�2T="�O��໒���EX���E<�
=iϙ�����H�w� ��<�>>��μZ�E�	�D=�ka= B)=��=�:�<3�
f�~�S�[�;�^=�o2=j�ϼ�Z��%�r���;�=J�7��?�<���b׻�E	=�qS�yߤ�!� ���T=G�	=��<V�:��O����<��m�̬Q�a���dHR��^�9���\�E=<A�Xn��C=����y-]�9C}�q�<�����;=���<h�=��.=�y��m�-��k7=wJn=��ּ��`�=@�7�_�q<�O4�5�{<,�7�u3e<N�~�{��<=P��P�=F�Y=�3=�9<ټ97=��ua����;������=��f=��8�L!.���;�E��8U=G�+=�������<�`Ƽ�;=���<�G�<�G�U�<�[�<��E��F����̼���d�<=�O���q=��`��3�=B$�h�<C�`i�<g�<����4����5<`)߼^��Q[(=���<�	=u�<�qȷ���=��= �F��}J��a��ɘt��X��'��<�/��J�<�q���2=_�N=R����2;�;��<��Z<9O��Ji=�T�=��:=@�5=�3����5<��N=X�Y�0�=�q<=?<�+�:=Ɠ4=�C'=��żĻP=���R=`Y=����=``�<zmX=_,!�2��;zSP=}�<���;f�m��9�z"�T���R4=r=�]\<��y��h�<l#=�X�����%� ]7=��m;͑�<}��<N��<� =�v��� a=�c�=jf(���ݼįʼ.�<�9E�A�A�=�0�*�
<�����q�k.2�'�I=���<�q=�=�M0�<�d%<a]�:��3��~j=��
����;��s�]/�D���><����Z�4���<=��=��뼵t��v)<���=���<�=�?p=f��fi=���<�C���<c=����B�=�q<p�I=w�=���5�)=&�<�E�)=n��<J��;=sc=���]�9=��-<��ʼ��M<k�4�6o=�{a=�$��z�=�!�:)��x%�<�{=[��;ԅ�:�o��ߎ�<�V=�%����<ٻ;���;�o��C��<��<�(@��ȶ<��/�f8��K_¼x�1="
��A�<k��<D��;� r�%<;�)=��P��{����=y�b�q�]�K-ڼ%��B7v<��&=�_R<��<�<%"=�N�J���VM[�i���J�*=�[f='{=��B=E���C=|q=HƂ<d�b=��N���;V5�<Ko��NO[=���<���;XPռ+K�<�ڌ<��ټ=��;6L�P�=�켯��ܒa=��=�	=*�Y<���(-�<�{ ��1]�H�Ѽ�G;�[�<lE3<��O<�$(=�ʼY��Ɠ�I�L=+����<�=�"/�<���"�=��<m"=s�d�n;cb�`�V=�E���;6~P=]�`���<C><nF/����v�,=T�D<~{1�kZD�a�^=�=�r<�Sz�Mb{=Vs��[�N����)=�2=�~?=1W����:y���x�x���=2�4��!0=�h=ܞ:��T<���<FE;*�=��7����;jw�u�ż��¼��ۼ)��<�����S�< f��T���<T0�<�T��� =;�7��
�;^j��Q'8<,�뼫�6=���#=n��;~��G^�<6dļ�\�`�Z=l�e=u�=�r�'G�<
���]\?�;==�}M<�L<��%=�`<t{�Ÿ=�_���0�<�ו��I�N��<��1=���<'�R���1=��*=��G�ʐ>=1�$=/�c=��,=b���$=Fh-�fG���K�����W<�7,�{A=\)��@�<J1�s��<�ƣ�wG,�[��p�����<=�(]=���
�l'-=����eS�<��<�.=�����I=3HS;H��<I<��H��<�B����	�ƻ|�T=���,=�io�ML�F&�'�gq,����f=Wh¼6}»AP=�=�94=a떹.�<x���-C^����;��O]E�z��<xe����>=�_=�!�<�L|��A�<|���S=F�=��2���B�������A��˼PE<��e��8�<F�ļ��=�ǭ���<�p�Tᄼ+c/=��=�̼��O��k���D��Cz=Nj=�'O�D"�I֜< �:}VT:���;J��<�ռ�ƹ<X��<��2=��2�������d�}�l�<q�o=����S<#^�<#==���f����"g�����x;=�]¼��W�r'ƻ��=�r"������Y<ҟ�k�
=�
<N��q�ּG�G��I�<�t�p�=�5�a�w����;,*��#�����»�"�<��O�-�Q��9��4=</����v�$5=I!<]��z�V<�A=dE�1�h<x{=��<N�#�K�<1{=��<�]	<����<?��*&=	�ༀ2=�=���<rN�����<�6=�oB=�|���>��`�)�%=a��<$K�<ŗ|=�_G�@[�<�=λH70=�?мn�W<��q=��I=f�5={J��<�	=��'�Opʼ;��<�6��=��ü��?=]�]=b�N;Y?м�<�<�n=�vM;�7�~]�s�&=�M&�W��<>�3�w�D=��$�(�59>��p	���O=_�y�0\��7�%�A����*=���<�݃<� <�o:b�ҹ�/�<�*=S�<V�	<��P��<�s�;������Ԅ>���n=:�=���<�y:*\
�΅"��V�<��;I�8=��%=L)üy���o��;�k8�z(�<+g�;�?=�gA��X}=�X�ˢX����1՗<���93 <�ȁ�����_o=����W��	-�.Jj�.|=��b_�:s�7ƀ�?��h�ı�<͉.���\=R��;J$ѼPO���=�2+�Pk��
�=�	��Y'<�+���;#�<
e��W��@˻r(=�W�hk�Xg?���=��N�q��< ��=m0!�G(O;�J`�?���B��=[�o=}��'�C=�*�<h��=[=��0�k?�2$=��a<��	=�����l�w=��<�:����_!�4A=�;��>�Ih��,+μڏ4����C��U�<-�Y=9��<��<����w��ma�� �=�C ��#=q�<~�ռj�=g�K����={������<�A�<W��<��c��m��FL��v�<�^�;r�y=g��<�g�<\8�<d��/=��<�̕<u�h¼V�!�N�=
#f=�Z=��Y=�i�<�9=�eW=t�_=4� ��:����1i=a�����d�"Ժ�W�U�P�.� �np6=�mR�bn����;�	���zw=H��=���.X<��(=�f=��t?�<@~<�;)�<�-4��j�;T"��Q'A��Eü��x5S���@�~4��;�J=�jp���$=Ԧ���ͻ�TV�k����w%=4p���c�Z�5;/�=(�(�in�<L���~d=��=Ӆ�<���X�<�u��b<%1k��7�<��b=���S7H�y%6=v�9�]���+
=��h��N:��6��ü�SjR=��_0==8�;l�;<�$�"ݻL�W�L�b�K͉<��	=����dD<Co��V�s|!<x�=B͊=�sO�B[�<���<!aQ�K��<�ݣ<&�=�d���{b=�[=�%�%���<K�����=� =_�<�����U����;���zb�1X�*�"=�Bb=�
��հ�T��<�w�<��<s�!�>`<ä����M��P/���l<���=��W<9c�<�R��`��~5=-����<��w;ێY<��ͼ��-���5��B�&��<�}a=���;�@��k�c8��@h���c=�e,���;|�j=e�]=��<Z؉�����f�m���ż���<��z<iHN=,\�;��[�/]b�M弌S0�_���Y�S�7~\� �Z=�����G=�(��]��>P<��H��#�<>�8���<���<��\<�������vc;�p=�����˼]�9�G��w=��9=��<9�t��,<���k<��8|�o�=�O:�(;�8�n�I<���85=S��<��L��$L=��_<��p=�W��j"��?M�<x��<Q�W�I��;�w=p�<x;��D��r��#�<�,��iZ�/��eM�<R�9=�H3��E��.<�<�
�<1nH=�[�9���4CK=��̻x����=���f%=���`���
)�Қ�<���;+ְ< �{=�il=��=ظX�=[���\����v�;��=�y��13����<Y$y��<,�Լ�ֈ=pʯ;�����:� ���;��<w�=h$�<a,����6=gj��Lm�<�;S=�����@�V�J�9\V=l�N�D[J�R�=\+�<l�=of���m<n�[=	g����<���壼i�f*l�N�=��N=/��<t�$=w|z=�_r��⳺2<�}�<ϻ���[亊�ɼ�!����<Y=@]=��b�a�2��.ʼw�!=����a�a^g<Yü��+� &A='m���g�����=�1#��%���E�E3�����N��;�w��#��K���s�<�G�M�<�uw=�$�;HQ�:�U��"�a=�J���;��<����wc�]=a"=T�;��}"��%!��囼Ͷ�<1�k��.�bf~<�蟽���;�-^���<6/����W,[�y���$1�<���<
%!=�#=�;���4��;U�P<Δ,���
��++=��/=���E�$����;}�<м���u�:�=�g=�"�<u�m�U�<�+�X輬u����>��ˬ��N[��_O=�d��f��E�?�Uْ���9<},��6Mʼ¿ؼ�3q�-{=s��7O
=A�C��+&��ͼ�hm=wm)=��<��<�¼�Q�<�<p*<�!$�LH�;�.M=�{�<�K1��U9���Y����
� s=~�S�.����<[s9��i��9�4�����>`�;�P=;�+�0��<��/�`]�<�zt��=��m="��2(!=,�n�ph=��fɻ�c0�Hkv=a�i<�<��׻��;L=�$μ�UQ�(צ�/<�;��e=ޔ�;g�+����.���,�G�����;8��<*���p;�@<=�ɼD���v$="� �j�^�[�<�
=$R;=��i<�{@<!CX��P�<ܺ�iF=NS��<F���,V;]	=�f��}܋��]Q<*�03����� ��o���qy=3�<�!�Ӧ�<���<�Ի�E_�{I�<j#p�1)="�f=	aI=�����=}�N�=�堼��>��8.��H(=x�
<�=4}N=(+l<��q��gd�+�_�Nm�,|�=�=g�i��:��E���=9�f�3=$M =p=�� ���i���:�0���t��Cڻr0��yL��3'�Io<��-y+=$=x�� �;�=2=��>�<=������?e=&�ü��ȺS?~=F};F�̼��}��p4�)^ � �-�$�Q=m��<U�A=��#=��$��ˢ����P���p=��!���<��ļ���XZ=Y�<f=�V�#?[��)=&<^�1��6����<�zB��T���<�8�<E��<5p��<B�xq�<;�a=�x=��<����h�-��<a�?��ȹ�E�"=o"���=��j�)�ټpY=�V
;D+��wﺻ�d����A�s��k�=S�Ҽ��ټ��˼�P=��D=����;�V*=wwH=q
W<=�o��V�<��=/��<��;�W=bY[;� ���Ķ�pl`;Ъ@���!��8<�\=��?=8��;�,=��E�YXL=?(4�݅3=�}G<q��f�K=���^�T����<WۻH�e<��;hDJ;g=׼i<�L=G5=J�=ye�<� �^�������0{��)��ֿJ=��8��.=d�=��:E�s�a��<�tO��78�p�0�*�;;��;��]���,�e�n<�!���5L=�J���O���=�Lܺ	6�_g[<)	�����;Wn�;Ӂ�<�8b��2<}��ټ�u�<�X�{�*�@
��߫ƻtt;�� �Nbw;�x�,��<��������$���;yw�u�!=:e�<�Ҽw_�F�?���<@]�<y��7[�<���rˊ=�ͼ�~�;̓���T�<��Q��*ͼ�����vn� �<�4��_����W��#�T=d�]�;�:��S<8>�<hw_=%��_�=�7����]=�Jb=��C����?�Y�圔< ����;;�>��8�=XV&;oa�%�R=?0�<�n9�	�ڼ	a5=D}4�ӸT���F=���2�/=��!=cB�<��X=� =N���MFi=�P<H1弊�c.ϻY��<�tj<ST��	6*� L�<;�>��$?���ʻ	���$�=[�-�1=:=�6<�y=(̼���<tĂ<����d"�.x�<��~�;3,=J%=�>=�8ܻ�'=ÿ
=�X���<2i.�����<!Iz=6u�<�n�9:r4<����!�<�g<{���Z�<���7o=;ۼ����j���R�;j�����?�~u.�f��:��;<�G��0*��b9��y1���=�a�ڼ?��F�4;�T����<�û<�f�<U��Nm=��u<l���k���3��h�H�Q���_�ɲ+�x�A�,.+��R���:��P=�e;�5�+W1�k�;����<��O�l|C=�:��z�I�L6�;ἃ�W=�⿼��<��\��+P�s�G8-<&���,W�<\���G�^�u��(�����<��b�y=��<��<�ɀ����<� "�'���m��3=�Dp���I=���<����
;=#�=9)�<��9=��?=�=�����}�
=N׼��7=�8^���[<ׯv<,�3��{<!��>���L(��!�<8=��?�
��<�b<ݟ<�I�;�G��en����a,�P��<Չ�<��d�7���N�t�ޖ�<�=O=��}��O���:
=�/@=�u��B��"+=���g�<q�D<K==��̻�S�=Z�=�2�(�A=���k[=���<�#�<�ɼ2�x�Ә4����Ak=�im��h���� r_=�@]�$V_=���ף��7=���;K�̼��L=D�<��Լ)s�<e/����+<�zN��Y
��&ȼ�[�'H=v\��ٻ�Q����<.I=]�&=�a=�r6�0���ok��1_=��
=���:f�<�;��ީ<@�1�Ȋ�,9��/=TNL�U�V�Iw+=��(����<	#=�؄����*��vߊ=��3=#U <
�d=�R�X{��P�+��/3�E5��}�U��_'��]c=� �<M�<_�<:Vܼ.�c��OԼN�v<�d	;q"��r�rɼ22g=_g=4�λ0œ�6�ļ��<:�b�d�D���<�>�<�0;��"=�);�%��[:=Y�<���<'=��q=ҊҼ;7�=��=�=��E<� �.UD�o?�<_�ۻԄ<��;�c39�j��H�;�m.���B=���;�`�<�N�v�P�D�8���d��=*"=󊼼E5B=���eD���B=5�伻e <�sU=Z��;uf=$;�<�I�:�~(�Q^�@_n<���vH}����=�F�<��2;��=2�T��;�M�<h�#��a�<��)���i�Yh�B�F=�{�<|�⻣I�<ȣ���T=5>�<��0�]��=��(�M1=N��<����z�	������2<�;Z==# Z��}=n�1�B�g�=l�<�V�<w�<VaV=t=�w�<m�<ӄ�</��<�.V�#=j�V<����� =�JK=%|]��]�N{���,?�8�Ҽ���<��<�z�;��6��u��O�<�3�b���@�86��%
=<i༰�1�0�o=
A��N�R���-��o+����<�=��<�u,�[/¼�!=�T���d<F�����j=�"=𬺻>9?��o<;V�h�Wؼ�,��8�9ɀ=�Լ�㶻���n.���(;z˾�7�=.k�%h�<lI=�ż&=�!@<��=�D=y���.�:��3=�=[� =.E=tZ#=��5�n	=}�;j�
��ּG9
�a4�v���K;�ꋼx�J=2*-=+̝�X(�<6:(=9�J��y=h���4=��K=
�/=��!7)=x�����<M�<k��;(sQ=�t�<�;��R��֓1�A��<�}���Oc���2<��O(�<�Oo�'�=�j-1;Hi =b�=���;G)$=W�.=(��PMO=���v�ȼE=z��T.=�v�}�=qO5=DW���U�2=���<M=�m��O=�(�����;\�<Z^=R��<�M�}�G�wŻ0P0=��<�᝼�b��v��U��r���_���K=��L=�I=�E:�����Q�u=�5�<��~=+<��2%=�����v=Ec:G=��<��<t �<��i=>o����:{�6��+�<K�ļ�,<u(	�
�`;���;ۿ���-��<=|��<Un=����x��)�Ǽ��-=������S=�1=wQ�����<y���X��.<<D%��K�;��<B-2;I��<W�<��=�Bj�|��<��==�G�<d����N=�6|���s<b�S��C?��_�]�B���<=��4�-�rI��N����8<޻N�{=1y<���<f�=���e
]�|�=;�<��
CI=��;�p,�)�<[�S=��p�qQ���Ѽِ�<�-�=1%l��='����;5<D�=�d=�M ����TN���w~��j�1��<H�"=�9�;$:�(�弗�m������g!=Xz���T<ܼ��s��]/�<�)����<����d$��� ;�@�u�"�r���x[Ǽ󣀽�����|9�4�w��u��9�ڼFy�<����8=Ɇ(�.��<ݹu<
��� �;a��<�1�� �R��Q��2~=G�:�ۆ�<5{j�`�9��"4�?��<8`˺�_<��<�=�D���rF=/s=y�7�Z��<OP�<�^.���;++��H��P"���:��D=|������n�<r��4"==0�;��(����<x�==��T;�]?��N=k��'�λ�(b���<(n�<T�=-�S�<��<;>�TR:=�����J��-E�&!G�X↽�K
��=�Q;ˠz<�B"�;�=}�.=�
=;��I=zڮ���=���<��<��;G@4=�'����4����<:@<F�;�s�����<i|��hjc;Ӳ:=���<��<S�ʼ�If��7:�~�<���ͼɪ�����<?L������U�&��ŕ<����z�<;�1�L�5��o>�s/X�l'��O=�K�;�X�=��x<Ҝ=�"�=^�';s+��h��<������=� =�yW��or<ļ��=�U�j��=;�F='䞻��MG��)�#=�W�;3�<� 5��D��hȼ6%��*<��ļ�m�<�jm<��_=(&�<�U��/!=��h<zX�c�.���=rbP�.ڨ��V(�<Պ<Z
���	�=�<�$���L�G1z��y�b�":O��<*�\<��f�^�(�g��<�G8����}��<Z�_=�DP�u5���~<i7�͑��ZK�=I��<�'���= �x<~6=\.R�Y���༎@�<:G�<��Z�=�=Rl��軼XK<G"9��8��|=�����м��=�F5�]��*E<?Y���F<)��<�"=t����>=سk�<[�����q��"�9�z=ip��Y�A�|<#����L�;8.�<��y���鼗�O��jۻ�۠��=���|���~&=�*���;,�b�ϑ9�I~x=�(*���<O�˼��<@f�%Y2=��<��P��=K�2�y�<l�<��o�8/���A$,�c�X�����p:h���:U)=�{� �<��k�x��
�H=��<�¼)��<��J�A^h���;��3��,=�!.������`���<� U�y����=LP=�D�Z�2�g{
=��ڼMhk=kUs�r�e='���F<����=�D���'=�b%=�h=0����Ā<�[!<��'�ۼq�o=��<��<����T��"�7���+���p��;C�r�s!���Ve�O�<N���$U�!�$��:=Ԭ+<q�һ���<��==��%�_�< k^=ے6=��V=��<��f��L�����<��!���m��{=t1~<�%���Z���׼���<e1����+�ٺ�Ϛ<�ol;��d<��J=�| =[z���X�폕=�x��>=�jn�f۰<��<d@W<g�=,QQ���M<|�2=����e�=����k�#H�l&�<*�N=)����#<�f|=��\<�/=�D5���=��=��>��*�N�D=���2c5=�MO��H2�Ja=��==~j��<o1=T�|���<$+l��
�=d�K=b �;7E=6aż�0C=q?
=H�J=��;��7=�ށ;���"���>�=��4<��n�&�<{��%�`��O�q�m�'S�;	Y��"=~���MT<�����=1��<�=Ƽ�r����=)�ؼ@B�~W+�	N�㩨<|<�;ԣ�R-=HKr���Լ�G��}�(=��(�e��<1�ӸŐ�<~���<CH==#���N=�PA�tZ=�	=ɓ�;P!~<G��;�J򻼿��&1��㛼e4=<��Vj;�#�5=����Ұ�<��q=�]=��?���?��45=pr�<;L����<�$<��e=W�;Y�߼o�)=y�3=��<Aj�<�4="���p�<p�=��<�ŻH!Ҽ��n�(����Լ��=��=$*��x�v��;9�<�Fk�sO��P�<享;y,B=������<���Nu�;�,���:�%����r��'0<PS�;���<�x���8y�^F��A��-<m�_��/ܻ�ܓ��@<x9��;��l=��<=��=��*<�1<�*=4%=�^�<�U�'=�
�<��x�j����á<Ai5�y�w=��켶HI=�ۼ��=K�B=�A=���<��$��_m=e@|���<��/�ʖq<���<aR=��ɼ[dO�S	�8~�'�s֜<j8S=���<Au��ٙ��cV=/]B����=V{��H����	�F�*�).F�&K�;GdA=��2=4E��-T���= <�$ɻL����Q���<܏=��d=�!!�c��6`�H'=%�2=�	ɼ*��<�"=��W=h	ż;7=>Lؼv�<� ���,Q=)<�������3=2�˼bd8��a =��R=�z=շ:=ku�w�;D$4���u<ؔI��a���U��+6<n[���C=���<`��9��)<�>==y��Lڼ<O.<��<��%�;�G*�"J=0.ἵ�㼵 5=0��=�.S��+T��M��B���:���컢q��{�&��i<����z�[���=�ߜ�0G=�ʽ<;���=�X=�{�kh�;I�����$<�/=A"��8�)��;9�!;_Q�<0Ӄ<�(c=��l<��<��üci{<�B=R/ܼ�52�,�����1�&�b=��'<��=�	Z���; !¼HUe=�H���E��vL�	v��|H=7��&��������q��1E��:���ժ��1�o�<PO���A��I��gfJ=�T�<��x<1��<�W�<q٠��_Q=����"�<V� =h�����e=�1��&<���:�8�3x���vm��m=A8$�0{V=gR=\�=3�N=��:<^�;=s�
=Df�<�H~���s��Ց<���<�U=6 �:�^�<*Y�<΃^���Ѽr=�(��N���8=ϫ�<�68���Ǽ��#=��߼L��;̤	��e=��"�������<��/���*<�ռ�0���ٻ;EQ=��<���;Ģ=��ɡ�ڳ�����j
���4���j=�L=��$=i�����'=�m:<���p���V�;������:[������<H�t=�C<$����E�x���;�a
=[�G���>�/]*��69=f�Z=���F��"ޒ<P�L������oS��R5�@5;��=�DQ�>B<⟼<�u�<�t_=@5���Q�ƑS=���&�>�N��X����6=g�ʼ�=��l<z�p�L
�L;/��\��=5�O�j
�<3+4=y��<�=g=���=�e=@���<E��i!�/4��įE<'�<��A�$��x��N�<���<'���Mޥ<�s�<��<�Z�<�<��@<�]�7�cM�<���W�!���<��ٻd�i<c�!=f
)��X=Կ��?�̼��<�<=�%(=�<���;.;@��f=蒖�/�=�D�j�"=<w�<ީ
<��ɼ���<F�_�X����'7�E�
����+�Dj�%6x�o������� ����
�M��{�<&f�����$f����<�]}��Ӱ�{ټ�!�h|����=� <�����Ż�Q;;�V�{R=A)=�Ǽ�7��(�-=a�5�-b=@��<��0�`}w<K��3�P�V͙��>�<��S=�*�<���<Y��<��q=ø=o�D�G{a���D=w�T<�u�<�T���7�����;�6�<�]��H�<)�#�ޚݼ�q=��=U�w��d=L2.<��!�or=&��7�}�82
� �f��:�EC�U
=d�U��7��O�<�:.���g�b��^͵��C�<ּ"�_�;�&���@� �.�-����'�_��<�B<c�d���+���Ǽlp�<7��<����im�����̜�<�p�v<	�:�s�;��<!A?�l�<�=�<�V�<\��<�{ż���s=��Ѽ��n=g�k�틪;	i��O�a�L=S� =�<=>!<Ks=�"^�����P�ȼ���<`��EҼ�sB��q��������=��=�+�;k\H<�Q���0w�`[=�l;�<C@_�7M"='g�<��=~��m,�h<:奻�^��+0/���T�0�
R��@�:�cJ	�ӿ�<p(�<|�{=�b�ZA��%=oIJ=@�c=��E��+1=-�z=6C���{�� =9=M�����<�CN=�~�<=Q���o)ܼ<�=�p�<�?C�_�;N�p;�P�<�ȹ;��U=A���њ�<��l��Q�<�Ƽ��ݼt�@�y������'=���N��<�a
�Xǰ9�_=6SҼR�&�e��"�N�<�;qFż霎�l�a��<�� =�z`=�#����>Q=�ٌ<��W=����q3=(ȡ�9�=i�V������m�!=��=���d"<x�=�i��0�6P=�E=]�w�<��<LH�o�H�n>=p�r=Y&���1�A뉼7�'<L�=��?�57P=j�ѻY�Q��:;����=��6��$<$RH�E6Q=�}�:0�\<����z�<ӓM=�	=ʨn�23�Dأ<w�<��3=�2�<�l�
-����;s��@B��ޓi=��B����<��<ja�<�\'�l�?=GB�f$�uׂ;1n��=���X�C=�����y�u�J:B��*=�#h=��4=kɻ<O�o�Q����I���X� p/=P�>=������*f"���R={P�d��<-2M���d<�aB��'X=� .��Ju�L�`���<����vO�k^�<��M�Z�=H�B<���<b���T3m�f���_���i=����T��~<A�#�v�O�"\= »�=<���ֻ�:*FJ=D�=uÆ��i8�"N=g<M=1�C<X�<2J�ݙ�P��<�˝�dûa�<K�N�?Tb=Q�Q�\[�u/�T1�;-s{����;U�<��<$֟�t�b���A��2<��:<��<Z;��</;&�=cGR=x�2��^<�!���?�>��;�i�<c`�<%f���A��S=9��k2=Q�#)=�2�<��]���<���<��Լo��ȼD<b���X?�N�7�𿅽��F�t�A��%����ҼƟ����x;�16�q�<�a;�4���0=�Od;L�<���[��<\R<ի�������<��ݼ�XY��tD�Y�7=��[=���<Jϼ��ļ߰� P=��j�<j%�<+x�<U���\<�==F"��߼&�F=�z���G��=�"~�>����]�<���<��:��A��<�1X<X=Q�� �c<3?���D��	�:2a+�A6�<�%�<�=��\�<���<��J�=�1^<ϐ��o�=M�3��e��$=)=O�F�{`�<˞e���i=�I <�b.��Y1������l����sD��Q�<�
�{yj=����b�c<5Y�<G �<qq����(=�=M-=�S�g�K���w<�B�4s��c�?0<�����<Gõ� \Ҽa%�<#�<JxZ=E$
=S��<l���	a�<i?O<�2��f=(��<�B�;��o=����"=l�/��zۼ�Z��2I�A��<����x�4��I����=?G���<�Tż����=i����<�����jK<�j�;�;ֻ94Q=~W���	����<z�G�ZP{�Z�==��<�M.=�� ��i"���L�+(�P���#��dKl=o����@=��=��<�m<���6��u=�{<��?���y=�R�(�, ^=ͳ=IB�=y��<i�:<S���JD�x��"5==�h�n��<;�n=.f�7�	����@9=��ټX���?��;�l@=7h<+f��gV�zr�������.��A.=�(��u�i�5�T=�5�<`�<g�}�v[��ʭA������<��f�iY=��_=�S:<�R]<'��x=�7ؼ�-r�zB��N=׽������~8�E�9����<��=�>(���<��=�r�!�4��t���|��:K=Q�M<��9���<}����h;=Loj���ۼ�e=�u<-��;ޘ漠=�G=�� �;�`��<�C�<�r~��F�<�i9=1=w%0�(������<�z�<u��<�q��)�g��f�<�\W����<3qZ=�*=c�=�X�<��=��Z='^�}�췼T=��#=�P=��T�e��<yA�<�{�o��<dZ��Y���F���R=��P��(����J�a��O~="BW�V�_�[C�yٓ<T�]��8�<��G�b�=7�.���?��r>=��T��G=�� � !�<�|�����:�<��M���)�ނ��#�<ņ����ݼ�;�=RL?=���<��=�����[<w"6=�2껊��<f�|<I[&�8!:=0Ҽ3�)��51��Ѽ�~�;�?s�(�=n�]�~2V=�?�<s+J��d�k���i��@k��e�<�Gc=�#�<��&=m�;E��/_���^��S�;T�I;�m�<C�%=W��ퟱ���6�Q��,��.%��2��~�<;�@<I��H4�<�]=��M4�4�����R=|tp=)=�.<�e
�_�=�������L��xE=C3�;�=	;x3���T���:|�<��;9�!=#���`& <)��S=����<=�7=	5�φ.�ʚ�|�F<Wx�<�yN=��G<�V����j=sEJ=�	l�.����:�P<:��'`�� �����~����r��޼�1���ڄ� y���33=�Q�����V.�=Y8:<��	=�n�;8ț��i=���Aؼ���<z�����(=a�a�8����<��y�n���+���)���
�/-�=]U=��\�!���0���=d=J��<7�����<����s�<g�*'����8�(�=ѹ�<*¼V��<�9�;qr =��<�(�<p�#=6����07=�F.<���:/*=����je�i� �P�4�l���$=?���Z�����.�ڼ���mY�<�m+�]�E=��q�q�?�4��<��@=i�<Q�|=�=l��=S�[=f,�<��<�=i�Ƽ>-��r�����E<�<���#7� #k=�=I�&��(�|P\��cGX�l󪻥� =���/�=r]P�6�9�W^��v�3�avw<�������<�Ǽ��5=X��.=�X:=n��<-"��=�R0�\��zf̼Br=�Cʼq�=�	�l���W��7��jhs���=:�j�f?=���J��<�O;(I���G�YAh���e��I'�������@=>G�I����?���r(=�Զ<w�,�1�<L^�<�B�<6� <�\��z>������	<�sW�OE=u�;�2�<�I=����(�<�$���f�<�V<��&���f=؆=�^����m�=�6�*/=��<�L<�D�<�V���X=Yo�<Re =���B�n����<�pټh��<dW>=*'�`�e=�G�<�0[�I;�=�Ԃ=W�*�f	�<��I=�8;��I�qx=��<��=e�`� =��k�iE�LG�8����9<)���<7=�ֵ<KR��[�3=��F=�ۿ��S=�b=:��<�Ml�!�����H�?ㅽ��;ɞ��;%�O6c=�8<W9�;�3�Αp���< �}��Y���8=���<��;=ta"�t>=eA=цV=��R=�s���5���:��<C�r;���ŏ9���Z�=�H9���<�
q=�iƼ����/��ؼ�6-���=�=_�>�#���t<<��d��A�`<G+Q<��>��~��d0�S�M=�c}=�X�<�� ��<9񮼒�ϼ�;�=�* �V�A=�Z'=�ڻa�H���<@��:3b�d�?�hQ�^�μ��B�;��1/<�^��û��C=I+=K�\=��.=y����v���e)���9=�ۼ-�F=
w%<�,�(���]���w3��μ'�=�9�S����G�M���A�����=�O{�Omr�q�K=�#Ѻ-`~<��M��=�==R.;v�
��̤��cż��2�Tf�<$�=�Z�<��=�FK=�"���v��Z3��`��l"=�eD���=@�7=d����'��6�;�h^��{=�m��]d��N�<hR�<P�<��@�o��<�M�<��:��R)�Q'H=��j�^;=�cr�u�[�_�<8GӼ����ͼ����M�8�=^�<,�;�7�E��|9�#�0�2:���_<�x=�=��;�K�u���a�~�<l�#=�}�<z�[=�r�=���<4@6����<kԼ��<��!��T�<��N���"��r:;�����u�$�+�X���Z�]�1=�߼�O޼��^���
�	=}=);^�q��r���T�l�Ű�<�j:=sp��:��U
�<� �<�7T���<фF���)�-�]���=�ּG`q��@;�ǿ<k��D;=��<)<<-��Eg=��Ӽ�!#��Ya�Z�xܜ<qM���=%�P=C���`�;��a���_=3�6�p�c��<�tc��q+�׹�<�G��F�s�d�
�F&&<���=��>={3Y=S�=���<���<��=����3<ۗ�;��<~��:=��9=��<�|=�y9=B�<>��<6u;��3g<�^B=��<e�;<Տ������1=� �d	@=�E�;^���V<bC�:="j�'���m2=��<��7�>.=!gF=��<�c=���%��"�㮲<�=�G�֭/;}D�<J|a�p:R��E=L]��I�<%���e��^��<��;#�$�Ma�����o=��1={B<F�<Y��".=<0�ks��
����*=�\�=ȱQ;�!ͼ�L�<��
==��;i9���=�U�������-ES��S�vK=(��c�:���=:��=z�R<l)����qTH=��P��c=R'=uFw<!�P��&6=����^s�S�;�:=�j�:�~�I!=
D�#J���5�<����_<��*�i�F=z�޼��5���"�_��<G|���=~�=c�[����f3H����;���<a=bּrl4�@I7�PL�;�Ke<�~��o����� �Ř�<�]�<p4ͼh�<���������M�lB=�������=LL��oҼ��n=ȹ�̋m�J�b=��8�"'��
�u�9��9D��1=�5=yC�vX��K=[ػ���<���Vҷ<��p�SX=�Fɻ�=�h:=d=����"s�����E'd���<�08����<�y��`G=���<�2�<�m�<i��<!`�<�r!��Y��Hڼ�t=�,<2�;`�s;�I���;��v�5Xi���=$
L;5��\� �/7<� ��7�w=�UT��H伭*7=�I2=�G<< �<�'�<m\�;��K���<ߚC�?1üK��<�3=�>t�8��6��=�e=~��սԼ�YC��5�<u�:�{ p<'q���g��q<�6,=�S9<�
&<�l�<z��S��<�':=�OE�xpx=���X�y�Ğu=ɡm��W=;��<�g���J=��<g�%=K8��&<=��*=�.S=�G=ª%�iU�<�?d�~m�ѝ�<��<]��<���:�f���&�Ǝ�<7�,��R�<T�<���|q<=�󁻄�Q�s6�Üü�0X�}�9vt���lm1=�J=7I=�C=FC=1X)=V����:<�׹<��2=E|$=̕=���s��<(��w=�.j�H�����NP+����;{��<�g%�����Jr�j�6=�N=^����6<�&A�-����漏�g<�=|��$��u�a<�ܼ
�`=��q��'��(2j��?g��<�<�ܼ�Uɼ)=O=��T�^��<��0�Q��<�Vʻ��D=ۧk��=<4<�ռ��/��x���7�m�S���<;g�<��K�R#�< Ἃ��;fC�<L<=B�W<���<�s=��l;�Z=zbE=f96�ވ|��HI=�%���q���P��˼�����H�~#_�f=�R=V�:N�<=ރ=�6=�+='ȼ�,=Л���9=
�"=��<�eV��^=�.8�	 ��=sM���s�;�|	��^�;��k��5Y=qK�v������<��ʼ�5=wCV=�⼖pE<�db�P���.=�P��N���.�=_��<<������H�<�7=��X���5�K5�;���:���z�<x�%�����A��]�<�i�;�q�<`��I��u0�:=�:�� ؼ����Mo<�Q�=�,;��=k�ּ~@=���G�7=x�;[<T�;P�=�H���.�.�=X�<N��h�=J�<����<&�p���;�B<��o���-=q�=��<����E=%xS��s=�T�;�?S;�����<\������<�7<Z�>=̶E=�2�h��;#=#��<|�Q=���<��7=%�=؄U=U�\�5�	;⋨�Vl<˾f�w
<5�Z�,�==];�<38"�9Ą<-�<*D$����/��<m��<4�3��u���w=�R��c=��ּ(�K�7�=׶��)7�q���<[c����;���<k�*=;�꼔U��=)�����E�$���v=�J�<�
��*B�z�&�zGo=�'=�|�9R%)��,Լº�b#�;Q�:�uQ=Fd���<R\���¹8�ü�<Gf��P"��;$=���<z�;=I����3=��X��T=�;V<=N���+�;(�`=|߼�	��,��4�;�FP=�P3��.���t�{�����;U��W�6=��:�2��=�X��#G��<�$+=�G|�B��-����<��=�����I= J���VG;#�G�"�9�2���-g<L�Z=�$�<�j���}a=��=�O=����~���,<A)x<Q�<?6=��P���<3Q��C=ɇ���=����� ^=��<�zm�F����}<zL�����E�0��<9�:��U��vc��+
=���<7�Ǽ���;�-ļf�;~��^.�OB�=F:8��%.�Q�=�c�u&=J�<q�=GZ=�?��#{B<�!="�;��f�<���A�4=�M�<�w�yZ8�[��;%�[<9R�=i=L��8%��O3=��ļhmȼ�=��<!#=t�A<�s(<ڮ�<xA���{�y�%=O#+����;Ĳ3=$��<���<���;��H<0fK��_U=ܷ��4��;+#$���0=X��H<~��;�P�("��1�<�d׼�=�9��<}1���$/��{��ػ0�=Ց>�a>�< 0(=�[=2�ʼ�#���];U�=����/4=�48=3�<�h=-9��8���:=e-��'c�I瀼O�u�JlM��<=W����:�<44�<��<�����9=�MH=GƼ�=����?m"=���<��=��R��w�;j45���Q=��P�{<P�<^M�<�P�<��U=c%�uk�<I����,=q#=���=�3h<E� <1 �<��;;���"c6��7X=v�μƷ=16���=��=i�Z�}3����<	�p=��<Z��ǯj�����ޘc�mEI�*�м��`='N�U&=��:=�Nc=<tO��A =��O=��ȼ!!���n=2Q�#��<.Ё;��Q���X�Z�P=��N�}�;��~R=r~8<0.���ST=� =��y+#=j!�߀E=�HҼA{E�J݋;N� �E������ݼ��<��:���<,#�
������.4�[�z�"�<:_g�&����d�u�P=��^=D����A缒wQ=�q=J(=lVz=�����T�������;�)�q��H�e=x�=��<S0@=�=<��b<=D�<�K�I�=`�j��=�����<��=�K���h=pr ��J���$;���V�$=���<�0��1=�6V=�)5%�D�
��;���~`���=���ǞC�B���B�7�����d�<9�׼.����<|H=�1��=�\=�ڼ��<K�c=���<���nk���f=iAJ=���<^4=j�=�μ�
H=ӌ=�F=�$��v>�@E=c�&�)�M<鳵<�J�<��%=��<��L�U� ���<!<�a1�1=�<��=�/���B���<�K*=�VK�򼻋wH�i�-�n8q=$	o<�
�-Lڼ�Q�<I5�<�V=�y⼿x���T�:z�+�b+�<��<I>����1�Z��<B�Z=�e�<��8��R�<��#�e�=/Uq;�>��Eܘ�]C�9�m"=\���yE��ц����<�c1����;�ļI�<����:,�:8Û���<t_=�WE=��$=D:�k�m=�==�����=ڞ5<#��Ұ =�l�<ڻd�!w=��/=�f���:=29L��<��a�q��N��;o<6~_=s T=X]~�V��<ђ=71�:�m�<rI�=^޼Q9;T!>=Iv�'V��H�SVM=�S�Ɣż��i���.�:�绛/��6ڼ�^�<�n-��Gۼ[����ϵ;�Hf��?=��=v�A��\c�n�*�]��<X̻�<�Cw==.=����(]�:`���>={�p��C]=@�]=G�?�ʛ���Y�<��V=X�c�.E���>5�k�
��V=���՝Z��=<���<
:�;��<7b����=K�a��JF���<�,+��I��IY!��~ټ��d;=O�<�=�G����)<y��<դ����<BSU����j='��<�@����<��=��Y�d�4</�2���)=�.s=��=,�_���1(=v����M��z=���`�[2<�T&=�r=H^��[8>�����|���/<�צc=�<cʄ<�9�<"�5=��J�J ���0��6=:��WzB=\%�<��*���-=�F��N�;��/��ߨ<���p�v��<�<Aɥ�azr���;XRH����<��<#=ܮ0;%�����)=lG9<3%���[
=�1p=R[=X^�a V�'wf��}k�>�G<�僼�D<���<*�p=*�.=�34=�S���y���<z���O����<ZD޻þ1���<ޣ��F�����Bx<�C;�{)��IM=7q�Bx6=�fw��X3=�,=�=}��(徼�.��qR<��^=1�:=�vY=!�:l�s=�c+=ՙ2=�#�;�����:�М��C6��{�<�s=]�"=ǅ<g~�fZ� W&�κ>=��|�^���\=˳���ö���ѻ�ü\h?��N��Џ<A�ż�H��>=`k�������j��7��<8����q<;��<)A=3䯼���TR��^�<�����<�Z=CD�Jq�B1��)#=!���yoo�;=�=�j�=�t~<��_�*�i���B�B�<j�=5Ӽ�%u=�#���F=���;=Nk=�p=0�;��,��U4��,���$=�Ϝ<3��;d��_�<�;����8�<)�Ļ�@I�pr;��$����;!X��I�v�<���<�'=rW�<����Ӟ&�V�R:�s =��<+
\=�E9=��!=D����U<���<@�r<�*9����R)�<��i�
U=�g��1�L���!�8:;;^�v��N<Jʴ��6'=�L�
;��R�&��=�hջLH����pX����<�mG<p�;�]<�F<��<�"¼{���"<�Z���:����)=H��^�$��=�i~=�-6��D=�^�N �;�{X=q�=/���P�<�L=t>H����<�黉{m�,T�F>���I���1=�v�;��l��u=$�<����ߘ��������L�<�X3�B�= ��<��-=v:]<w_��񉽶Ԙ<z�/=]�=���;��^�nK=�:���+��Fa=X��m=�q/��v��;MW��k�;��m<��=Q�=�-=�B=[D=n)�<r�=�L�'={�C<H��<=��c;	<s�z=�H���@;����;�L�;��<��L=]	�<�]���=��$�&>4=a�<[�=W�>;|�%��"�W����j�=��;��4*<��9�t9<]=:���J=�}&��)b��Y1�\4=�P�z�|�~#�<P�_���M��X=�iy��7�<t^ <mI"=a����d伉9��gJ�CR`=��r����<��:=����M��:�t�<�g=��=�;�\<�x=�6=�ɾ�ѹ�<`=��V��1�<DH=�#�'{r�j��<�G=.�^�\*;�`G�;^^��@=�&3�<�<=���<�h��
���8�=3�B��� ��T�<�c�<�=T�S=ל����7������>� � =�m�Tiɼ�b=r|O=�<W�D<�<��%��;e8Z��7��~�`<��弡/"=�<���ߦ1��-�cw0=�g�~⼗Ǿ��ۻ^�Z=�=�<�������xv��l�����<v7=��Z=�|����<޺�;OD=K����2===�5<�;^�(���d6=��7=\"#���= �R<&3���/=��c���:<��G<\!�<�T=��5=?�(��3M���F=[�=ွZ<Ȝ��JW"=�%��䬼1",����z�7�=���}A�ڼ�{9�<��1��28=���<���U*: �-<)�ؼ9r<Jx�<X�.=�3�3�8�yD<��7:�y�mFջY�P<	�)��aA�8m�<t�"=��L=�窼[k� ]�<t�꼬�<{T��@ �<+׼KK=��a��-O=�3�=�Y=�)�Q=Z�^���s=s,b���=����i����#=i�<�L<��|@�"@=]�=+y��e\�*:i����H�k<k`��a��uD<��K�<��<��<^g�Ҳ;�6=��F���=_/ �e��;����|<��=�͂<lS��2*
=�l����&�wo<=��=��O<-����=g:= �;=��>=�Z=�������<S�<��G<�2��!<� ��|U��IF)��:�R�:�s�s:��g5=�+�=�B���Eb��Ǆ�~s�<qC�<| �<P��<"3D=(O��8*�eN��[Z����qN��L�h=Y�N=6KK��fb<��������t����Kc�&��=��C:pi�<� �����OV�<3m��XK�m�Ӽ��<�EE���
<�Q����T�F��<%ᶼ�
=�=��N�(�y;��&=��4=
����5�!�c��N�<u�D� %<�{=
��}�7=��=�~�LY��~d<�a�;%9׼T�;�K=���<�Zg<�;E��<F �<�����=�.�=�i;:2�j�=��+�}as���2=h�<eun��^�<u~ �>�u;��?�Wl=�2;���;�<_3{= u�<�"=�1@=�P�<^෺�ݼe��.R�<��_��zQ<_k����h�4=�}�*]7=��@�@W�A��U�d����]�5�<o!,=ѼD=�<�2�b�U=��N=��<��'�x�{�k��<�2<�$��vAO<�M��~�z��9*�P=#k;N���*<��뼝i���<�S=��\�'�p�?�y�*�B=o.�<�h=0��;��<=��<�$T=�c<��<�8�;:����L�V类�s>�Z�I����
?��V�<�7�<��;�m�<G�F�2��>,���v;��<BE�;Lݦ<O\C=2G�<"O��ݐ=m�Ӽ�+<L��Q)�<i����e��ۉ<�5=qy��9F=I7<]��<�
S=g�d=��H5T:��=ڥ�
�L<�:J=/��6ݻ�T=cO;DIF=`Z�tP,<�����Q=0
�<o�g��ڌ=�6='nQ�n�����<�:q�yC2��X�<��}��M�#�c=�y�:\=S���<�g���z�*#���1<�K ��͖��D7�_z�R�=.��<(�<�I��q�\���$=�I���<�<�Y�+��=.62=�X�r��N&�<*�?=�5�.0�<�@f���W�d#�<��=4�<�+��,TP�X�f��-"��'�|'�<A5�=�JH��t`<"!�C��0�I<���<��K=��!<�u�=�A�<\/8��R�<��)=��Ҽ~E.=�K���<֑=��<񪬼@�<�|=B��;��=�zռ�=��@��t���<:����j���(=�Y=��^�z������<�V�F�:���޼�c�<�v=���<�$�<��}<�i�<�|�<���{/;��u���<�v;�Ț��sg�&�<��f�V�R��"8���z�<�D=v�N�|�y�f�<ii<?ܱ<�)��=�4tc�$�F���<o��:ם=�r(�̓_�R�&=�t
=a�	��}+=��<鍰<�Tu<�꺥�K�m�<��;q��?!=��;�Y�>!e=���<Ҽ�c=�Y��%�����_Ɉ;�
E= S�;��n={�P<SI���B�<T�=\BG�����<M� ҍ;?9�a/�y=��,�~�+�ʊ��O=v��<�i�$0=@ =�fx��*==��<S�I��L�;��\;H*��bB=��6�����@��}JK�j=�<�J�#�k��5������a<7Ƨ<��]�#�L=r��<�N=����m��O:/=�9��Z=�-l=n��<`�k�?�i�bk�?xn���<�0;	 y=��1�֘0=�z=4�������f~j<(�.=W'��w��@�:9�2<u�̼��
=��,=��A=kp==%�<U��<�g�<)4G<lh�<wkּ�&#�w�_�^h9<9j=�]=�e�ո8=V'�9/�w<j�Y�E�"<d��<x���=ȼ�U����;&��1F�=�T=
{K=2�N�I3��j�=Qio<�y=Md=�XF=�J"=[�C=�+@�$y��<r�;�"U �Po�<�=��=65<�nUq;��P=�E=X�m����ک&=Ƙ���:˼D��wT>=c���:��uN=�V��X�=�Fe��<P43�2܈<�}��
�< YA<��o��x`9\_#=�C�$h��aX =J�"=MV˷4�2�a���*��cC��X&=,�=�����=���<<:G��<�~�=�쬼d��<y4^=��A��l���=x�����=�ы=.�߼�\�Y�A��Ѽ�_D=�;�U2=Z��<HJ^�iU<6�>��P�IҢ��+���y;2rr���<uk�ߤt�'�^<��c�<L����帐���="A$������43���޼�u�p-
�~5=M�-��y=��a?�EQ߹�)<4o��b�������<uq*=.��<�9ü��=l{B=C��<1>�:�=3=� n9��`<���ˮ�<��Y;H{K���:�!j�;�j={0��̏<�w���;|�;R@(��	=�%@�9G<[�<�u̼
*��4=�[�1n�=j�:�F=v���j�<
�v��g��S���uм�E<�F
=�cۻ]�&�ɳ�<g�'�����}��7�;��&�y<4����==љ��>J�8,<��m�-���$�/����l!<ڤR=)hR��$=��9=�R.=�M����Ǌ�NH����@=O6<��~=($꼊C��� �T5=�|���F�H:�v�<xe)<�t�;��<�Ќ��$P=��H�T,�=h�=O�5=w���)=¼7=��=�V���ϼQ��bI��^�<u���s*���<��Ǽ��.;Z�=U�!����<���<��O�˔��t2�;死�y����=�|Y��3�;�K3=A䑼;�<Z��kw�l�=�t+���D=��������;j=�σ<M���	=S}<<�����r�c[=��q=ʵ���I#=]�=C��<
2F<���<�&�2L<��D�I�=?��<�$=���;���8�����i=�h�<T�;=�Ƽ=:<��ng=O�<��<�M��)Q/=C�<<�b�m�j=�	g<,4=C;d��ĉ<����t2\��g���;���n�^<z�U<�U�0�л�*�43�<�y��;}5��μAns�|J:�**뼛����J���<M��i�<��L ��=��d�N��1����u��,^�I�5=��J�(�2=��E�X�g�6���$�;E z=9Ct�ѵ0=��-=��<��=��=�FU�b�Q=���;V�J=�-q=`��<�uC=
M��)�Q�=�I=��n�lJ
����%�;��,��W�`Zպ���`Z9<M(R=nr�b�m�l'A���=m}k<�7�,ft���9>�<޴=�-.=pJ�0=tm����<ц�<��=�.�;I(=c����<W�����2=�i��F<;�Z�:�S����>�i��.yz�75�*��<��k=�VU=�����<�F=tif=o,,�j�5��"Z=�%�ij���m�k�=_�<�8���(�RK=�µ<Q���<##�<��d<Z��=��0��Ʈ;�3�j�\;3�_=˪���4ռ�}q<I��<�+�;7�b<&93=x��E�IM0<�=xz&��,0��d=a����=�/=Jlh;�c#����`��=g�X;�*���b<N���=s^�<k�=�6T���8;~�`����<�G<�[)����;��"��v=6Q��D
=����l6<cxC� �<w|�;��h7�����P^��EN<΃_���;�ݼ��D=��o;��� \
���8=){W����;=v\��"�`<�d��Pb�(�!=���<zy��>V���<r,:�/8�����e�<N���t=����5=���/���
�<�`=W�=����ijd�!mL=���8@�L=fb=��� ��<�����!��q�\;�^`=4._=�b =D�6=Wat<�q�<�w���j���=�_��J*=�$<�sS<�  ��T�ۢ<���<��<W����'f���<K��D=r=7�6��5�<���<�HM�PÏ��-�<����<aQ=1�ܼ�j��[a<���(��u�:=ŸL=�7<4Y�<��C�:���<,�(��&]�S��:x/_;Y�B��nJ�Ӛ9=��h<G�<��û������	��ü{wh<l�+���u��K=�<�Fϼb�c=v�=j���/l��1�'���=>��4��CX�;o��<��=����f�<��<*��<Y�?=)�H=�<:��1�<��;�m��L�=���<�]B<B���FK<�Y=�qw����#^�7&�9��|�ZX%�Ɂn�rW�<��c=͡�x�_�OF��"�<s�<�������ǘG�}�/=&z	=X�9�5��=Y=�s���ּ�zn=��鼥9鼴�==��:\�=��_=<Ԓ��l�<�r�C��$�� ��i+����<��o9�M弼z\���6��s0�|�<e�ż!+=��<��&�<��?��*<��<�.�<BE=�F=K�����<y�<r@�=��<��=4�F���<<�:=�vs�����<���=p1ټ�W��x�b<-2��7ŀ<��$=@NA�-S<�]�->;�a,=߭ü�/�<'�Լ�; ��<��e���P=��l���X=	�`=i���C=���&�;@�<��&=|�=z��������<���)��$~�<�BN=�g=ϒ�ݳj� ���a�8ކ�(�,=��}=u�h��6<M0�<��P��� <b����v�0��<�ü�"O=O@1�d�[�o2�$�2=��<7)�DA%=ח�~tD��&=h犼�PL���G��
M�l�7��=\=c/c�gp���>�4'�:ֺ�<���~��<� =@!I�<�,<O��<�tX�f�g�c���Msk�	>=�Q���!�~��<����;�����խ�3����/=�8<��F=�;<{g�.Q<2�E=��M<t=2=Q&��VM=,���N<�r=،������ƒR=��Z=,��<[<R�1�5M=s���À�;Y�<C�~���n=_(�<hч=nL����<:tk��\7=�{�:]/8�
�j�.c}9�B��W�;���g�Xcz��W��Lf<>u����_=���9�Z$=�Ѽ��=Г��!�;=dNѺ���<��(=�[n��9$=N�D=���=XN�<N��;�Xy����<��P��:�:G��<`=6y�AiT=�1=Y�l=��=� i�,E�id�=t�_�>�{;l3<Fc� @=iz��W�=;Zn/����<����=|p#<Ժ�x��;L�+<ݱ��u��I^�z��;	[G=Lb�Y�<)�<��=	��"�=�/Y<�_�z<==P�y��dz���0=��?<5�ݼ�Y��좑�	2�<�+=gfL������μ�`G��6<�C��b�?X�;�����F�=3�ż����]�<��=c�=�����<&4]=h�ּ3I=�A <,u8=�Xf���@�]u�<[�;�Ba=��C��S;�&l��}����t�M�<��=�s-<�o�4Rf=�'�>�q���<ާ#<�o=�u=B�L[F�aɼ9@O�$x
���I�����F�<d���	�c=Q��Tk=�1�<�=�!�;RF�<��.��$z�j�N=�"M=z�G=`���1o� ���(=(
=��K��L�<��<Q�M=d!��]Y�Sxɻ��G��H=�F=טT���;i���jOz<�ʻ�;<�qn�i��B�<w�\�r�&= К<@�#=]�"=��k�C-�J�C=c��<�Gh={��<Q�v<�M��P����<�M�G�;�u���R\=����O��;�P�G�s<�^@�nY���_<��=:��<�o.�҉���<ȯ4=ai0=�	<X��<03���b�ֿ�</=EY�<�ػ�A�Z	C=�;��:�<��9f<�̇;���:b��o�v�=��V�f1�g^T<|�+�'�!��ǎ���/:�� ;��=l�<Z��;Sռ�+��p������:<�o<�(=� K9Pm�<�����=�LG�XX=:��E�:A�<��X=~yH�D�Q�T�&���;�1%<�A/��Ԙ:�X:<{f\=�t~��!>��������j�;ϵ<:m(=��%=�i5��<��ӼzB�;B��'�>�E�<g8�����C�><��U=���[=��)=o42���~<�;�j�r�^7ּ�\�<�B�.��<
{'�00���BU=�:=���g<c}G���2=fF =�_�<w�%=�9g�Iwt=�%<s/�>=i��<1wԻ�좼�J��Q^<:Ǽ�MO=j5��*�]9��'�}M=$_ȼ,�P=��:{T��LV=r��mZ��\���-��.�Q�<��'��6��6����n=���<��(<�H���_�<�c3�  E�ep#=�=�;�0�6��eC=Qٸ?U�;�'�7�;-o���<��U<.�<=�=l=b9T=���<OR^<� d=��G���m=͓��^��#�<���
RT��_E��ܼJ�	=p�T=��=��)=�<W�d��l=��ܼ����|=�}�;i��<�^e�Bg)<N���P��:����ނ��X�<9̪<-���\U)=L��ި<'�l=�b�<*��<6]�����<�9�:TCi�Lʴ��eC���<��/��6���$<���<��ǻ���<a�$�lG˻.Q	<#%8<�R<�O��8��9��I�]���Y<����`���*5=z��<rm���?=�\�`�<�@=o�=D�;��<��<'m'=[�B�mLJ=����ov��;���$ǼI�5�h=8S��	�G^=�-w� 	%��tػ�h�<��<8Ǚ<#>d=�S��)�=���<2�`=�*<���<o^N�`b_=�p�by�<D��7��弞 �<�BN��7�<�� =gZ��
=�\G�I�����v=�J��] =�XK�a�=w��<��=@��<��>�μ���;5�!<��D��S�=�0[�+�S=0`�<�.ɼom3<�G�;���;���ݱ<�F���o�F�2�9�=Wp�<���6)�<u$=�e���������;����B���]T�xe�W"��e�<�&�HH�n��;�nN=w�<���@�G�yE���<#���]<`j�=79�k��<���~�S�yǓ���<`�h���f����?�<-�����+=�km����<�*0;�7�����;z�==���
�I�jy=9�1�"��B�|=����b�;=m�>=��ֹ��L��� �K<;�㺭ɖ<�ټ��=��c<W�C�K'�X���1	��-�;�c�;���<G����6=�=�#��"��%^/��=���xmr�/9=�*A=��D��'ѻ0�T��)�5�Y9�1"=gMh�GP<=�K$=�Ԍ<���<_.��v��*�`�^3���7=��@�<��"��9%�:;�4=0Q= �:�Y���=$(<��@=ߎ�9ՙ���\�{;�:'��<�`^�����^��s[��=N�F=�$x�|��R\i<6����y�H<�sg=_<|��;7����=L6�;�K:���#`m=RDH���N<�:�<���<%�<��Q=�+[<@�<=�=���켂�һ ���h����<���^mg���-=h�x=a-�BN7= �;K7=@��:��X=�]=��E=a'��!j�W�D=�����:��!���Nռ �}������`�<|cz�-8�J��;&V�<�gn<Ь=���<P9[<�8�)0]=Px<=���;�
J=s=U����?=R���ؘ-<F�^<@d꼴 �U�k��ڼ��D���7<J��٥a<�yf<-=�h,���<��c�iZ=A�=��o�D�k����:Z���]���k=:�t���x<��<*2�:���;&��<�g��B�Ӽ���'G:=�d�<��;�V=��<��~<�Q���L=<-��<kk�	|D�fC\���	��8=h/�2�<�9N�<v��P�<BS<a=�;M��=�#6<*H/��!K=��|���%���Սf=D@o��}:=��y=<�)ü�]<Κ[�{��<�;<�*����<J\U<�4X=Ɗ/���_�*��LR4��=;�<��c��9=��`=O�%�7�_=G.�u!伛eW�"�<߼/�輷J���A<<:�	:k��<�� ����<��r��nl��m�}-b=��<�m2=���l������<�]"�r0!=��A�E���R�Z��`S�����Ua�F�S=�� �k��o�0���Լ�E=t\�<�P<J�����Ҽ�;=�\�.g�������<�Ec��T:��@�<M)<��c���=�6A=`X&��G<�I��i�A=�%��C�<=�o9#_)=�#���2����<�Rj�q���0=�n��vL�!R<r�<�)Z�,I�<~=�<�*���%�%P�/O;��R���Y<�,D����<J�=gx��^�<鍀<j�����>���eeZ��A���l<�) <&伛L�����<
*R=��D��j�������O=�ۺ�	;�+�X�[=��(=��u��<�&=�Ѕ��W=9�(=� =��꼅��<sY���`��=��;i�H=I.4=C^��a�>���;���n0#��1��);��=��*�O��<���y<��G���=��(�������L�P��<T��<���<n�<�'=T��&����<�3*<=��=OO �ڵ�<���<�=�?���L=	*J����:��_���8=���<��P�8�J����<�,�<蛘<P�>=m��G�Z=0��<�w�4�	=��D�G�ۼ/A�V\_=!<�<=Hj�����m=ip޼d=�g=��x�`s�:=㚼^�S�e|o=d�< pݼY�<(��� �9��<�>=.�Ҽ�2=!6�;�����<�)�<l ��gN�5�'�J;�H1�<#�t=���;���ǵ+��t=h	�"����X=Tq_��q =��
�R>=��<�Ġ���׼��1;I�߼��O=἟���fq=�@�<����k�Ȁ<��=ϥ����Z=8�@��z��~;=7	<�:�}��<I@���=<>�=�=��<�<3�y��j�4!�<H+�;��N<H�5�A;#�`���=�[�4v�<����1�i��p=�&��c�</�ü'�<� 6�#��2+�$U�:/�E�;�=x����ܼ�S<BF��'S��� ;�hӻ~[T����#�{�T=��żqSM;kɣ<b�Ѽ2f�y%�E-���)<�3Ӽ�0;=&kD�D���t�g=�ņ<!�<=�}K��J[=��s�v��r�_=�U˼�ɨ���=)k�I���D<�� �=��B?=�rP�F���;K�<G�޼��<np�<�I<ؐ�h�+=�X[=����'��?[,=�`��=;o6=I���QL=��<E���y���@���/=x�V= �����<J�6�n�ʼ0x<?�����V��:ԇ+�؊������eb"=Qv���w���TлV�G=�=r���M0=	=,C7�Qe%=�%���+������-��A��M��)*=ո#�Q��<��<߲�=�0.��j=�w<�V =�=B�Q=z_-��r�<W�v��J=�A=Z�3��V�<˭��(ؼ��C=�:��
�<A��d��=���;�̼�B��V�&�9���t�
��{=�}{�H"�}��E� =?1:��.�.�<=�^={��Y�9=t�O=�y	=����~�S�(��ؼ�w�m�<|�<�0��Z�<�j��욼����=ɉV��Y���m��0t0��B�=��1==��s���E��{=�U=e�$)�!�$=T�W�]�<�̙;�S=�ݕ���4=xV;�Q�	Z/=$��<�aj;,�L�G�9=󟠻0ф<`�S}h�]xt9Z�ܼ?�H�K�<=]`�&%Ѽ��5�4�@���$=�`F�������s�i�C���=|�u<z�N=j����üu��2�Q�=B51������D�����A =�3=u
1=����P�;��=��<��.�zc�Ѣ_<Q��<�ݼ���<���;�wG=��R=һX=�f?=DI0�a���+R��ڞ��4��NC=�k`�8�9�Z�����j �J��<
���G=���<s�<A�<M�;�?�=p��#	N=Y.F=܀��J `�!%6����<"�y�4�y����r�-F��l��Z4�=��;b~�������5�<<z=�\=?����<܋�E����'�k}���å<��7� �<��<<�8= <K=Ø:��<z �H'=�#9\87=-Oa<%�?=j�<Qτ=J�[�$#�;�J���n+=:o�={3<=�fI=F/%�rQ�<b�={j�<w=���2����c��$��<ۅ�����i�)r������y�ʉ��qp2=�I�=��t�}>���k6=��)�A��<�i���=�"�=��9��)���=+��i��p��:��#�:<�<1/�{�=��:���Z� <��<�g�4��<MY,=�Y=D<���;�(=J <�Ka�^@����s<������<�5Y�Fh>=�CY=���<���<r�<=8=S4L<�I
=5C���ּc-
��O���<�D"��JR<W^�<���_��=�<�9����3���O?=�
�`/ļ1��<�=]@�YfK�/�k��DȼE�e.<�����=<�缻�[;vT�<���sDP��^�u�8=�=="�=J�I=��h<{�̼�Q��`��<fly�O�4�-83=�����Ά]���=�%~��V�=|�;=$_o;���;�=%=�;�b���g�RŘ��[��A�z<i=��g���<5�#=b.��O���]=��<�$=�-��7�;��=l�5=���<P�7��R)=e�z����!�Υ��Ԭở6�=t�
���G���L=�p1<���`Gݼ�?�<�M�<s�䚧<L�)�'``�)��<rT=��V��f_;�����<�٢<��\R����:����>�ڲ<��=���<�k9<Pٗ<]o�<�������k^�żf�=�*뼝������< ż���;p��<^E�m]��lR=��=�-P�x�������S޼j����#�=�T=(�7=�@����;��&=)��ӺI�<�=�1O��=�g_���?�]��;� =�=�庼	=�e��=�� ��=4��<��=Zs��/�>=�B��RL=��&=���<���oy��|k9�k���X�;[v���!<�9M�l舼�Ȭ=���<��J�1�V<���<�� <|�<A���<������*c�Yi�<�?=ʬ���G�<Gb�����<�;�*̼��X������U={�M<�<�<S���&�<)|><���$��
q;dLA�*~)�/����x�!�;�&=D�U=��7�<X�D�����"=Hn��
���#��g����%�^�5=����!�<��cf�<uф���E�,��l�<ڜ�<�iܼ ׾<��Ⱥ�a)��i=:���!-=��������=t�=X�μ߇��B����U<m����1�~d=¸�<�I=g4=xYɻ�|*=E�^= _�<�L�<�X�;���<�=�#=�K��� R�����F��g[��!�<���<�=�4���a=O�ͼ�v�â2=p�<��K=�z/�gU�����.�,<X�z<�O�:V�R=f=�~&��(\;�r��jj��e1'�М��Yl�2s_<%��;7�p�.]8�hS�<~�v<�~�����ȉ<�R�:�=���;�=<�V=*�(��W�;ڎ	��88;��n����<�+=Ġ,����<O�/�J6�<��F=�7M<:��;иj<��Z=[ka;j�L<���fTg�ES"<�&�<JI2��=s�{�[m=�τ=�r=��d���	�;{�����M�.�U0��O�X<�%ɼY?�<�q�<��	��'�� �<T=]z�;l��<�5=�s�<F�:��b=�̼�]8�~$=� X�+xn���f����<�硻�㺼y�g�$*=�9�<�\�<�۵< C=�@�����m��<n�L<W�J�r6=qy����X=��;���<R��Zd*=��<"5]=�hf=���[R;E��+�����<x�Z�1@��2V#=%��;�<x>&���8���j=F(��}I�����iV�<��;sVg�6g���oS� ���O�<+��:��=D����^}�;;=+.�<vļ��;a���"�<p=p�=k2=�ז=��<�u�<���<�N
=Y�R;���;("����;=T$��T�*5���V�'�O�d���������<��fP@��
���w�w��9!=��7�u���t�R�̠��V�_��E���^=L���x0=Ȧ=���=�,Q��!����0���ؼ��1�ã��ͺ<�U=�D���_;�a�<l�C�Ӵ*=Z¯<��4�
�8=h�#��B�<����6�;�f�D��Z=� ϼ�Q4=��E�@1�dr=�X7=����YG��D� \�<��'�9�u<�,�;_@�<���3~=��;��=�,�:!�b*Z�=%#���M�5( ��_S�J�J=����6ռ�4;��4G=-
h<ޅ<��	=�z��;��<��;h�;�?"=9�=xI=��;��=���<� D=��<إ�<�19�va��L��LR��)�8N��|=�t��T(M=�4=��E��V�L���`����]-��i?<[�"=
��/;�u��xW=kDB�a�<y�w=l�=��U;��tN]�a�z=,�m;�5-���p�+�%;�<�_N=��=�B����=p}=}%�<p��K�L=��#�ԕ�;�L/��a;���/o�.Y�<�V㼁P=�<�F�5�`=
��<�p��]<��~�t�=�nO��� =��<�����*���(=��<���0��a
k;W�<O�~<��Z=CN�<Ȼ�Ƞ�C��<�
�=��;��"���L�J�<B�=/��9��V;�;��^�rOJ<?X�<�-˼���p��<�hI��I�^�D�'�<�l.=3ļ-�8� D�;к�Q[M�����:"=
$Ժ����~�<�����$���3�����;�<T�=z�d��<u�ռ
�漦�:=�w�<��<�k����;cQ����<��":��<e�!��RC;���YY~;hC;<���<�-8=_P���<}�$�xF=�'�<��ͼnr>�� �*�E=)<�<2%=�zм�=d�����Ƽ��W=���;�rӼYڑ=I�^��R���G�xT^=�༉0=�n���f�s��e>e�g0!��~C=cG���FM<,�F�1='����~<�����<��:������}"=�^"���q<h;�"t7=b2n�؏ؼ��s<~M�:L�!���d=�z3��(Z�݄(��1�<����A�pEU�w*�;��;���<m�_V�<{NL=�$;=�d=�$=��L=��L=�1����Y�g<&���7=Za;=,F���@�QQ-�h�Q��=4x�;xB=�����=)	L=�IZ<#�n=S⹼�=H!�=_^=������ռ�%�<�;="^6��\��e^o<�Zջ�qQ=�4�<��;=�2`<k���M�I(��t�<�{)�K�E=�`����/���;m��<��R=l�<=R������P�<�R*=L�=,Ѐ<��̼Sx=�<���;o���<(���:=�� =��;z�4��¹E�<B�<� �����;�m��=�@�fߑ�.�j��A�'=�eK=]q�č�<�28=
�/��*<F���l�	�U�۱@=/����������K��1W�%S��E�<���2���$���;����;�D\=�5��
�<Ix�;6)��ἕ�n�U%����eƸ<~�׼X�=�Y.�f��<p��&��<c�<=+�X�O��<.�<U�<2�{�ڷ>��D�<2�>=0v�<�x���=�-1�����)�����H;"/��I�<7h˼n�'��<Hݼ��=W�<8^V����=-�޼�vH=�Լƈ�<��P��Ѕ=N�Z��6]���7=sGF��a<U��>�P=3�= ���;h�_�W e��q:=J�=<�叼� <��_=UQ=�0n��@x=���r�Q�&�V���,=;�c�53=s(=R�C=��@=��l���"���!���P�/�=D�=��?��0=��<&Ѝ<� v=U6Q<'�/��y&=�W�v�٥���Rޔ�\��;��]g:=�:�<W��<T<�k�<�"�<:Z(=�j�;��W��Dn=/N]=��Ƽ��:�ij<ԨI<מڼ�dI<����&%=�[;=k��D����|a:S2�LhH<�}=���T�;;�=q�H�m?Ƽh����<%nм2:żIW�"�<O��<N���u;,@)=�\��ݻY/�ӣe=���& �<�Ϫ<���/=��� ;m�ř��&l^<�Gڼ1�����72dM=�*.Ѽ0��缕<ˊo<'�6<{m=E�~�u鈼��8{��a�L=0%���Ȁ<I�S=b樻���[�%�I��<�Nӻ��:<�Z���`�z���?�0��<�-������C=�81����<a=���<SXK=d`ż��o�r��<Q�q�x�Q<�X�<�C#=��<�#=D�?�_�]<0�׻��!=�u`�Q��I|<��	=s�<�i3;�p=��_=^�=}��*��<�V<8T��G򼂶���=����8G=�5+=O���|=i�_���3�R�=�Q���U�v���So(=��k�����ρ=�t=&��kP��9$� CD�G�P�];����O���]=���<&,��v=x����׮2=����5V��A�Q迼�Ё=r�/=��B=����'S�={�<��L=\��<��D�!"Ƽ���kM�$Iw�נ�<z��<mE#=p~�;O��<,A�ٰӼD�g���R<����&;<YrB=����ļ������Y�$M�<�7��N�h<�M,=}�=���=N��2ܼ���(�~Լ���@����*<FÓ=���<��<��>=k{����<՗�<�]`�AN��'w6������.6���<�ȼ%�2=�	=���<G�a=?I�9��ʼ��%;�%�<�MA�k�;�OM<?�ϼ#+=L�9<��=���f<��t��P/�T~�Qu�L��<da�=&��bE���b6<��|���<	�Ѽ�		�/�b:��!�o-�os=o�;'�_��=7�[=�`��c�=�;��F,�;�I��ǡ���8�<KT���\@����<)�m=��i�U�Xü���=8�=�G =_B=���'#D�K��x��;�T=�̥��T���<+��;��B�O�ۻ�kO=�!����d�e =|7�wm�퐕;�J"����:�,��<��$�<��< �!�v�?=P&����ټ9��<hA<w�Y�+i�<o�6���o:�Y����R��y�,�bR�Q!=����������!����<.W�ց�<c��%�<��`�H�F�$*�< ��<��C= Q�K�s=&�F=o?=;H=��)=77�;WOC��z���j�s�j�1�<�JX�F����c=��a=�B˼�_�<������<T�F=-�v���96�=cd@=�e%����<Q�#���~�"��B�=��:�5!�ˆ�<8�b�#A�;2\��m�P�X� ױ�j�ڻ��)���G���j��3O�0��;��O��d�<T<ɼ:���K�
���(�,<���<(x<�_�$��k�ż6\��P�T���<���<B"m<�Y�;�d��3s����"<(_<�&%��V<�"ռ����'ܼ�&�����<i�=Vs�;mU=gA�t�����м o]<z)%=��$�r,��[86�Ց�� =�}i���-=� ;:�u�N��<%5^����~V=��U�J�C��o:���M<�����,;�'��|9V<�<�n��w=u2.�c�żgü�=��<��M=]���A���/�v՗<^���i,<�&8=vW漈�m����=�e,��nZ=yo��3�,=5�:򛗼Q�0=��l��S=��B=++=o�4��B�9>� =��ܺiC=�Kf=A��<)�L=���M*�8μs�I=�8=AdQ=Ќ6�un$��
���,�s����$<��<��=��<x����Ƽ/{���"�=�	\��N ��F�<�W�O��<e����:�=i'!��o���37��q�����<��<�=a=�B����ZEZ=��=D_�<��< 7H=o�|=!X6����f-?<E
���W=��<��=<���1S�]�\�ƠB�^������:
n>=�p��C�����: ET<_�<�ڷ<K��K��9ai&;_qP���<����<Oּ��=gY"=�0=v䡼#��:��*=/؊����<���"��x�<,���&�&U=@\�<19>�b�e=ab\=���;nnG��"	=(8<=����<����Q�u�C=3$s��B�Q�<��(����{�=�� =Wt1=���<����l@�E�=n#��Xx���)=���<������=a�؄��y�����wo���<S"��O6�1/��E�;��1�3ޅ<��8��c���=�A��C��<��k�<����I=!U��D4=��(��B�;F���l=+;��m=���ɺ�<t��=Z��+#����;�#��K��<�v<+=��0��"f=�Fm8	l\=�٤<�!,=�#��h=��/�ڼ\�ü��B���ͼ�6��d��F����=~V�<�_=]�׼���<�8���:ʼG�?<�z�<0�<Gz:�{��`��:!6��Z��<��;4�r=e� =��[=�<���2�W�5����<n�ܼ����7Y�`V���G�_�7=�9X<�s_�7zO=o�;*1��:K�d�hf���Vb=7���E,]�i2�<�I<�G�l�<����;����X'�<�"?=7�~�6=PY���4�;W	��z�E�h<�~<!V�<�v���|=�!�9���X�6;I��f'��{*=b�M=Z!�x�<����;�f(��u�G4ܼ�4=���"CL=�:(=��<�0=B��,���g� ��<�7X=h��<i�*=��;�E��Y��żN�n�[��<(Q�<󼼉�;$y�r@)��!>=m�|�����P&�D�;��;Z/��r�Y���<f:��< &!��-�<
=�Ϻ8��ω�ޛ��×=��<�N� r����<���j��)/�N�b�C<_$=�_�bMJ=������</�K<�<x=1�-����;�W����<����V=� <x������U�0�e������'�/�
=�ϑ�	����=�@��0�l=�G��o,=I�q���i=��*<������;�. <c{F�Ĉּ�M;�(R�t���������a=ڄ����;��1�Ig�<�@�q��0���=�8=�'�q>�<d=D�)��U��� �<��<㍽<4��7,=�J==��'�����=��P==7�伟Mh=Ҫ=ݐ<kﯼ`�<	g=�1żum�<9����`�=?��J�I�T���~����E=���3�/=L;���4=���Y�����<��U��9}�<�<�п<e� ����g�K�;�X+=C�`<&�I=Ơ�<Dl�i�,=;�H<b�C=/,-�>'�;n[��6�K<��8=��r���q��ȉ=ެ&<�+�=�:�ƍ=�ռ4�C=wh�ʄ�<�c�g��<We/<�'�<�!6=��$=@)&=Ѝ=�Y=S�)=I6=d埼Vz��B͇=��:���<O���cN���.=!O�9������z������=Yap<���`�3=�����=�;��+d<���ij ��4=�}��	�;=�.�< q4����<���<]IF��Gh=�ј���K�(�"=�\��Ň<�7=qy��N;�8f*�L�0�sE7�?w=���<�_z=�<"�d�LҲ<�d�;7�h<1��n]|=�
��%cJ=%e=ݔ弢�h�����U�M��<4o1=��<��$=hq�<m;=����w��yt[=���;�����M�,F�<X�=����`fn��v[����<��-=��<g�U���4�_'ἂ��=�:�;b���:?=d����<��=���=5(��<�;��_<	�E=�w��a��=��{=\g=��f=kˀ���H<b��;�8��o�k�)�F�M=��#��I:<J?"���m=�&�<Q��t0=o�V�J��<QV��t��a˘��ܔ�7P=<=�-=�I=\�:�?=� �;��B��=z��[�=���b�=���:�f�P����3ϼ���<}0ּ�<�s;=�:=\IƼ>]F=f =�G�<��T=;�z��-M�xE=���Or���h�������oZ�.�ռ,g���Ү<5Dּ%�1=ʆ5="MƼ1J#��=5��<Y=��U<�I�=�T���]�<�.��*;L��<�Oļzdֹ?��;��u<|#?=C���eO=kY�t�F�AQ��/�n=�_������t='pA=i=U��,k�v�t=�"+�FI�;�=�y�UV9��=N^=0j����<W&K�b7�kx¼G��zL���+<΋��4=:�k;��^�S�%��o�<�7C�����qk��7=��<�.�Ր!<ar_<�ٮ��0��)��L X=�2=?�9=�ᐻ��ݼ�r<�=N�]�g"=$%��|����:�2 <�}�� �<�+��dϚ��,M��lk�Q��;>=�3�<fX;I܏<����R^=-O<=�qۼ�ƻ�ռj��1Z�<*ZH���μnh���Ĥ<j���gC���<�ҼG�\=!�)��C=
��<ݎ���='�n�y@Ȼ���<( =���>�l�=  ;�,�<!T"=һ�P�ҼW^�� �</>]<�
���!��.t�<������;4CE=�.��:	3=U�{�j}=~��;P�&=Җ��O=��g=�*�<�{@�n�2�q|=mʼV[�n�X�=A�]=���;B�(���<��Լ:rN���O=��n��<ah�<?<a�ez�:�K=)�<��?�{=<�Ի.܏�c'���c��w-<-D<�D��5;E=���Hw�М<��'=�2A��=J<�N�-=�$�:/Ս<n��<[y���X<I�n�y͍<��/���<�-�ǼO�j�т�3�ֹ�I�<���<�����F<���pg=�~��z
c=~X����L <ީs�0�&<��r�·@=`�l��<��O���Ae<�t=�V�<3�=&|��?)���T�O�8=��p�8�E=A2��e�O.�<`���is�pt�=�='<Ɵ?���h�9|=>�A<c&���_<HY=)	c=/��:���g=��<��=eE�<bme=x��;k���o<�hԻL�y�C"_;W��^�Hi��yݼO���+m��>=�������Mg��.�<4�;�N��6�B=jn���5�g:f<��=K�.=�~������%=�T���� �<��e��6Q� {j=f3i<�x=�T;��������)��P,���)�d̓<�i<�n�Ǉ<)�<��}ż��l=�$=5l`����+�<�Z��SL=�S�;�P=���xi};?�V�Ƕ}=�T=���ƹ� q�5�=<���y#=$k2=�b�<k�=ۚ\;����J(��[=�[Y=HO2�<�`��� =
:=7C=�<S\ϻ��I<�Mc��b,<�d����������̓��l�<�r˻+Z����Iޗ���d=��<��=�)=�G<<w�?=�m�y#�;I�<Rx���=��<���<��K��,X=`Ğ�L�;�	�=�k���
��צ��$�i�F;��<9n=�>��y�u���_�ռ�Θ=c���
�\=T���u�%#ؼ�=r�M�<9�=��s=2#�<�n�;'8=x�����;r�,=�Z�6�;�˟	��4��A�=�no=\\��]e�<����TZ�������;��~p����<���<�5x=X`�<��K�|U_=6�=]��;���˟<�ـ��ӹ<�KD��_P�I爼�\�N��������������<�X��D����=��m��m��*�U=�Ї<b�4<��X�W$��v��8hd<21����<9_=��=�LQ=���"�@���}=����a<=������0�R�!�������&=�;�ѹ<�c�<�#�5-�<'�¼v�<�IO;p�V�s�\�?�׻��{=s�D������X=���x�R�\=��G<S{a�-;?<zμbkV�5t��m�<�٫<��ͼ�i��52�S+S���1={��<�:�<Z�<0�`�0"���"=�0ļ�CA���c����<F����C�5ꍼ�D<=7����<��K������<탔;�g����<�X�N8<1 +=�pS���:�9�.���PW$��`�<��_�g<ٞB=M�=+�3;�s���=���;2X��L=X�-=�<��j=P�ļ�,A��d��-K�;�-�f�<�S��)��<#.=?V�e���Q�$=3��;K�@��z�<��&=��L�5����U��kQ��=:�F=d��<J�	=�.	<�v��>y�<o2�<�s�<`�4�ټ�W�=	I�9=��Z��=�V=T]�<�N=��k}�_��<+�׺+��;#[>=f$Q�4�F=�e��t ��d��up=�F��*�<�x=4�<`�Q�� r=���<�ܼ���y����Y=� �;��$<�la=�C0����ʒ�<�Gq=�c�<*o=�~�<C|s��=�<�pR=�Q�Z�F=u[d�hӥ<�?����;p�{����<l�<���<��<�NR��Z�=��x1X<H��y�=[U�0�����T���<��$=-�E=K;��_�`;gÔ���`�kvg=v=��;�=�mu�=�A<�QM����*=��q�p��<oY��J��[�=�_I�E���G���,�=���a�=,!��^*=7��f>N=�i8��pl�u�(<r�����[γ<prq�)�⼾�ܼX�4��8�Ը��Lq0<
��<��6=�ri�Rs����t��,==���gv���ǻHZ�<h���@�<��L;?�_��<n_K=N�w��x]�u3׼<:�;�WԼ�惽�+�.�<�wH=i�'<�c��Y�;�_����,=��C=��ݺ;F�<w!�'�<=�&=��E<�#���[@:΀<�=(��;,D���f=~��<��2=!V?=䆉<��9=j]���
�:o=%�_����&`=�zf��)ؼr��<v�����<��+20�w�X�x��< ?,=-Ly<�e��؟���B��v�;F�/�V=��ZSF<}�(�����n,=S=V<j�T=-Ǌ:Z�޻�9i=?�ϼ���\�=���;�d=�S=��e:�۶��c= 4�ǘ�:��=�b}�n{:�}3\��O==�=?2���.6�QT���{� g�,���=<�ۍ�Q�U�<% g�2�%s�<�`=8x4<·i��lQ=^�!=�5�����ځ�;}B�����K�<�MY��9��dD=
�={!:�KF;͍�< ���IN���EH�=�O5=�V9=��8<xi�<i�<��ȼZ`
=��t<G�;R��j��<�j|=�<��r��L�5=�L=�g��ƭ�*�x<n�X���S=��C� ͑�m�;=O�
��)O= D�� �<�+M�n�+�ƾ)��I�<�t�R*=C�a=P_���W��3��c��;W:�8F��|M����<�_�<��*=��� �<4�.� �b=j�B��R1=$�,=�#<A��<��%=�d�B�H=�C�=����LA<�����>=%��qW4��);���<%�Q='�I�R�U=�X�<n�b=�B1��œ�0$=e`	={E�<|'1=���Y�0<�i�; ��lK������)�f�]=S�M=���<4����Y�P��<gu��of�:.�!���x��UC<��=����D��8:�<`[����=�QüxX�<�f<҂�;��T<�lA<�=H���Ҝ8��T���|��2=W:�^��=7��l,y���Z=��;��<錽x=-�=*��r�<RI=/==��3<gi �9�0=p}k��=��`�<�B/��C/9f,==�ּ��|�J**=n(K=�5<��<��8�M�yJ=Dį���F�}�I<@��<:�<b۝���1�k'�:ك2�6Y<d�9;�+�?��<�9<Br�<�P��#h<b�ы�ި=�5=.�3�s���i�9�{��¨<%k�x�J��yf=X`$=���=TL�:^$�i{?=��<\F�s��7�����0=�Ȣ�zT�t�*�Z��<����I�m|<��[�7*��Ǖ<�Ǽ�= 	��O8�����X@=�6 =�X��7�<z\��ž���� '��Z�=~ɐ��u4�wڼ��<�g��e�u��)�<o<�3E<����eR=I�2����<=`m@=h=7�;=̻Z�l	
���<=��=|r==�h;(so=��;�0_���A�9�s���f;�/Y<�t:�(�[��߄=�0%��"�:���E��a)<���(��<V��<��ռ�}=1�`��jK��s�<�q=����̼�5�Q��]�E=:*�eBϼ��򼻓9�7�u=�i�<w�6��=`��;v��<̑=�h<%N�1H�<�_:�Ò<�'=�n�мKt�<��<L��<���� #ݼ���;Z u=��J;�G=���D;a<�v=C��B=ʘ�=�:^=H+q;���<a�4�"���i?����<E=�<�UƜ��V�;T=���<p��:�N=b		�35�;����@����M�F��<ּa�YG&=?(=9<ܼ�W=ھ!==/��v��.���?o�<鄽�1,=r���P�<��9����:G�=�w<Lh=Y�7�k[��׶���K�������<&�8��
 �;��a���<3$ؼ��
��BS<]j:t�ƻoO	=�<�o<}i�<>���\H=���d�N�{=���<z�O<y1ʼ,�&�'���oK=�X��5��Ic�����ϼS�X���I<�Y7=@Y=-A��99<&$M=ݙ9�������<�<�t'=��:�@;�c4=���-��M�e�f�	=���<R"��ؽ�<Eu<=�I��%�|�ԣ�Uq�< ��<8�<�Q�<�R=<"w��w��D!�\g��8���ӼE��5�<�9Z���I=A��r7�:0W��/�a���4=�6�<�yZ�YQ;EE�Wo�<!&=�� =�g�S�n��Sy���#=tp�<Fb=E�w�?�~<Ze��k�u���?=��?=Z�����q�өջ0D�=)a��̼��_��W5�%��<�=]�/�i�f=v��<��=ٷf<#�|=����?5=�z��@����5��A�<���<-u��實<�xQ���5=2'�<i��:����-|�j��<򈂻ߓ�: �;N����̼��=y}=�i7=��7�?��<��n=a�y:��S=�Ge��=@=6.D=�*�*���g=A�R��Í��m<m�U�G��i>�tT�<5��;T_��L���8����m<0��;�u��<k��︿<F�̼{�d<5+A���i�������|o�I�Y�8h;[M��RϘ=�@��F�.��<�z%<�/�9&�<ech��y1�\�b=���<�*�K4=�ȝ�BԨ<�T=���<��1�H����GP=۱��uDk=g 4�SkF� ��;����=1n =f�/<��μ����d����<��9r4=,�<W�<e5 =��.�Cb�<�T<=�o<��*���輔%��	|;1B=��0����.2G��=К�a��Q�l='Sg��,�<b~�<h7=-�0��]B�!_�<�
뺱̣<�����H�*�v!=�s�<�'¼=�Q�{�o=�Ţ��*�<4��W�@=!��;n%��`M��O�<���kS�ҳ#�Z]�<�*�m��;�J��Ǌ���.��sԼ��=�q8�����x����X<{\ؼ��<h� �̕������<:��;��M����<�D2=��%=F*=�j�ߣF���~=��I;֩P=qH=��<"s�<1-�� =�
���f!�b��<睵<s%мQ��<�.�<�+O����;�i�<k�I�l���"�b��	*F�#�*�|=ĵ�<<�<��<=n�<�`-�I}���M�<�W�s+�z=^է:��d��P6<��+=gv���(���#=�(<�zI�SDn<D��<�x<���(|X��g<��޼��K=%l���yg�y�(���=#�o����<�w�=��ڬB������)��?d��0K�;�=�ܿ�
����!�;QS�<@��<�囼?�B�i��;	�=݉�<w6��tB=��G��÷���S=����"�<"=RJO�M�!<��f<@�$�n�.=*��<� #=HF)�����+=�������/&=��a<	P=�ّ��d��=ȼ6��2��I߈<#���q�O�)=�)@���D����;��g=%�q<k���m�<d^�<�ʥ<ޜ#�욺<��/=0�"<�L��� =k�T���<ezY�}J����<��$[r�7���?�=ۭ�@-�<B�ݼ�~=������<������=�	<�C�;�(C=�q=������ ��� ��sa��T��8�V�e	=����¼v�ϼ��@���+��̅�� �<�=U�"��6��|=L�$���=R�ּ;Gλ}_=�}�<W�l=	4=��e�T���L��K��O}ʼC =�G8=�:�2�={��<28�(�T���=P�/:�[�<��<�"I=E�<������;�^����;ª�	`�<�B��a�x<��e=�����<.��羅��謼�E����^�Ӽ��=+�Y=�N)�K�69��<���;��8tD=u.�������<�*+=/�r<�4��=\}�<�=cn<=/���R���77�=ވ<��<�Q6=��),�=%�&=�  ��3�w-�.N����<�z='¼_@�!3̼3�=��=ZR);�C1�*9=#"=.;=��r�-A��4B=���=����\�x�6��R�;.fl<�|�;#H1���+��� ��35=mS=�V9��l��\�=��W<��J=�Wo;}�f<�<=S��<�r6=.C?=��0=:���;=��<��;�s#=��<�� ��=1�:<?ʺ� =���j��;�%�<�Ab=�w��=�/=f�;��=	�w;X^�2ό;=)軽��;'Mk�������D(<���G?�;{'��	=y�;��K��^Ἵ���o�� �+9H�'�t}P=[Ҽ�[���1=�{R=�;R=�";���~�>T�����ea����L���%�h�����'�����0��Xn��\<�1Z��i<P?����<�	�ҧϹ�=�=%[4�%X�<F8h�w�e�������;��N�B\M���`=��&= ��drw<�,�r^8=�慼O�üIǰ��y:�o<�He�m`���4�9��</�=y-&��%=6�=�0x��i=g�����J���gb��|[��b��\��22���o�dc����;�o�<^����}=80��(
��M<G8="��<_3�=�w��Ҝ;����!E=���� =�.�J�-<E.<:g�oƽ��fj���D�6<ۼY��<���<I���k9N=U��S�3<;G׼�!��?=?�k=P�_=�T��]E���ɼ�=ڂ���f�O�L=)8+�ʋ缰�=�S����-�[hB=~���"B�:�e;��o����;ZV �/�<��Լ�=+Q����<+���.�d=��a=,�
�3���(��'<��d<�P(�y��<[L=��Ku���2<��Ǽ%)>:Jb6=�#�E3��`�~�uy���<�#C<��#-F���L<@�����<=��Z=�Ԉ���<	􁺳�@=t�L=��,�~E����ռ0kM�v�=����M�=y}�����]e��y<��=Q�X���-=�y�<kq����ʽ����<$��<�7��?�����@p@���<ʺ/;/n9�-m�L@=;�3*<-�<0�Q�����qc2��.c=�=�<�ʼ,|�nǬ<���<y����=����
�H�������!�,��e�<�(:���)�%=�T�<vd��Z�6=�ͱ;ڛq;E�&<��R=��A����W�B���:�&����;�Z�<�^[�)��;S�g=�7v<���[<��Z=�fy��UX=�Ho���s��rQ<���;tO��=�G���<�eA=�z��%N =�:`=5*$=���<���;�re�)CL�f��`1�<�P����޼�K����C�����7�-�\��l�lX�<�>���Hr���;�5L����<7D=�WH�� =��ּng�:V��;#=S��O�=ꟽ�&m�<��<k���~��C�����(�<�2���7=�%p<*4�����<I͔<�l=(�A=�ZA=!M+�����Q��;ü0�/=���<Ў�<����-�^�Z=�I"��0�<GDS��&���e=����<���L�����u�˨;��.��3Y=�i�;MoA��(=���kJ�;ʹ(��� =< W=���;��]�	�=���<��<r�F<�Ra�ۗh=Cl=τP��3��a�D=fW�������l*=�u�=���;Z�<�O?="�=��n=x5I=��'<c�X��׉<�ig�s!=��ż��8b���O�I��j�z����<˯E�qTE�h�X=�&�O
�+�*=�lU��`.���f���<��"��w7<.��ͼRi���q<�4M�J J=
�[��=��Ǽ�v˼Q'@���
��c�.�<C� =w$E<젼_7Y�%ZF�޼���3t�)��<Nh���D6��J�s��<��1���I�S�;��f=eF��H��h�;��<�p�M���`=1�$<Z;=�!���c�%iy<J����U<�]V�6ID;ω�<�)J���@=v~=VD�9�&�<�=���<�g7�oVB=��R�<G�����9g�H�=�w<�o9�i�G=��<��#=�(��c���==6�����;�I�<j
��I<'��;��<8����Z��^z=�Z����<�I��,_��f����;l����3�v�^��ѵ<�L=�4��~f����;B)]�Ơ=�x����Y����;k)���n��1�<&𜼼�
�+�<�R＄��U	�B�R��<��q`��V<���j=��<���<j�5=�A =EK�<�?Ǽr<�Ǽ�S��x}�CPp<p��<��<����Pi=��<S�*��6�b�%:A�0=Nk� 	^���w�tU���|�?=d�3�[E�<~�(�������2?I��/V=��+=��;�c� =��c=y��o�;����L����6�<g���;ܢl=L�X=��Żv�X�~�==�r�;��/���;6�V���/�JWN=z	켏h���~�<)�<��<�Î;�����b<C�>�ei���`��?	�'�@���<���{\�<a�s��K���b���W=
���ol=�g=�H=�=@��<^���.�(=Gc��µ�<Gs���"�,�<}�J�	��<��b=v ��<_=�===�M�@m ��]ʼ"=b=]�+�<^r=�D��<o�5=��)��mz<YrC�<�'��g�<�?n�#՟<>W�<9�:;�F�m�P��=��Y=V�i=8�w;4���]�%=G栻/\����<�A�<�ļ<�D=��\��߼�ݗ��	<��;�;�}ϼx���9=)����d<�o[=r�Ӽ��Z<��=�Ȧ<�|a��_Ļ�]�\�:=����J�p=�#n=�oB��|�;�6�"Ƽ6����=/i3��Ď<9ԕ=�*=T�'<�@=O�3�/���`�����<6���M=3?,=gZ=/�u<Q�Ἃ?W��'3=\==a�=iSj=�`
<�?��뼄~�<ۣ��%����>��,U=�Y�<9�U=��D�pAz=�L�<�d7=&A=�р�d=E�F�-*<sF-<�$�$�Y����(<��<��I�D�H���<o<N= (�<I�R���<�=t�K=w'U=��=��+h��9=kAټ��<�r==X=#<Q�O����R��_e��T�s�<W5�<�l&<V�)�3U�=�Y�M�:��л�8w�u�=��~<��弚�D�����`�����-=�>0P=$:=I�9�EO��i,=�W!=�%R=r����B���=;⌻���A��|=k��<tֻ�S=�3P=��_��yZ�b�z<.�q=�=�.��;�1=����\=3N,=2x��%��;+�*�x��3������"����<D��<��=��� ��;Z��6�M<�~-�(�Q�n�r�9<�N[�I�#��%�:q�w���=؟-=��Z;"8�<!s$�AtD���g�X�==K2���,V��(�Z��<�.��W���F,=��O=W�t=,5=��Ȼ�i-�-2���V��0��ټB����Q=ǲ��#i=⠁<��C=2H��[�<�H���K=�nA�0�<���<���;���}����h�<Q�&��q:�S	��_ {<8�G�3�9=��Ǽ�~�<��>=�S�<n�T;�=���<,w���ļ����4<�����b����<F��<M�������j�<�;=v^�8��1��L<h��'{=�$9<LV�;`m.���*��V�wWK=�++<�9<�ҵ������$+=6ۼ�l����#R�<��h	1=E<L�sjg���9=��L�?�+=����q��V�n<O,2<TGI����;������=���YB=YD�ָ�`P�������)=N8��ъ�5��;���t-=�X��de�=fg�;�p=P0�L�6�.;��O�=����Mq�>�>��1.=�f�;R,�;f����`��2=!L��A��:��=��<M��<u�Ƽ�;�J/=�ݼ�(X<���; ��Q��y�%<���<�L���1�PP*="T�;�H��x�ռia��r��<=-�;'c�9ׇ<D8��8�X<����xF;����f=�P=�%�:�OJ��؇<�B5����?<t�̼�T[�l�[��z=��<=�;�/=wY¸�(�ސ}�E��<�h=�K��Q��<��μ�1�Y-D<O?=�"4�gN=K�M�H%g���μچ��ԏ
���t�uN�<|E�:��1=����Ғ�<��9�ʭ`��͢�<�wu=}����Z<�i༟�.���q��l��@���S]=����g=ͩ�;�i޼�p�N�&�x$=�����;�j<�	=Š���+�<�c=i�E��m0�U �;D�5�se�<u���a��<V��\���DN˻��H�9Dغz���e�0	��m=!���6q:���&Jo�.9���܃�<�V����=�ʧ<L:=��U�b=�B?=��; �������=߷�t�:=P�R�7�<��B=��<%�e�_�G=�#�<��=?�'=!t+=�&]=.�3 "���=��E<Y?(��=�`j��=5�x=���3�*�<C�=�ػ�G�;Ђ����-�}3{�F�d���=��<���<�l=��<Y�J<�@�<K-=3N��B8󼥊~��ׄ�����d��&=�o��a^]�����M��Nhd��<V3v=V����'k�� P=C�������,)�]�Y���T�t~=K0=(�<=�߼�K�+��=�9�=f�<�ޣ��T@�X�ռ��8��%ռ j+��'=�����]�������,��<���mY2��VλUTF=��Q�N���i='n�<���<34B=�:I=Ȭ=<�+�9���k� ��\ռ!$1=�ü@��������r�<���M�$��&�;�>�Lx;Kb��p�"�һ����S5=�_<$/'=��a�+��#eռ�Y=��^��r=j�2�PR�?*=�cZ�n�<���<$�ּ���� m=�#�t�$=`/J=w�*�!dD��2�	ĭ<��<l�'<������ۼ�[/���=d�@��$@=6s=��C<G˼�s:=G�M=�;�z>�xo	��7M��Q=2-��X<���@=��(=��o=�01�?�=��=+��<�M=l�w=>K=4n{�a��y�<z�ɼ�YB=4�B���N���]�| [=��a=y��<]!F���%<M�I=n2��H�X;�����;�I<=c�����?]�i�<D��<�I=

4����<�(�����#��f{��:=Ù=�bv���ڼ�y?=��μ�2���L��&��ռ�fY<�|�<�y�;(3R����<���;��<�h���H���=S.�3'2�0�%'�<'�;.E=9���`3=��ż�$i��Y=���<Wz<��m�;��|t=�5G=W7V����e�B�n,�<�h̻�Xm=/:"=��<O �<��[=j�S���B������y��1=Ҋ��<��<��=����4��*�Ʉ�_c
=��<I��<����I��<�=#�?;��6�s=:�a6��e����2o�[a)<�<���;�3�uе<��M��ml;i����:�U=2l�<�ж��A�<彈<a8�<d�J<��9L?Y�o��rF��7�ټ�2�=���<�A=s�]�^�|�=��&��<X"�<Z���z���I@�S��{`�Hn��9����9=�Oj<�~�='>=j3�� ��U��굼��;���<��;�L�4�)��8 :��<ȼ�<�ՠ�E')�.��<+QQ��oۼ�aB=���<�o�<M�1<	H�d�z���<�<[�S��H=6=U<�f�C<,	C�*u��2e;�=�+�Z�V=���<7=/�v<r�����=�%==6�.⼷����y)`��wF=�=I�<���OD$=h�|=Z�@�q���d0�Q|�
�n�����ɻY9�<`�7;GI<��%�Pk��H�`��F�Z=�D=j.�;κ0=x;��)��	���x�<X6�g과�/?=C���X�������<f��As=px�;��+=���(�<�ظ��<ܾ+<�i�<�������-k<�����/���S=�$޼�; =Y�伖��<�n<>��<�g򻫉�<��<���A*=�P��ՙ<�:+<>�<���;�Ca�� �<�0�!�Ǽ��<Ƨ�<cH=�G�\���H�0��[ZE=�мU�F=�,]�_�k<)C��5�xp�=����2{�?�=��N=�܌<m�<Os�;�n�:]M�<k<y���H�<`�k=��	��"�\��������-�M��4<	kM=���V[9��L=�Ra��2=![
��{3��Lg�a�<�=���:P�/��bǼ���=AS0�ڥ��lʺ�0�<i�Ƽ!3���M9=c߼<Ê,�:��H�"=���;(,#<gX����<��"���e��T2==�JH,<��@�M@�<qB$:ݮ���I���P�����"�~�=n�=W��< �1<�M�<�5z;��=��<gzk�.��;�3?����x����y*�eq�<�=����\y=o�S�t8���<�tW�gW�m�JF=���F�<Q��<<��<~[<��'�N+X��P�<?EM;���`h�<�@�<��p=҅I���!=�[x=�8=I�	�j�z��u�;RX�;aZ��D�<:���7��~�ռzK^�iF�<�<�1��)E=��=� �<��o=M�O=��_�=@��<B�(<��_��B��d$�Et�;B;�<US���»�[=�T��(��+ȼ�|N=A�=����*���
��ST����`�Ѽ�<�2;�3i=t�E��f�;^�@�]EL=�T\=Z'j=&J�<�,{��ŀ��k;=ev=^��<��;�
R;��
=ڥ�M?�����ٶ�<!7T�3�7<��Y����<��H=a5�����=�5�:ю��#�<1�<�=ģ����ۼ�^���v�<8	 =m�<�λQzm�|=(=y|X����x0=`��i7=���<���=�P�<n�=��=F��<�L=�NM��	k��/=��T�o	=�U����=XM7=�L���"=�Sx<.W�<��:��������<L(z���<��2<Y(����]^=�=R;�
�=�X����<�{B�M/v=�=�-
$=�o� <�� ��je�>B�m_�3��D�>=�<�E��(*�g�"�8�漹�p����<&����=� <��*=�
��м[��5�J=�m<��<n��� ��`�>�.�1�4F =&Շ�5�F<A��<5ǼBր�F<���c��6��U����K=F�<c�)�^!�:�~!;/�S=[r�0U-����=)��<��==Z�f<x:=�끺g'.<��U=��<z�A��Ѽ��ӡ<}��_�<���;o��
�ּvc=:١<E�a=�v�f>|=&�<��d=7<"=�a,�ܚ^=��_�����T��ZQ��4i=�:�<_�V<B2C��k�qoV��2=��7=7���H���b=��;�pj&���<?�(=_��`�9=��=���<���<	,��N��=hW�J��=km������aȝ�Msѻ!�+=�`4=�I9=���6c)<q;��:?�׼z뙻o`p=�8.<$�R�A_K�C����6�Ig���R=�PG=�*�<RH�>`�<A_	=ύ�<l��;�o���ڷ<�<=W/�]�<��L= Q�J."��L&���ܻ.7.���(=���=�L@=�`Z=ss�9���4=�C�S`�<�f?��u�8�uY<�;��6=�Z伪��xżl��dk=K��;�s��%���0�!�d=x�<�"V=�jU=t�h���9-l���f�=��p;Do�~���ϩ;��<�ܲ���=<��L=��=�Yu<|;�;h�</L�<��S�����H;d=��I=9�=꫉�S��<WE�<:2=$8�<��4=�E�<��P�I',�Y�Y<�A�<Bb��1�<�����0X��\,=�ZO=��0�<A��[4�%��%�=�B��|��8Y=�(="|?=��
��8;���o9=�<��U���S&�D�g=�*ܻ�<�<�9�w�����<�_=Ģ��>S�c̛���n=��j���(�\�W=��\<�W��R�km��ȧ=���<^��<����B���޼���;��E���<�"缡B��:�<��v�:Q=$�=�V��k��<���<��;d�O����=��<%���;
�I<<�2= bO���"��I=����S���<9g9<����_�M���l\=���<���K{���<JJѼ�R�Gqa<�FH����$��D�M̺��?�f�r�� ��HI��}�=}[z��fY<�i;��`��-=�d���<�5�;&�;010=�Һ
��<E`=@i>��$Z=��<3�=�c�<��7=�5X=����,���y<�˒;�\����w=mj:��<�;;^��S'��{<�ܪ:)B=P���/�����מ<=9�ȼU0��F��Y���<�)=��a=ч�;���<�ۼT���C��<��^���I�fS<�<�W�����O�_=���<����t =��<؆8�{�:��W�sv��i59���¼c��;ڛ�h���sA��2Q<�cG;g�6:�~���7=�=�h��G�i��+�~=X�ļC�l��O�	=��<��缄�H�5R=$5<�Um��?G���<��6=���=s���M���,�3f�E�r�>�Z=�g�<�Oo����<�G=u%-=�CM=z�廊{�;��{�P����;=, =S���j�<�Q�&��<��<*ң�O	��x�Tp9=&�<�x<�� �<q�<<v�;<
hP<�a�<�(�K�z����<�:5��B�Z�����::\b<@�һiYN=��=��S=&�J={;�����e�3�G�}�=���*˽<'ᏻ�!�<�[@=��-�c�g=����2��ݼ�i	=`�
=QCn;�=�sp;3<�5�����<���<��r<Lyw�?�����<�0W=k�<8�=Y|�<]�E=��A%�Y�6=̓0<6�g���<}���4�;��W<0H�<ӫU�:�5�:�<RV�<EN}�l��2��D6(=�����;��E��8��<>D�<�&�<AV=IɊ���U=t O�2�=jI�?�8=A(��ywa��eC���<�>�'�輴K�����0�8�h�;_��;S =ַ"��I<�����;�)=�SR<j��<n�!�᫑<�	q���b=�i��Oq�H�a�-/ͼ6qU=w6~=pD�<_��<u�T�A{��� �;�"���޼)v�}|=5f��y�!=z =�R@=zO�����`.���Y='U���!�<@�ߥT��=��Ƹ+�����(�<EU =n=�Ǽ腴�3`_�ζͼ�<���<�Z<T���5��<�`�8F��y�<-���>��<�&E=�����O�}�Ƽ9 =ߔ�<5S<;=�8�^ɱ:�!<09;`�=�u�<�["���q=u�<��U<"��;�;;=߀i���X�4!�T�]=v< ������{��kt��P�����e���d���pu�}��<S�'�:L�:�ia1�@q�<ْ`=�!�%p�XFZ��5�<v�i=s�b�&Y����P=>P-�ծ=�w9��D޼���wl3�}H �9NѼ��'�=���<��\=�fR<�	E= ��Cp��׭�\�<��^=2�e�H�ż^l�FQ�<m�$=������G�<���lF�<� ����=�<�$o<�B=�fR��?��u��p�g=d�<��1=.��:�Ra�1������<
ȼᏓ��t��2��@=��p<D��!��� ��y;.=�����'m�;-�[=d���)⼨�G<Bo�����<{�8����<��V=V�8=��ѫV�r`3��I�=��Z�& �Lm=/�=m%���=��,���>=��}�H=_=#;_=��H=^���y�<�z:�ٜ�<9�=�`F=��"�p:#<S��q�����r<.�p=d<�#99^&=YoD��߱:=m�<�,�<�}��m<�Y=���S<ݶ��m#=Z4=�I|<v�ѼYl"����b����G=��<��*���r�����ˢG��r1�5ۅ;~���N����=�J5��S�<BTպ$</"y=/�9��ɥ<cR�<M�<I�]�,�;��<��6/ =y͏:SL<=N�5��;���<4$�;� =��=��;��W� (h;d�w��2?��}Ƽ�V;<���<t��Wy=#'0=��;���<�~�c�0��5�<�	j=\PW<�6�c7�^Η<���6|?���=J�L=���<�,8=��y<��^=��E���=��ݻoIi=��8=Y7�]��<`��9�\<cR�v1=�`�<[�=t�3�._+��p`�zlt�b�<��<I�<2�����==�c������v$=��8��G.=��;G���.��ϰ�^k4=ƒ)��s��/?����*y��vWμI(&�mp��1���m9�g=!��<-�.�W����4=�C/=j��"=o�4���ߺ��D�H���Z��<H�a1<,'=�!=(:<�̇<}�<.J���=�.�ڼS�0�E�n=��<�49�������<&f=��}q��%�a���<�ټnq5�&]!=�W=�2�8��<+�ټ�;�<��H=�6�<%\����_=2��7(S=^��]Ni�LM���N�Kl��ف"<�:�<��3=�-k�$��<,�+=��>��ψ<��=�6={����w=�lӼl=[=��;�r=}�7���J=a=��;�s�.;����H=�(?�g����_�z��wg8:��F=�=U=�?1=h����\�<O&�&�f��Cw<�˼�����F�wPm���Լy߼�J�����ݼQ�i��1<,(E��=�<��<*Լ�'2�g�W<y�i�W����
=��=��<�7=>IX��/=k�,��/ļ����������O-���7=���`�<p�㻬-��6���B'V=>O]���#��t�<�N=&�<��c����;{7�<�3 ���)I�&�V=��+=Re=�w���r��'=�˼��<�4�<U�=*�b��������ރ;6�>��(=����e��M��d�w,=���<��	�BU��]��`=���+����?���G=�H�<�$
���p<�<��;�����<H�	=�%S=���<���|��< �G�O-<�w:=��-=e�;:��;G��3�f=��'<Yy�:����*��B�%=�w{=����<'I=8�<�祼J�I���ۼF�(���Ｃ�Nd��~v?=E�{<�i��s|</O�A�<�@=<壼�-u�I�<�д�c(�<��A��M���V����<P]w��W�<�f=M�&�1=�S��\���a���M�<i�=C�;<<��<]�8=_�]����qL��j�?�C�軓Gh<0#�:��c�<�o�L4=�w7���<˙���n=C��<��<�D=lf�2�7=�h�<��=��:�j=o�h�<�y�э�<�H���|c=�6=�g�<�=5=��R���\=< [=����  k���F=�=��m�Q=\i=�̻�)=�i�:l�X<Y�»����H��2�t�"�~�r'��"6�2낼
���~b�;��D�jڟ� <v�_�;imF���(���=3 !=y=TT <f μ�V#�K�O�T<�W=�l�!,=��_<�#<��<���	��Zk�����&�<a0=�����9C� �=���3�$��w%O���=s��d*�� m�<7�h��I�s�=VN#=��W<reJ���O=\�5������m=��;$�	=9N=֒�;�WV�����h.����;�y=RA����O�<mר����<�[=�m�<3=�n��o�<�3����;�;���߷�||G;!�O�3�"���)�C�=e��EDY=ȩ�R<�[���h= I�<�}>=c�6=�f�<��0��;�B]=K���}���=W�˼!��<�xQ���=&P^=;"=������<���<�B=�jü���h�<��<Y'X=t�C=6�O��<�X=�����|D=���W���<�o?��HZ�ʟ<�A=+�'=�E3<�s=�0<�EU�Lv[=ѳ��� x���I�Z�<R�E=p9�<�̻߁��xz��X�<�s�G$�����;�o�;B�#=,��<J'��W�<��g<��<h�?��1<�=��c.=��#�6=nN(��O<˨�<-�*���v=c=��@�_b9���<ґO=l�r��2v=t�=Hm�k�6�1����.=7Z�<~}=.%*�^�<���BNy�ExG=��T��rM;4�便<�&r=�t�=�2�����<�����;�1�ۻ7<��$c�z�; ���P=V*$�V�+<�Td=�N���I�W=e�r<t�y=�M?=��E���Y���<w�0��h�m߼;���n�;c�W=��H<V��<��=��B;�n�;�V=���&o=������<�����d<��7��6�=6X�g�	�~�F�^4�9t<��=�i���=���=�(=��a�'` ����<�%����FkҼ)�T<�g/�������&�0=��<c�7=?� �ӵ�<���@pG=ba=��\V���(�EN�<��u<v�u��-�;��<84=�KO=+#q=ch=� =ـ��	\=�6����[=fa=V���<0�3��d�<��'<����MU=Ou�<���<8��;�c����ռ��<�B=B).��1/<�=�n2<Oly�r�<�	;&���>��?�d<���<���3�0=s�M=nw6=�HG��I|�l��������=��J<;��<I�>=��.�E)����_�]=_���xG=���a����d�r<��<�KA=�.ܼ'N��uթ<����Nn[�q.������[vy;9�y<A=��
=�E=�=�ߍf�L�7=70�Y�W���Z�	��H�b=�s�<#��)d=�ƺ8[G=� ���,=mԊ��
�Q�(�6ZF�$�=� �
ڼK!��#|���O��U �K�5=TY=f]0=�>@�a=��==,����?0��r�g,�<r��<��E��qC=��v����x<�0A��b=7�_=(�/�<�=&pZ=Ř�<��; <f���6i�9��;�L��q�:�X���eؙ;�S�����	o�����@<G#<��=����<n̠���<Y�<M�=67@=`�8���&=�ٻ���T=c�<3끹�>Y~���!��c��9="�ċ=��T;�R�� =��������M�h��<~�G����<�-Z�AI=�tB���R<��C=�<��,=��0�<1�<갫<a!b�ЯO<��"=e��=az˼5=�;3/,����=)d�צϼ��<������;��T��\,=5��;$��<�d��&�d�p_�����;(m��甔�g��A;{켊ϩ��~�Ћ;��]ƻO@,=t�L=�S���<.V!�P�?��4���(=I<��b��*x<F�R=���;��8�dR6�Hh�b��<r>:�{(&=�4����g�o�;��>=�'X=�jV=�V=��%��|�� <�#h=��ȼR��<d�C��]7<�(<=����v�9��<���<y��<+a�</#^=�:$=����I=%*=�=�M<C���+�t=�4�9�O=������*=g�z���;9����>�X
��8�֍C=��=_�A���_=k>=�<�~ʼ�cq�b6=�	���?�f���=�b=9q�<���<%͊�m�'=��=�����?=�!K�C��p���TH��#t=�6�zWb��!��k1=�y���=M!!=1 =�X�:V	���m=H� �Sx�@{ =�L=7O=�ư�B=�D	��/8=�=ϼ-��b�K�%4���U��P6�O�R��R��3����<hO��P��<\�=���:H�	���|�$��� f�<���n�G=��=���Q���n�����;�(�(0B=��b;$;��<�/p�{P���s�<�<!��*p=Q�v��+h=�N�n�*<6T"��/�<;�:���;���A?����w��(�r�G=�� =�sQ=��9��� RI=C|Q�c༫�����Ʒ�<��=8�<��U�<o�׻DL =�'���'=
X*�h����=�) =��:�l�ī]�v.����Y=�<f@=(�*�W���2��jE=�p��=.R���;�b|���!=��&��<!=UEp�V�W��;��Q�<�d�ֳ^��Z;��=�54��:�i��EX�%��{�=;�/=+?�=�X\=.�O<޼НǼR�=�#'i<<�����7"U:�'X�e�5������y�;�:�`�8�e�-;�t󻎱�<�xb=�gt�n����Dh=T�ͻソ��nPP=Y�K=��>��U=�׻��"�j�6���r���%=}V�<T
�A����{����k�j�J<�1�;��-�����Ƿ�����A<��=�F}� �_�u5=����o��}=��N�خ=; �%=���w.;9=U2��߇c�Z 7�o���֎U��>��@��<O���8T<��(��x|=���<R�*�xF��{n)=nA=W�;|^a�	�n=�B��b��EY=h��
�ȼ�c/��&Ǽ����4"��K����N�P����e=þ'=�k�<�d��sv@�P��;mx;=��r<��,;%�0�H~��\�Q�X=��"���u��v���l=.���ŀx�P�=Zs���QJ<4$L=`�˼ot��l���.��ٰ�I뫼�'�z��<���������<c?=�u�<��g�OՈ�a�9=ك��ѻv���<ݫ~���:�f=���<�(z��:=��	��C]��{�<��Q���ļ��d�w��<"�)���eQ=�Ԕ<Ԝ�=& )�Vl'��DC��'��@#=[0L=��d�f˒;
J��rX��X[��!=�V���b=i���޼��'��o���Ve��{��V=��t���h�[=.��<Ӱ0=�)����;�3=�xw�����.��i���y/�n�Z<uA��x�:9?$�|��W�=FF�-�b<�����<h����nl=�7=�y6=6/�<7A�;�ܼ��<ȉ;�v=��O=)�O�m�D=�{��RE�Ҟ><�Ã;��D���{<)+�c�<��M<gXu���=V��<�*�<,�<��+���¼0+����f�D=V��:��U=I7=�� =����o=��
����,_|�Aց���<�� ���=(?���<�o=�\<��R�6�s=tγ<�Qr;��F<F�l<r(���=kL��.>=Q� =������ 1��h=��;&0=d}�H=嬧<<Ɏ���6��j�<��p�U�$�^E!=���6�;�j�toU�|�=�
�;L� �!��7�<c
�m�<o�����'��츻d{!=�<y�ټIO��Ű)<�3�͹<����M��*=��żY�=;Yx<����<��L�T�,��'���3=��a<�`=���<i��<�ޠ��J��|Z.�EYH���7=k�*�U�gkn�߮��m�<5[<��v<Y�	<G�ϼF	���O��n*��K�X��<��X<��<'�2=���<k��Ji=���<q�<�%����<��=�h�USy<#�b���;���<,�=�	~=LR;�!ѹ7v=���=�֊< �l;a�u�h��<qfN=�HB=�G�4��<�SQ�{5*=5�r<�e����/�\b��'4=M�b�n�S��Tx=Xu�:��(=��5=�ҷ<�gv�ˍ;���<5�E�G��<�
)<=GF=*@�H�W�_��͇���[��m�<�D#���W<~O/=�bJ=�"�����8�*���:�\(�=Q��!,=�<��N=i'+<��.��)=վ�;6��`|A�x��7|tɻT�z�(��<��ż$[7�ާ�}Q�u�<�䩼.�ļ&BY=o�>��f<�Sc�i���;��8���p:=C�9=��6����La=��E���6;T�S<]�R��z$<����="
=�{���0=�O9��ۻ��D=�Ҧ�E�=I \��o�<�?=��B=���;s�>=�齼�g�<���;�7y=ܳ��(�<o;	=�*�<�v%���l�`�伣%s�2&��q�⻪e�f;��;��|'�<�\^���U=��6=�a=fr<��m���;�q�=$M=� �<P�:��`=B7g�����ڈ<|���x<��<Y�=%�l;��<��E��F<E"�N���l[��n����=?�M���,��0Ժ�aռZ�������Q���򼲣!=���F�0�Q�;A!`=��=E���4����<�ES=jv�ৡ=TM=�����}���^'<XgK=�7J��P�X���n�;4���p2]=놾<,�A=�������<YH��p�"=/�7��逽*u+=�Ne��7b=3��<u�bG�<�����X�=���<d�<;t��<������e��<-�2���'���P=W��<��<��u��`(=޻�AUa=�>=��H=D��<�&ͼ�S<2f!���H< &<��ֻ_EF=�l�<?ɦ<�t弔���$�<�*�!�ʻ��3�4�$<<9���,N�/{[�㛩<r<`:J�v=ކ�������P<�2=\�2=����m=�Oo��n���P�;iK=�ޜ���1=�UE:�;����Wv�<��׼vÕ� ���N�<%Y��|����<&�j<��$<rp�;:Ǭ:��-=+Tc�6e=sC�:���I�/��&j���;�8<!����P�ρu��p�;4�=B��4<�Ѷ��4\=sR���/=�M��ļ��3�=�X�v�=T)=ր%�tF<m�=4
��=�~=���p�;<2�b��u<�&;�&�;;21���J=�������<��_�lӻ��.�Y��:���&�F=&�;��<=��Ā3�!������W� =��K=�i`��т�5�<�hL=�~^<�%�;�\���h���)�]�:<�A㼋�-�R��<�=��l=^�<O�_o<��-�f�lVb=4��(��;1�[�$.���t��V�<�=�;��ּ�Ņ<�@��H,=f�5:0<������u�<=�D�0.��x�l=��J=� i=w'�<8�="'U�fN�<vI��ʫ<!°<8�g�="\�< &�<U)��Ϟ<ʽ�<.���	Ӽ+v�;�k�<�K��NP<�7���vh��$����<=����`=�XM<V�<A��<=�?<y`t=O�\�@7�<��-=��<=0�C=A&<=�e��#|ɼ!Ѽ�
�;�r�:��޼A�����ؼ���<ҷ�9����;_4X<Aa�<osh<Ȯ�;;e;��=�<�<�ݹ��*�ܻ0Rt=�@s�J�Լ��3=��R�!�=1�9�{��<�K�iG�<�8�:�U=��+=�6<�G;*��<U�<:@~��R���+7=]	5�+QU���P�����p�<�sY;��:��9���<��,������18;ݓ�<JJ@�P"=M�9=�3<?���u�<$�W=��m�r0!=�,X<�\����	��b<4kn=Kl	�VP�<�5��aX�.y�|�/=�v�<��<G�����-��=ÑA=���:�3���Μ;�7v�S��;'fp�1�I<��y=�<����D��h���/=Tv�=+�L�[/M<��-��[=�=�d��1}=�Տ;�/=�@��E\=,�>��yI=Q�A��<Y\�<�^��\�<o=���pg<���<���:;��< ��<~����o<�;�?Z<Q�;H<�8�<�9T�9M��&ּ�w=��=^��<I� <����<+�OKX=�"�;r�����߼��<�'=�&߼ɥ�=����|�����G�F{�<״Ի��;��4=bc��6�<�)=^d����<: ���1j=)_�;j�:�Eq�}0)�yK�_�]�ϙ�T�	�l��;��<��.<kd,=}�=Gۻa�M��º�� �M"	=��s;��!<�=m��<i�;=u�k=�μ����d��� �%Hu=����GO=^�<1����.<=D2�U��r�&��`<[�e��Cټ��6�A����=����3��|�;z��C�<��:=��ĕ=c>r�شe�.�=�.7�.D#=��/�_§;3�U��.�$ {=IN�;�oZ��f����W�#$�a|���]�����5O�͸�r=J�Ou <�D$�@ �d�&=��N=t_>=�S=h�l<}9*=�~;�u8�y��<���:�����N��m��s���w=UB�:�bN������ϼ}�.<g|~���W��b�Qs�#�<ʻ>�떙<'/+�}u�=��<��M�9ܺ�L��[�7=��ܼu ����ߚ;=?�����޼�#d���<����J���n;=j�<l=�:�:ܻ�<x���ŏ�O�:=��<U��<�B��F�<��; )=t{<��`<���<��~��^4=��d�w�;=� =_�Z=�桼d-�<�=�+Y=j'��mMi�*�<+T�<#U�����B�r<�*�<U�e<r9��!D�l�m=,,������;������D���<���V�W�(������?K��(=P}	=<I���'�(M�o=�:�8<l"=N��1���)4"��[ļ=�<sq���I� �x�`�EyG=0��˶����V=�TZ=���<ic��0��>g<��ռ�D7=��c��-���<��6<�A�<-�L��W���ͼ`i�<
�<��;�}��C$Ҽߚ����F���_<\�x���9=H�/=:���9���xJ�[�q��<�W���!2=�&��Y���� ��k8˼���<��G=�%:=YYv���<&�6=/(=�PK�yy��K�;����.�9�y�\ؓ<�P=�=3� =��_<�)�<�
=�{/=B4V�z�O��LI�|�=���<�U=��<�q��ܟ�:�	=���<��D;=M��=<��EM=�+��1�0�<5����ļMW���,=��A�W7�<�҂�i�`=�9=My�,l=�kU<���<?�i;x!X��0���<��4=�GS<��;\'�<L�<�8�<-&��Z���D<�'����j�J-=h�2�J�=����)�2=�@�<�W=ܑ���f7��J��L.�®�<a�[���-=y�=�����8=M[�<1�=��$�F��<�̓���C��
:�h�G=�_o<�u�%JM����b���h<;�K=�%��j��$5�<'��y�S��=88b��-����="���n��]�˦��F��$�<?r=�9��Jջ��G��@�*�	=ݣ�<SQ�<�м�xBh��a/=�6=��<x^�<��<��#=K�7=��=x��O�x�D<4=��4=F;�͓	=^5ټ��i=� ��6K��q�7�ٝP<eko��Y�<U��<"��;P�a=o�+=Ye����<�*����&�e��7</��<|��<��S=�/=cH ��vE=�=���x��<� ;R�#;��Ⱥ$s!<o��<%$=P:������o��$�v��8C�3�+<g}'<"���*a�Ml7���9=���<�Mi<�=�}��-P/����<�Ɨ<K��9��z�KZ�������;�_ܻ8�;�B�4;&:����x�W�t��_��;㺤���6=��=�9�<�8b=o�l;�m����Z=sN=��	����<	������<w��;�N=��0��4���)=�����{>���=�֞;r���F��P� z�
B\�s�@=�i5�B��<w42=>�=�{Z��Q���y��;=~�|=��(��,-�M�d_k�r�D�I�����c�� �=X��=�-�sO�qT�=lCI=z��ԙ��.�6��[���=�F�<?=U�1���g�/��R�L�H�f�,d�<��9=ӱ<U�=�E�<�V
=��ʻ��	�e==s:x��X��<�?=�l�;�DG���"i�<;��ܙ��S�;"�I=@�t<*�-=��@A�;�]���ȼid�<s�����J<�mZ��=�4��-�0��<h�|�;x)<8�;��c=�b6=,�T=k~߹ � ���%=�Z�;(��<�L���=|U<�yu����<'��;J񟻟��u"|:��=�V���"=��'�<u]޼�1(<��	8������M�6�ͻ׼�<ťh=Sm�G��;�˓<R������Sc=�ڼ�a��1� �|�:}�P=����P�����<h�@�@�Ҭ��k<m�u=T>�d�e���&�`n"=wg;xܙ�Dcݼ����|���:<�y=Gϯ<1�3;�����ԕ�ƒJ�ŚP��e�<qL)�"�.=AY=�yC���=m�q<��<l#={��<����`=�F��3_E=0�<�M��J0e=]�l��mJ<�t�&ۏ��V=B�ּ�r�:��T=խ�;�*<G���==���<�(=h�KL;=c�
�j���U��w�-= ��<��<�k=#�=�z��b.=���+޻鿳<@�;=
�:=8m��P~<!�ѻ�� =��(�%A����`�0��;����� �%�.=����k饼��'�6肼lR�N�
�@��<��<�C�5T2=t�������V=��R<e�@=
L�5�;m	���L�<�}�b|���(��R=�!W����<P��e�I�����{�X�r=�@����=�8Ｊ��;\�^=��I=߅���2"=�%�<�X�� f��'@<�2���<��X1��啼��Y<����@����=�=?=���� ,=>Aq=1�="��ꑼ��м��M��oS=����}=�����h�����<� �<#�<6��<�(`���Ѽ G�;����S);�]�<�+4���J=����<<�u���s=��G=�g��il=`�����<�7��W+��J8�,�j��ߘ<+�����:�=�-!=}f��䪻�c=٩�<���;��o:#|:��+0=�.��tX���p���g�\�<4ĺ-ZZ��q��'��t6=� =Q����"��4�:�f����Nc��4�"���z�B*=�6߼��׼(ʼ�P�<Sl"��~@��l=��u����<,����	3��2����N���و��
<i��N=A��<��r:#�=�S<z�`<yo%<�ڋ��<�t*=v;��g�=έ=��=KZk�D����<1?l����Km�z5�_$=�{=���;�]J=�c���E��m�_�;8i��g�;���_�B=5�=�c=S�[<�(=Ū�<��C9�I��!P�<?!=WD	��V�<�ػ�G��;̨���G=�S���$��m�=�bq�MC=�8A�u�=���<ǬD��a1�dY�4��;P�R�H&=�WP=���<~�C=Q|�=_޺<�I�;�\p;ݙ*��==����Z!=�O��錯:�2#<�[���=��$=�E�<�%u=�1�<�T��^�OL=_�3%�<JgQ<�y�=���.�H�Ca=�v�Bg+=,�����=�ez<��=��=�'�:٨ =k,ͼ#�U=�TǼ���<<�ۻ�
�<��m=+�P��f=~!=0�q�7e�<C�#���q;��	=ܣ�<���<,\J=��o����*:9=}I�<m�U�I	%��$���\��M�<��k���1�k��Ls<���<c�$=i0 =�|<���<�.��2��}=B=��r�J��;����f!&=�UP=�w���Y�D|���A�ug=Y	=�@T�@�s=��̺Y��<'2���I ���̺�B�"�;�������Rb=<��nJL�Oһ:�^=B�p=8��;��Q<�*;<��2<�4=(�&�J��'�Ҽ�/=�x=K�m����qZm<M�c�w*�<�m_<���$;�=3��S;�����)��� �yZ,=����r<=�j-�8�� �%w�<	�<�O���?(=�m�<5eI=%5/=W��=�#�"{�����<���;Pz�;V�7=J-����Z��j��7<�L�2o�:׃=��*��US��C��C�sLF;�I�=sg�:01�<�=8�@�<���:�.����<��㼠��EC��Z`���	�3�3=x�+��PM<�	<5�[<V��<C�cϾ<U)�����ۛ���=\��� �;�=��@�����S=r��eQ��_�-I<��S=�o�<��_;|3�>-.��у<��=�k���<�#=;?l=�2-�7=��QM=��T=�[3=&=�^?=t�<�ټ�05���ɻ������<4�<G���i@$�R弄�b=�Ĭ�_�	<v���]��<nv<s�ƻ�ߒ�[t�<�/t����<]���g=��'������|�Q��<A-６�=P��V�2=)�K��4<�]I��d�������<�=�<�E�����L�<�{=n�!�]< �x�8佻����o���%=��r��
#��s�_TK�Qf;+�M=u�&=�D9�������'*h��c�< � �?� �H�F=��=?�a�-�a�Q<���Hv=�~<���<^a=�ET=�����������?1t���R�}�ft;�*���E<��<6��7�
�e�K�d/>=�w=�<�;�){���_,�dB���S=�K�<Q�<Iw�đk=]�I=r;=�P���<��@x��k��<&��f}�)��<��K=�_��cJ=��켺Ȼ�C��8��<R�<��8���I=A@�·�<z@9=A'ܼ0�V=�<=5�<���<�&=��<<��<譳<�t.���D=��[�D�^��l��Dмީ;h�b��"��e@=٩�7��*�1=�^9�aaX�L�F��z?=��W=�c@=�^:<ܜY=`<�[�T�=��	��?j����з=XH�U����9�G2=c?�]¼ļs��ͼXF�x;��I����[[��9�Z��=��P=<�޺]�6=��nn���>�#���A�����>g�<��U���D�C�U��L�;��S='
�}��;Lf(<�D�<��ƼG�G;��W�B�v�Ւ=#V=wE<�V�+�<%�I��;�`
	��� <���<�������[:�G(�}���l]�3d=�@=`�\���'=7��<E��:o�S��b��t�<	�=4p�=�^U<� 
�V�u<�4N��ht<9�);�+=ޥ�;I�<wNͼ31=�\=��|���'<�9-<��B�ɥ��/Z�=�W=U�����<���.E-�h��<�J3���̼}�$=��<<<eJ<�����4����Y�~� =��<��<n���n$�;.�X�Z	:==�|��`�<:�G��8.=C!���#%�H�����;f(=��:;DSN=%����.����^_)�
�?��6#=� $=��c=�C`=Q�V=&���������=��Z=�����<��=�J����<Sa[��-W<��=�͑9��؊<?��:c�
��7����?��հ<�^���=4��<�()<p�`��f������Φ<��9د=;֪<�C<E =�y�=�!�����<2mü<RB=�;&33;�m��}�S��/�E�x��L��p�q䃽�5=���<:ԃ<�H=�.����;lK��e�
=�
��[�� X=�$��i���޼�O+��h<�rA=˶=��ú��/<�����ʖ=G��<��˼�,ʼ��Fṩ��y�<	�b	:��¼��=��$=�Ӽ�n�<2�����T�Mx�<�
-=	Ć�`������;aK=\�<�a����� ׼=�u���<��<p�����9
	�������/�<�
�0Ǆ=6N=j�~��c�
鏼��=�=�m&��1O=5��o�];�u�<Y�:����;�=�-��{)<���;�ͼb3��U�<0���=k�׼Ms�<H���=:��V"�$s#=V]"<���<Y��k-<}�=go�����f�T<Βּ��ݼ�;:J�9����B��2�V����L=�[��\^<jO=�����03�e{��l<��Ƽ��<�d=�vs=^T��*�J<��
�<���;�*�<��:�6A��ļ�	�<�{�gC�<G�&�?��T(�MߺE:����9����<d`<���<w~,��?뼑�j9;���<@'=x
E��d�;��$<$/<�0����|�[e��ʼ�*$==�/��@��G���`��&=�*=v��<-�<m�<�]A�~%�������$=Xg�� �<�J%�)� ��I�L�<ΐ�bW���7�<�P�;a|<��H=�@�<}��xW=Az=�[���^=��(=�8h=��⼽勼$��3Is�lB; a����,]
=��%<���=��N���ڠ�N8�e�w=ߕ�|H��q��
���x����P��.�<F���MH��	9����<��?���=\$0�C�d=x.\�&�E���<[I<U"<�U.�vu����<b2�1W��@<�3=���<b ����d-��;E== 	b=�[;�FNO�.�>��1��@<�"ʼ�i?= w�$�%�g�%�8��;�q�<��ϼ��ü�Q��@��(#=���;�"���2�,�^�	�=�%���!�;�=�F�<"=mY=�v	=�Pc=���<'Q���#4��f��G������<�'�w�#��B=��f<�<�
��AF��C��Np��{?�y.\���%����<���<!�&<C<��KQJ�3�P�+�2�����<q��;T�<�H�<��E=��5����	c=vἧU���?-=[>��惽��1=9:���� E=�$���k=NC(�R�=�О���J=��<?&}�(@4���"���E���[�=Ӌ2��������:��X<."���*��-�8:�S�<�6V<�a켠[�-�i���N:���<8��<�:�=��!�@EW�l8�<�I�<�� =�Z+�!��<���:�B =��/<�8��̛-��I��}��N=y�;���Ҽ*#x=�3I;��*9�aA��A�rX<=W���
���=7{=5�%=�?��.�w=�bļ��
�hy=�� ��F<p��<���<�2]���D��m=뵡<��<	��k�<Nc=����T[�<;l��D=<���=
6M�!��9c=^=V!)�����ҟ:K&�)�=y�=	�$<��#=Cyi=�uM=:�5��<��Njr=uF�d�7��m=ډ<��b»��e=AzQ��� ���I=�HG���N��XN�{T<���n=FxW<�C=���tS��J��<T9'<�$=+=@=��Ȼ�<��<��q���H=mk<֟M;��"=Dxq=��w=\_���=?����R�x�5ռ3v)=��=.�O7=l��<�ټ;�<�"��E�q��u)��ߒ��b�<�h�<9�O�PZ���<�ݧ��8�f��>VǼ_i�<��G=�yZ=��6<�2�<_�=�|���^<-ju;\X�<[��<:ܜ���ż�<8�3�LV�����<�P�a�<^�=�C��QUd��;�=�"E���@=�e����v��o�wL<sul<:	;=����r�>=�xR=A]���'���� ������1�J�$��:H�ݼ%�N� �v=�0<��<�R���	i=k4��ʃ켩��;�/���^�J�s6��S1��=�\���e�N<8@F���<��N<�*t����0�=�W�g"�<�R<,�<L˰���=f��:I=�$Z=�xԼ
�<�b�<�9𻭺j�2�O<�����<�6���I=#��<�<���;�$�;���<	r�<�ip<�<�ɺ<?�<�N=�).��f
=�bW<��<b�A=��n=ta<�u�<1
��	=�2=�j)��!~�x*=�.���F��%�<�V�\�M�u{P��I�<�E�:8zϻn6��T-�޽r<����e=��W���W=o?=A�=Oa��U���s�?*��-=n��<m�p��%�<D���/�тD=W��<[�L�NJ.�G���q��8O���i����<�7��g=Iž���<ݺ��9IV=�2��֌�<�'J=�R%������<�fI<�,=�]��ܼ�b<��0����<�ZI<ש����Ҽ��
=Hg-<?s�;�S=Ҁ�<%4=��f���>=u�=�]�
�p��=�f��G=�.���?%=Ay;�S=��|�G=����ty<�5�<@=�i%��%<y�C��8=�g����R�C<���#!�<��ڳ�;��l=�fW��a_�?B��1�;�$��>16=Ք|<D5<��J��Ỽҁ�<�D>==]=��=N��<� �O���x=>�<7_����
=���<���M��,�=�ͺ��;�B����<ɠ5=�^G�3�<�p��05���j?�L"�AA�)ǣ�L_�oN=��&<Iq����>�LB�tQ¼�-`<�}�h�.=����R�J�!�.=�*B��Ӽ�A,�:�]=T�f<��<�o��ce:=��<S����L%<�b;[b�<���;�Y��"����=j���ȴ'��j��PH=�71<��(��K���U=��=b$�<,�|<W(=lGU�NШ<��;$�=�aT�F�<}x�=`G=R0f=�;�D�(&�>��;1���Oq=Q =	�X�ޛ?���*�:`�;��<��=b�j��᰻X� =_<=/ؼ��*=Q��E=�����5�B<��;RL;5,�<\@�<#���h9�s-�H���}=�ں��)���R�̀
=C����๤��#�<Z܊���z����<��:��T�1z伉ņ����}!=k�J��G�$�G�ϨQ=J�=�>�4�M�B<�>=\�h<�������߼�+2:ɕd�S�<T�<lB=!�¼�&G=���<���<��1�s�y=�vC�w8=�YL����:�-1�2z=&�<.���󼯉�:HE�<�?<CuZ��<�1b�3�&��-�<�#a��<�����Q�<V�����E=�$=B� ���#<��A�[I=��<c��;���X�?�~��<npѼ��.���<6jo��w��V�<�ɦ��w�"��=THE��~V�;G=H�һ§R=�k)=9}W=���tѼ�t�<�7=�q=�[��n|<M!¼ĕ%�N<��JmK<[<;=��<���֞����p��ʣ�y�|�;�q<�`l�Э�<Fi�0�YV�<�uݼd�`=\��K=e�Y=����<%��Ĵ;St�=yji=Ȇ=E1����q#�<��<�^=��<��;6A=�He=�����?�Y�|�-D��?�=�j��8���7����:��<��b�qQ�U���J=�jh��b�پ�.�:��j<�?�<�"�:icE=�����;��_��gQ���O=���<��r=�S{=��#��v<n���_H=�Y=72�<f�P=��s<e� �j��=N���9=�!<����<:K���F��"�<%*=#�4<��S��[���y�1 =݃
=��ĺ(�
<��< �+=��b<ET�я�<��Q=@�X=s(�U�5=�n��x�ʼ�;�x����2=nWS<�-)=$����<#[ =���|�;Am�<\;��(=�x��Z<B��<4�ۻn��<.=d����:��I<�6�<u6v=���wߣ��-;�.��s�M��g=��[��[��a��*�a;��z��5��� ��I�jn��;dZ;�k��)���G�<+1�aw��N=�j%�_��;o�<�T=N;P�{B�= Z-��N�<-'=i�f������b=�t �W㿼|��&�=�F]�.����|�>=�	�9�G=���<� �բǼq��{�;:7o&<;I�<�P =�\;
S�<h�=��F=s{�A���=uy>�((H�;ky��Ӽ�ؔ<h�6��s=�u����:�*)������<gk���G=�/�d#-��;d�� �B=�@����B��\�<�;�<u}�ص���M�<���<��T;�S:U�A��=�%��Q=�YL�3^Z��x�<�=�z��t8=״��Z�G���:���|�o��<1�<�V�;?���K�<jxW���,=!PZ=��*�
Ҁ=|�,��T��g0����x�B�� =='�<*�$��45=�A����$�{���� o���I<j�D���Q<���<iW��s@�<$T=kµ<C~�Z0���@0���B<�0=� ��-8��똽$tA<r�c��2��pj�l�!=)A�;S��=	4���x=�9��A�<k] �[�ּ��$<�n���Fa�7N��O�7=�����=r�=݊]�Ĳ�<4��ێ=JtB<����[�/<���<�N��0=�=U'���>���==?ޖ<n�<��D<��M�<�q����<�1׻�ʼ3e=�75=��<��[=>�C�<��_=j=x�H�=��q<荽Y�����o<?���k�&�rq�[�,�2�l6=�"'=N@��t���f�<!|C=`=��x�F�=��ֻ))�9�t�<��_=��<x`=-��<��<�b=�q���%�܀�<z�;Za��(�f�Yc�;�r<n^@�+�ͼ��W�����f�re=p�1�&�;@ۈ<�'=���<�M��v�:pf����p��.=0�<B����$����#$R=G�s<�x<5Բ<�~�<��&<;�R�@�=�p^:��V�E=m;2=�
��������<��=�w��VjW<(�3�|,�<���B�:w=�IӼ�&<ٜ�=+=�&�m��<�q���r�����O��~D&�>I��(1=	m��TPU=�hs<N켧8N=�a[<t�<�=u9=�D��;�z<��	�ѷ8�ݝ=��d�� >=�ۼS Y=�*F��������p��p�s�-���<�D,���=�0�=@e\=�j=D�<���<j�e���O=�=�^¼׊���=��L��'�R<HI=��>����V����{��(�#Wn��+������;�`�9��d=GG=�0c�ޫ��$7�<8�&;�W=ޯU=�V�<�ڹ<4=
y��A��e�����P�����<U`��}�`�L�<(��$��<�K<<Y:<K�s<i|b=����ة���wi��n�<�g�<��Ƽ>�L<搐<Q�<v�;=�U���C�)�O�n�<�ܼ�ή<�z���V>������A={����C��K=[]����o����^�<Z�(<M=��=�!p��V=��ɺH����=��0�pj�J��:��<�) =-����[=�3���̼��;��)= 5���f0=�����{	�E���+�=/�/��~=�)μ�y�<��<:���Y=`Z�<5�]:f�(���=��-=a�K��'=��o�x;�F=T��:t�-<և=N���{���EOG��&]=H�<�嵼s�������.�\�=��,���?��6� H�����<bk��C��΅<�D
=v"�fi�<�FҺ� �FfмYQR=<�ب<�K�;V)k<�c�<�A�|G���fp���ʼ'R�<\UU�>��<RT�<���=�������ݰ�<�Na�.G=�%�3#��c�:��W=�b;߃n�1Ȟ����<4��;ط<Y"�<*m��р=��Q=�s��SK�=��P=�g2=bC`��*8�f�=\�W�q�;2�O�q��h#�v����gX���;kꂻ7��<o���=���<�L�҃B�����:�ǺE:Ỻ6=��n��ϼV"=�+�<6W=%�<��"�6�=h�A;	�<����ȝ�ۡ� eU���=�ἓ�<f0I�/,����!R`���M�ٓ��x�����O=F���&+�=��=3�ݮ	���=��#=4�<C��6Ze�<.34<��y�Z��ށ=��&�^�<�i=��Q�?3�=S�<TΊ�;�V��Z<<��<@��<{�]=qa;���<e?*=wM}=��T=��*=g�"=���<�~��h(���O�;!�se!=�lu�&�%�p�<��I�t�h�i�'�#�z<��<���<��<�+=�B=��'=�;V7x<V0p�xT�<��?=&/q=�_G�b
f=t<=�˟<�7�<�=���<�`<k�l���<�����!<��0=�A�2x��U�<|6_=bs,=ČD�ձ������'��8�/=�Q(<��=K�L=m���y �4#=���<��<�s<Nh��s?=��w;�#[���P=���;0CZ���F=���98�
�J@=���J�%=Nh?�*g(�����~�<�F=F��<��&<�(1�Q�V=m�d<�΋�0�==�ʼ�8����$Ɇ��U�;LY�<z�K��L<�Y:�M�92$�<��P=�������|����f=��ȼ	hc;�u<=v��#��<���_]a=M�׼�o�<�	6�fRZ=��O=�BE<l�z<�K�# V�Yu���<*�q= ���<Q=J�@�:;5���(���n���;?g��p�<2B�<?wh���_<:�=��?�E5.��TҺx^P��:�/�<�[�<ծ�<�K1=�u��Uft��ܻH&%=��>=r-~�@����:�b	'=�}=�F�<�A��$v��?L���=�ч;��,=X�R�xS�TF=�L�rT�ap=�W<1�;=̳Z�p�<�4�<E=��<4�<����"�|; `%=D�!��l=�U=]�F=�y��7=rݧ<;�ͻ�a�à$=�q��b�=q�;�/�PhL��$����<���;��<Φ#��2L���<���;���<��I�PiF�3�<�.=�%�'��<����QR=N�
�Zɼ�G =mtk��d|=��@��{��밙��pӼhJD<�|0=FS�|�=?UQ���=�_&=]�5�*@��Q=�<�1|��b7=��d=��;�<���^ͼ;����x�<��#="� �_˼�=��%=�F����F_��
�[;*����q=��=��H7[5��R��?q<<k߻C=�`������ =�`�=�I��<�$=�j�<ߛ;�a$�|g�<�<���<��X��/�	R�<q�.�ͿK���3=h��<�s(��Y@=iN����O�ڼ�\H��S=<���mo<N;j=M&�<�k<V0�=�["=H�P=OO`���a����;1�A<��=%1S=�=w-f�b�=81 =6�ڞ�<��8=���o���ؼK�N�ę��K	;����;y�t;Ec<�=���<�c�<^>1=x��; )ϼ�Y�;����&�b2;+P��`���F=���s�,=��*=��_;�Y'�?=�62���7=��<T�q���<�A=�6=(nq=V��K�;<��?<\~<=m�=�3�6�,���<sݰ�R���t=u��<FP���O<D~��b=s1�<i˔�ͼy�'=�/W�Ki��g=���]����ڼd=�ez=\�!=��L����8��<B)��Lp=B	�<���1���lg��b���Ҽn�t=�!=����ꬼ���އ2��n=�P=�^�<���r���r���]ټ��k��{Z�ܩ�<� n� r<���<k��<�g��?���J�)J�;$#ݺ;��<��<ռ8���K<c�#=�(=�*�!��R���?=c�5���μp=�W�<O<MX=�:'�b��z(�;�V�y��t���P=��=[t��މ�t��������_=oFe=��=��,�:>�_=�7=Fd=F�ټ7W�<���&�<N��<l[O�:�U;�V:��U��<;H�< �M�և�<_Ur�۝g�W���OK���;B�*�4��<�O��jk<�-l�E�=�Y<m=1�1��i=@`F�QM���<��<{�<��Q=�/���A��<J�g�,M4<�=e<��E=�!��>Q�����1]�91��-�V<�����7̼����x�+<)<�2�l<[�׼��+���|�j�
=y���D�<\)
=���N��z�<X��<=�X��85��<�#Z�i:�V=eb-=����'�����X<��������<H�A��h=�=Pk=�V�`�2����d͟<Fa�<�/m�|D���'���=�Eu:�x�uK��D=tM��b�U�;H�<���<���\�&��!�?w�<{-=�ڼB\�<!�<��ʼ�Y6���n����<9=ɍM=��4<���<_'N����<, ��h�&�n�=��C~=g�<��<��<�B�<�ć�_
=49����<E[���;�<�9G��~�<1�.��ɏ<��(��
!=L�K=3=�R���$����<�H=o�m�X��;������0���/i=z�a<�:=�5S;�6=�:�f�3=��.=�m\=�D�;��;�it<TO9�iʼ����:��BT<J0;���(mk��=n=�%�;�S�;L�^�F=����P8=^�d�� �TU��#9T��a<e��<�d*�V=k:Fr��JE��1�i���CC��}<>d�<�NU�i&�<l%���U�<!���$� jg=�iƼw��Ĕ;�֣�<�>=����n=�܁<� <��!=�T(=��K��r<�*}�°������x��<���9�K�;5�5<�/����:bA<�gP��=�m��H����L��.�<߭�����K�R�kN�<>eW���<�^��A�<T�8<Zڻ��7��ݯ<4P)��A#�'s�<G�9=��<O�.��e����z�k��Rw6=�B���"��;b8�:e�$���ļ�6�<���<��߼:�j<D^=�a=��<�9��B?p<���[x�=���s�=��$= lC=�/=%@�0��D�*=���������<U�H;�+�<�5�<BP�<��K1�$=ty���zx=!V�<�u_=-\0��T��Sɇ�F:�o0�<�~��<�
����$�u񼵀.=�U<���~	��8<�ki<b�(��=�7�;%Bۼ�C��: =�%_<�(���<B(H=�C�3��m�0�5aZ:`kA��R:���6=E:=:䘼K� =i�$��<U�g�\����#/=�h�,кM�&=�s�<�W��li= �*����¿�����":-8=^>=B���~	�;�޾����<�¼���k�=T�_=MRF�9�p�Bq��$- =�^��Z�;^9�v�>��-=ǚ�<C#��`��IV=O�j<9�F<.�ɺ͆G=�z5��ZZ��)�;qz7���H���L\��p#�˭x=��'=v��4?G=!k���1ݼnb�Yۀ=�%�}w����;�4^��e�����<�#=�/ڼ�=�L=�^�q�N��0�<&)�<k5��YV���=o;=��n<��;=:XԼ�4¼�\=��=�#��8�o��I�=���#v�<h,I=��0=�B�D�a=߼���:�}���h�<au�<���<�H{����"^�p1��<TL⼆W�;cɗ;[�=��j<`U=�@=��?<F;��b�B��Dr<�h�&M=�BN<#|��^0=�f	�,|L=�i=
�3�,iؼyn=���P�<��z�S��<����
Y=B�h��G��Ʈ<r�w��
&�(̺��z<��,=^o]=�$�'.�?�%�I���z�-�Ǽ�;���� =Bn<��B=� �|�=��	=�}ջ-�q���u�'�w��һ���<��<�!=y$<M<<ht�:�q�;h"�;�m#�}�=gX�<�3=dU�F�]= �A����==�'�<n~P�Vм��N=��P=�ͽ<�w<�k��<�mj<��2=�f�;F[-�u7=�MI<'p�;5 ��|:�<ݳ�|���AF���JM�@�%=t1)<*Cb=�9�}�9�R=ה�<�`���-��\�<��{<������+=�4���='�Q=4uq��<=L^=�5�jP=jx=�8��ɺ�3�<ϲF<{�¼ɦ���=�c�&���=�i�=��5<��<�M�Yu�<�n��M 7����<#`f=GC����Z2^�$,�%��<D�=9�s���+�U	��ڻ��~���<
é:i�<� =��=�%=[�(�{lD����R�<T
��S,�j��;�t���=8��;T�{��w��.������+k�<��j�>A=���d9G�$V�=<�>=�`���SX<v3�k���Jg�����f����@)<����m	=���\_
�TFa=��=X��<�=�D���|`�,�+=�Ҽ�P'=S��h!?��>;��1�>�W=]��<yMm;`Í<-��x��<���q�V<
�Ӻ?�A=��=ʠ.�R�y=�I�;��<#1=6@K=S�X=�4=�&=)=#/i�t�<17���+.=[~�<�v��?�$=���<id�ha�xT/=�T���J���{=-�i�ؼ,/��~�815=P4<��=�#ʙ: �y���i�j�����=ރg�থ<��ɞ=4�3�W�ջ�|�;��G��|I=��&���<"�l�|=&=E��"�<���<�i\�	�l<G9N�i��<��=����(�<�Q���7R=(�4<��d�ӕg=+�ؼ�"=�V�<$	�<�6<f���S��dT=Z��<�
J=#w����
�>A�;n�a�ڪ��f������G</�$sn=s��<����t@�O =SƵ<���o�4<a]�<R�S��O���<��;��"��1)��VԼz�O="�S���'��h��/���n��;/=|��<;YU=Ɛؼ8餼���;�#�iQ�.��<�$�<�D�# <��e?���<Z��h;	�\��;�켫?V����l����`=�<)=q<s��
�<4cU=��n���ƪ3<�yA���a=� <��=w/J=?&��G�<J4ͼ_�&���Լ��p�[a�ϐc=��<ϗؼ`�m���?�� ��]�=�䂽a�^<z��?�=+��ґ����(��u�;��:�s����b�7x�;�G��i��z���H=B�.=B�'=��Q���=�%����;-�1=�-��*>=�	�iU=�x�;5�-=[' =�E�;6�<\�z��˳����ڏ�C�*�	=���1���*���N=Y�8�H\=]`=<=[<%�$�&�v�\I����0�؏�<��l=C�x=NCH�gc<�ke1�D�a���<?z<@ʹ�4�<��9=P=:� =�Z��\I=eq�� E�eO8=��<�=�=o9=�m�dr0=�Oo�?pP���&�G�C�C=�19=�o���5��V<"�<HWƼ	��<J4'=�^=��$=�v�<������;�7�<���<�nt�2�߼`^��r�<�[)�F"���2=+��<S¹���:�~�	=��e��20=0��(�"<�^ۼ�d�=��=zH�y�,<F���9����/=J�S;#�N�p��<#LC=���=Ss�T?)=r5<�M���N=�P<o]w��<�<�V��i9�r<=�Q=V�G��j=�Ӻ���;���O�&=f��%̑�E��������=�3�����T�3=x"�<~�F��d<Z��<S�<e�=�M]=������A=ך�<�K.<6��<{@軠L�<��G<�١<Ե��b�����f�\.��P=>���=�=�4Ҽnb=2zﺇ.8=� ��(Μ;1��ۻK���|=8�W=wf�<C�=�P[�J��<�E<B��;3-�|I	=ٓ[��$=
t�;|W�<��<K����x=�fk�  �;�Y=�2�<����B���2�<�\=�D޼]�S=�f�Ĵ<ĥ �7o�Xݼ�b`��rW=j�<FD:=R�?=��G�)Ǽu�'=́�;��&=��C=�i<�W=���%ż�=eXg=a�_=�x@=ط]��1=1`5=�� �4�u��j=�F�;� G������i=��[�¼�<��b��W�;���71a<Ăj��5T<��<�|�*?�;��<��E��<�k\��+==P�-=LnR=�ԁ���H�b���0�=�ܧ��������[d=	��*�~�7�1�S=dZ
�a�;<�6���=<J1�W�E�c=l[=B�Q=�3Q<�UW=I�G<��=�S�)��:��<���<�G�A��;������<��X=nN=��<x����U��N���1ʼ��=��>=
��������<:�ԣ"�[B��4�� м���<Vl�;~hO��ؘ�J�1�i�����=�"L=|���/����A"�	1�<V�����AI=	��<��<��=�z�"�<|ij�����v��1�<4� <���f�<�Y���< �	������i�kh�<����U�ߋR=��k�bPD�{U=���W��Ç=>��_{	<*8���'H=��U==]�<6�]<��d=(��<��)<d���<{RT��-�;~b`�t�%<����&���N<b\<=���#ؼ~�<�r�<����X1<�����3�d�W=����t�<��U�]��RE��C�<�3Y�f<˶�<*Z[�b�*=Х<��<���9�<�<8�4=�V=1�1=F-C�ؗ�<XC8��p"��7=��.��=��H�Δ=?P�o�_�o�߼�|�\�<n��<o�����C�a�����%�W(��Uc=�v=�K�<N=R~���Td<��Y���㼼���-��<�8�����<���<7�=Լv=�F!=���㼬�Q=�o�a�<�\)�� =Yh�<l7�0)ʻ��y���=�(��}=�<h�"�G�~�<�jB=��9���V;���a��;#��<X��<f�漲��<)��<�>�<r���#S�G�<���<���)��e=<<a���;�"><�)��AT����<��c��=�M=�	�;���=Vo��'Z(����	˜�ώJ=^n�<Z�=�#,:j9�I���@a�:|`=K�<;*�4�2=u�=�Q�Ru�=����Լ�(��`i����< �H<�<��� 4Z=��=�b�؛�<�,��|��:U�<F���	/�x,H=S�=<ʟ���j^<,��n��;� =��*=��<�<��>���#=���bY�<�d:�`��<��K=&ռ��T<\n�<�����I=P�Z���/�1eP=z0�<�KɼE�������[�<p��<�&%�9=A�==��ȹ�='����N[<��=��¼�zh<��==U�?=\�A=��ټv��D;��=����<x���0]4=y{=8S���X=���;CM���.��r�<�Ua�J�-<7W<F�|<�s�<wl:vc=N-=땼�E�;jl<�u.��R����ұ<��껨�@��[:͑Z=R��<��T�������-:���<r\�\f=��e�a=�x�<���@�jo<��&$=U����D��c��?0�p7-���=��=�Q
=Z�������<n�:e�<��`���<D����xS=����rl;�=�#)���;=��=���-�K�pQ�<�*=Zt=���?�KZ�:�B<<�V�5A�<��c=]�4���~=
���=D==����t�<�d�;؊a=ٙ_��z
��x<t� �"�ȼ.�<��9,�G�&=S�����V��� $�;`k;�N�����&`�:JE�[��<�=��=tS#�����/�=��A=�X@=�YV�u'=�>��üˉ<�3�<���<��w<�K;��<2O[=ؤb<e)S=�7��|���\X�F��Z���]�g}�<�	߼8��9F
= =�!=�ء�}n=�"���<Cr�=�v���r=��<�}=繈<g��%=)P�>G�<�l=��.d��P=�Y���@��e�
F:=���<G�D�#m�<Y���8w]��z<��̻�)�h��<c���(�<Q럼�_<~�=v�=�'*=��m��*Z<%�$<&�<X/m=�w���f4�:ͺ����Db=� �W��@�<�(�(LO���٦u<r.�;f��s϶<q�y�U�0=nC8�����<��=p]<��J=m�n�U��<ĩ<ϭv<�5�:��;=dQ=N�=������_��I���%F=�bH=�,��%`ʺ�[�<rٰ<�g0=҃	���B�o�y<����D�X�i�Y��K�=��׻Yx,<����>���=��q�������<#�,��e8=`(=���
�׻���|=wx4=��2<��5=��߼��T�y�1��Y<~5�(�X=���d7��P
<�<�-x=3�m�	 �<��=�D=݁v�
@I���M<�x<ƅZ��zm�Sf:=-U�<<�;0�=x�� ջK��<���s�p������<�+�<��O�?=f$�Q�&=����'�Kv���=<��J��R;{G0=0��w���h�b=��;H�j<4d&���7�Aٱ<��=�EO���c���?��������\���F=�V����
�<��=����r��;�p�;�V3�u�J�q�<)����T�</=����5��!?�|a�<d�=�0!���J ��&+=�����<"��ɍ�xa��B��^�<�W����=ު��H�j��=<>Y���k���X��yE<2Xg=�r�=�*=;�;&=��j�W�=?5=���<��=�Dc��#:=c����=ii�<��8��ŝ�¼�Ȓ{=s����՜;D�<۸�<��;��.��=.{!��7A=%�%��p�JHм�d4=ya��L0= �3�5N�<�X=�k;������O�X��<�żl�7=�v =,�	�(�2=A����X�;��<��H����}�i`�;��b:�$*<X9�������h,�:>=E��;��!<:�����0��<�����;'�/�͏�/�Q�a�J<A/1=f�ѺƝ�!9�<d���Q��9=�n2��&&�c�=�
#�bEl�s�<A��;�`�+��<�D=o��<�����<=�ѐ���<Bؼ<M���:Ւ<+"=2�,�2E���X���=���ݨ������>��h�Ɉ,��$u����ы�<�Ŷ�& ;�t<`��<��<�
=u��<�Tj�ZR��=񏰼vD�I��y	=���	ί��\#=�Ԍ����<gk;Ea=�A%=v;[�y>�����亙�:�	=tIɸ��Njc=M���|��<c���m/��m�<�O=�"E�{�==���<2M'��*j�2�ؼ��<K�C="��;:z	�?��=&�¼=�	��R;��p�Vx=�g�+�I=L�4���,�@���f�^��R�<���:�<.:�F�<���<�d.=P<�&�l=��C�zҰ<6ky�)_��l�=C�$;�;��'��<�xF�K�<hҼ�ES�70�<ml=��̼o
���n�K�k=T��<�6�~̺<	�7�s��߻�͕�r���d��;J	����!���;�|�<�u<qʅ�mgX���;�p)=���<)O��y����=jɫ<(��;g�c<N}9�	\)��Z��;�;�<=��)<���<�����<�-<�3 ���=����-��<#]����S<�\һ�<9�(L�<oF5<�05=`؄=k�F=Bf�;4@ɻ���������ӼV,�<u�"=��b��}���C���_�!��<�D�<͕7���;� �<��U=~J��vJ=��ﻴ�<<�</���W�;��N�W��Z@=Ư0=	
��0�C��XP�?��<�]��	�<_{c��W= m�=U��<��Q<Ty��=uOE��#K��iE� M�<����=�Z�-e-=h��<S1y=
'=�;8=(�\=�g\=�Ĭ<aS5�t�4�~�m<?�<=v�A��U߼��<��<��<��-�X뺄fM�H4�A
*���<z\=ޡ����/���[�20�:fĔ��k=y�<�f��LT=�k<DE�<��D=�X�	帼WΘ��؃=�ۚ<��;�����c%�	l�<�,�gV�L9���7�<*���=���¹iQ=�a�f����Y�<xG=C4�<ń<�h�g��:����aD=� Y�׿%��;J=F�5<`R={�=��I�ؿ��J�����ڼ�b;���W[��2=iaM=_2-��G=..���9=�i���bn=��Ҽ�H;�T��M�<�W<ׂ=��<�����&��b��<=	�;`?��� =U�=JS:��<S�A���=�_�t�4=�!�����<U�)=/A<S����==��<=�+�L�=�I7=u[�<>43�Ԝ{�T���x����<+��;M�-���Y���9=�=���;�PL�?��<�}�<��@
U=�t
=xP�6��w�P=-#k;D�<_�!=J,^�NP<�꫼A>2�A =�<=�4q��ā<�f����|<��W��NA�_�=S��<ݴD=pd=;�; W�A��z$=�9�<�0���(=x�!=#���#m�=A5H��b*:�[:��љ�t�=3�4=�����3=�ax=EV�N�,�ŋ��_=���V�<����NZD=1gV=��\�N5�8�>=c
��s�����^=�/;�L�<N3�<۷w�#���58��8=�(��������7=�
=�j];N+=�V���dE<)MY����c��O7 =&K=�"=�d��4�� Q<��4��<6��9=vq=9%�<���I�>=|zn;�G =G�Z=�B��"/=��[=��<�yD<w<<�Kt�=��=��U={�����<wa�A8E<�g=q|(=dz��J>U;�$�
5q<�;��?�����_�qTM���=��<���㚽��+� D;��R���������-Q'���d=yx�;���Z�<�c���Z�<4w�:�^Y=���<p�����<�2^����<L>�9={ߣ�����_������,�o�_j������5=��E�-b\��41=����C�0��>��v�<�
�U��;�׻r�C�sT��̨��[=4����<œa�pJ <'����<J�H<sr�=�%���¼J�D�/��<������W�:=х�<�)�x���ħ1=���<�o��1�;��)�"K�;|~!;|p�Z�B���_<i�=K=5]��O�a%<�l/=���<>7=)����>�F"=Z�6��@�d"E��4�o�/<� |�%�k�U��=*-6=�,?�a3=}h�<(�;�J�T�;Yi�<,�D=#���i=a�����S;D �<�"<�������D��I���=����[J��� ��=u3�;�%���m<�O=*ڝ<,�?��^Z<)ٳ���c=-�>��-��iZS�r���<72>��<=�8Ƽ�먺�C�����;�{Ҽ�9}���E=��i���<�����|h������o=�y�=�q�<��9=�Ϡ<�W�'j���<7��<�X�<U�0=�'8=bv���Ќ=y�\�U"-��AO�8[N����=i=0I=)ü�3��3�<'qo�*��<����P=xG�Yݎ<��޼�P=׆=}��<$�&=8�&�0�H=��=�ik�0���o�;<����~<�Y\��7�<�9����;��{ �-��e�<.ۜ�*b�<���<�A��]�A�l?<z$P=�м;us=H<����������:�n��>�/�b���J=*��<�D��-�>��0S�*)�<�W�bk]=��z� =�m���8�<�Hf��A#=n�)<%V_<�B�<���<�׵;�֣���=��<Z�G�f��u=�M]=J�=�Xr��v/=������;���<����>U�^�<��C<,����;�(#��W=Fj3��3κHv<A��[K���=Q	<��q=S�j<�%R=�;�5j�N]���
��9F��8�<�{K���伫z.=�^=?!��P^<�+�;�{���%A��f�<��xC=}�����=N=���;�BN8BQ�=,�Ѽ�=�=2"���e�9��FHؼ,9=Y��<��;.=�14�v�޼�}�<t��<��5==!��l�<��=6=����ڏ8=,�G���=%TN=��<[;4=D�U�,՛<�
��c%L=����>�=vkT��r�<j=�,"=�_$�]���J�<���<� �O��[� ;�;U�:v<r?"=O�;u�H=E�b�HK)�*�j=j�<��9=;�<����m>=�l���d�,<���ռ�K:���g�Sg��1�Y����'�������꼃f:=�;���x5�ߏ�<f]W=��x<�K�a94<�EK�5?=�l ��$b<� T=�"W=�	E�H��<� =bO=�y���üE�#=��Ǽ�j���^�E�����t��)�<n)��6<v=�2-������?�ǼG�k��I<8�<?�S;@Լ<�̢���<sX��6Ā�r�X<}��i�<�%9X�3��g<���߼��k=���ơ1=5�-=�S=�Й;
t���"��� +=3�C<���<.P[=%k<4A=��1=b��J�C��9�o=PK.=p��<I��<I��<�z;k�o~='�=8}�<�9��g򡼟�i�G ��t�<�N�=`��ټ3<}v(���;GC=�5�;�~��+iE���<��<��=(�j�ċY�7:~=4����<�<$�e=�LM�5��hZ=��Z=��wV���`�<y�<N�μu�9�Xa��u�+<f����РZ=�ˁ<��=��<��:��;�z�M2h�:Y�Q�<7ż8Q��;`=���<e�"=ZN=�k��",��P!���mP=E��<��ּo7�;�\=%wk=j׮:�9I<�ڼ+���`��TT=�#�;��5=y�I�R�+���5��L��=c�=�1�W'�%&����<k~`��5��J�-_��(s�٨!=�ڂ�h�Y��Ա�;@	T���S�3�I=��9����<��*�}A1=��R<���<`��������?�S] �/�ļ!t������<�v;
=6���S=��<b�H���;�+=��<�J����@g�����=�`W<����y��9�;���j =�m=W�)=���<�`
�k�%=�=�ƥ<Zn<�J.=��;��W�*=b4�Ap�<ӳ��"�<=䔼J,�����<��`�;�犼{�O�`����,��N���?=���Ir=��̼Ʌ���;!��<�w#��"<*�=fLH=CT���V�_�	=.���lN�9p��kk���vU�Rb(�-�<J�<�%>=u���%�<J�b�vSԻX��<��\=$��<QLW=U�]=7"���=�>���M[���;��ü0CK��v=ey=.)8<W .�<@���!4=�-=����~�=�b|����<�Y��+0�����7{�*�|��
=�>���8�� x=��<d�ջ�=�`C���7=���<�Za<���<�h����.��#�<��I�PϼSq?;�=�A�`� ��fh=YA1=r�	��p�;I�=!J�:��O�n윸���A�<���<!�<�.D���4<V�<䩼+C��]#����<��"�M��`b�<�ϼpL���������K�'���	=ZW���=�h=�`D=�����z���&��c=��=�O��<�j=r�<�W
=BFt<��8��;�18��һ#��`KJ���l=���$=-<����r���:g��`=8�V����<c�Q���u�x�3<�6����8 �<�FJ��ּ��K�-Y�<���:���<=� ��ڤ<�va��:=$�&=j�V<�u���h=�iH�$=�p]����:f��;��h=��c�S�U��;-��t��g鈽�K;zyR��u|<��v;:Ϭ<�n�<��#���G�\⧼na��z����o<4%ػ���YZ;��<Ό�;��ȶ����<�^� �^��b�O=��O=^�<��<@ =1i�<5|c=}7=1j��)���Aչ�=���<38[=�[;�j=��n�y`��!���w�9�pG���<�2�����;�!1�I(̼��9�� =(<�=I���K<�<�vs=�37��?�<'���LN��5=L=�tr���<�S��y���7�<��N��d�`㼆�� 0��'�;bc<�
%=�x�<��5=R�ƼڍJ�+���Z�<�ȿ��#i=��T<,�����'�-z�;k=��w҈��CO�U��KJ=�i=��:�.�a�N=������0�	�+��<����/=�<�U_0�p�%=��=��=v��<_������Y4���`<��=[+U��=�pS�
hE�>���6k<F?|;���$�ٹ�G-���<���OM=�ۼw��v�"<dY�(��;��&���=��_�^�<�<xx�w#R�%��u»��=�<>^5��)#;�zU=QxX��VU;`*�<�H<�=��:P�<#�0��\�=r��;5=y����/���a�n�*="+];BO���1=�\=,E���t�$D&=>&;���<������<l�U���I=�����w�/	�_Z�<��K<wI-=��<=���Hm���<C��<)�z<DB��KA=+�5�,��<��T��m9=!ʹR����H=P��а5=(6�<��F=�Gl��X=c�;'�\��;�<��<,�Y��t6��G=�r�<��p�ܣ���$�<2�d�,��F���I=����<4�gu(��0��M-p=�Y��^
ܹ%~,=l���(���S�l�=��=K���5c�;i�ӼHÜ;��==漲��;0��<	(<#�'�Z
��Y8=��<�5�;J0Ἆ����E�<0�=D�t���<i�"��G�={K����<w�L�c�a�'�g=nK,��;��P=�#=k�@4=�>v�"82��M`<���<��r�Xu=���<��p��S;=T:=�^=],&=�&<��=DK��[�<Ta=�i�n}R�AB=YPv�i9��L;�qh=�h\��w�<]�M=u @=�]��%�D����9Y�c��\���Rt��3�	J=�	=Lw=.�=!籼雹����<@�s��j>�Du=V(����:̓�;)F"=�
�n@=�d�<�7X=;��V��e�<���_ƅ�f��<�����e� V�<� �ĺm�2�\= 9�=��o<��F�<�=k�u;=o�3����*��47=H?=��<aqU��c< 1�<��;�]���#=�{�� E=�!=��<۟<[��Z��)=֥��S_=��<�޻��D<L�roA;Hɯ<=��<i�f�Rߛ;'�(;��L��-����;�7��%=�O�<!M�"=]��<�<6% ��du�|������=�PS=���<r>=��t�1J�<~=����#6�\6�E�)��;�<�$-<�!=�`��}4�<C&\=�y���=��m�ӈ=�� �J�?��<Q����!=��<�e1��Ȃ�'豼��*��ż&G��1k�<�<%��6&�ژ=�	+=ݥ=��*<�Ӭ��4��]���=�<���:�����x_��nw=Rb����;V�X=i7�<���;��3=M#�<�o�<��6<�Lڼ�Z���=3=���Ҽ�q����$�>��ܼ���<"G7�Kw�;w"<!��<��=ǒ���#=?�<�yҼ�ր;~�g���4�6yļy=E�׻�݇=�0ټ��g=S|l=}ɮ��o@=��c��{0���=�՛8�;��O=�9��6W=��=n=�j�T�k�/�<�ti�����?�<�I�h*�<|k<<�!;�2=b�	�GqY�K�D=|�]�}z3����;��S��<�4=�s=BB?=m{�;~�*jf=e����}Z�du���(.��¼��=HҦ;W;�<��=��f��M�< �=��꺍��<�.=�0=��	u��=.�-)n��D���J*=!�=��ټ��!=��<��ty-�6|��w�<�2[��aw=$�M=��?�-�ϼ��=��%=�MX��I=0_�<��=���<]�M��p<Q���a��qR@=�?=��Y=��+<�)�a�<y4Ӽ�3+=4l=_P
�� ��-�d;��=u�R;���}؇;y:=8
�<�Ix�|dn=��9�$��;�Qk��<=�����g�%��;KL�Q@Ƽ�l.��.���(=�-�����;��={��<ܑE��/.=OF�<%��<꒼w�<[��<��Y=�=��K=^�*<��M<c�)��'/=��:�@|k=DI�N=��u@=���A���ch�x�0<�dX�G�)�ӃM�;^=!�F��9����=.��XX�<��1�E�'=^�<2�G=�|�x�<�`=k)==I8,��Ԗ<)�8��Q��|;=�3=O伟oX=��g�#F;0�m<0,����<Vh��P�-�q{�:%;��h1��W����\!�<={<����F�<A`Z=��+����;�o���kM�/�f=���*��9�$�?*=��=���k�����=�*���"�P��9��BL�u�������bY<Ҙ����
�:���?=�Cϼu ��w���W=�� =�5y=����_=�,�<�����aI<��<�-����A=G�<h��2"I=��~=��]��!<!=M=t\�����;�	� �`=�@=wv=�d=슎�AD��N�B=sL�s�Ƽ�`ͼ�T=� C���ּ��W=�v�<�~k�������X=V����v�R�d�~�>=�kr=�6<����Y�]܁��s��U=��)=bd��8�	=*W=*X�<����.�<`b����G=�xջ��8=�Q<~#r��u˼\;��G=`V��|��KP=�Ł�*�1�4����5=�\�<e>0���ܼ�j�4�=}7�<<�=H�=��ڼU3�<��4�
.0=y��<�A=��<ƭ�<�
鼹W_��%5=�b����*
=+ =_E�<{SL;��d<}�b=�"��W�����@K=x�,=�	=}�\=��㗂=�Ռ����<B�3=g�<���<Lyh��=��/��Ү<��?=z�;��==�1t;�Y��Z�R���&��\�<1�
=ݾ/=2�ڼ�����<4Y��D<�YK�G��N�l�,<�Nʻ<B =��ڼٲ8=�+���?�ɮ�<�L���a��Ƽ�0�g���(�����<#�G�zVҼ��&=�[���z:��0�<{=i��<L�;{����t;ڿ<�Q�;�;=d�<�s!=�R�<��鼐C�<Z��?A9=\�<)M�<k�W=}�<|��<1��<i�<�-=$ϼ���<?f]<η
�v.���9=ι���l��<��=��S�\�'~��=��=�]^=tF�{o�<5�L���Ҽ��=V�.=&�J�:;
�hIl��A��s&�!�@=5���K�<c�<�L�:S�:�j�;��<A<؞<\��;.�F=��ü��2=*�;R<'���;'=0���L��0���<M'�<�����k^=�Q�<�\=��9��F=;&�<�;0���Y��C=�=��;Vd�<L�P=�����aü&_^=Q��;N6f= E5���¼�}<Ĉ�<���<�
�<�Uw< H�^v����|<u���6<���l�e=�/1=ޚV=�$Q��}�<DQ�=IN<�l�<����z^=Q���u�����<��;e<O�}��w
<�R��P�=3�ι���<;�e��r�<��<�7�0w�e6�����k/$������g��<�9h�,�t<��4���b</lX<�J�<��Z=�8�/�&=#�|=7��<�����0�R��<U=<��<md�<XM=�h�1�2=�!�"��;�b�%)=/?K��Y=XЊ<�t�d�;=���<k9F�1R����J��e�M|9���׼J<`;Z鼛>������mѻ�!�<s�@� 0<&���<==��=��)��^¼�-�<��d;�.=������Ȼu)��N;���M����;2�g�n<E˹;ht=��:��R������=���<`�<"��<��=wI�c�`=�@=N�o�k	�<�� =����޼�l��7�:L�R=Uu4�v�^������5<#�]��,���@=켊;��nT=�t���m�L��<�<<Pjܺ�$<��~�0��7_�1�i�.zλ��弍�<=��M�;=@�<������='��<m�<l�6=�"4;;���*	=��*�;:A��=:J�/cz�u�G<�Ɔ�_�B<0U=�� =�}�;���<��<2E'�C�`�K�a=J�	�-�T�`=�>�b=��=p^�<#b��E�<3*�<����t =�I���?����9K=BUa���5=��M�������<d�_��(/=i�Y�zfE=�IX�(}R�F��=�S�<n�ݼ��5<��H��}���S���f���
���=��m�$7<��b=��<s�&��uS�۔(=7U;�F<�A�<�=�<��<=?�<�0=$M<y�<� M��+�<G!
��Y@=��9h%=�����N����'��<���]�R��{�:nvּ1,=�0=ʺ����S����m�<��7�>yi<�`��";�J=�C =e��8�v='W!�ȧ���h�Ϥ�����U=�7�[ƛ���=X�J���o<U��<iN��Zh=޵�������^5�\��ބ�d9ʼ��C=��<,�<��j�~Fl<��_�{�7;�s�:kv�=���� ��".�Vd;C)=���1P<_ů��P]�q�<����3�<i-z��Em=&l�<o�2=�t��-t�����(�:=a�)=f�1�z�<ҫ���U����V�B<b�79��}��H�9!<<�<��<�"S<(�<�
P��?���=�#=��������5�����Y��?H=��-�N��ߜ{<s6;�|�;�sI<?q����=4X/���=@p]=b[���,��'���H��P�A�<�n!�*|p;v<8���]<��_�;NQ=��?��=�?��.L���	=�e�=�g�l�;����c=�s
=��;`�;<瞧��w�;�Ѽy �7k�=΢���<PA༆c���ɼ;.�;�|S��.��f�R���／�,=�3���ϼ�D̼o�=�@�=�(����3�8��;ۈt�	�q==�B=Ot�98=R�<|$�[���K�!�J�`=���#�����c�>��<����������4F�R^���0��pY<헯���<z��<Ͻ��f0[=c�"����;�ͦ;���<�w���D�<��.:=�4<Tr]=*1��({�D`"=��ѻ6~?=�輝�V�p�<F�ͼ*�;��ECY��2�<�ך;�U>=r���[=�B=�*��#C��m7���);ts��l:=���GYb<E�ݼܬ�=�$`=/z=2���3`=Kֺ��v=/�c��2�<X�켥�ͼ�y:<~���<ա:<��`<)��<��{=L�Ӽ�᤼��;I����.$��Y=��]:奻��;af=Q`X���Ѽҿl�|,"=N=�:R��<�w�<v�<��i��=: �|F�J2���
ļ5�����<��F=���<x;���,=o�7=w#��f���!L=D��<p����<Ce��@='�\=a�5���=��< ļ��!���+=�O��~#�{^�t�<�~��D��޿���v�7Iy�!��Q�3<����=�I�<�MN=;Ӣ�E�8=��J�10��O�;�!/=󤅺�y�����<E�=�Ђ=��
��I<�3=w�/���<ׁ4�Rn3:�%=sX�;P<�<���;B'+=��ĻU7d��(=��Y�u�<�=�g�=j�ۼ�>=/�4=�����B�e�}=h|L��S@=�4?�B�]�����	�#�ש=�
<=�c��+L��$�E�%%F=�ɼ[���p< .=�`a��fɼ�e�:�����K����i�L=��<�<a���ս(���D�'����A�)@;����<z������$��<T��;���<.X�)y���;'�<ʯe�]�ܺ�=߷Z�M=D�\<UQI�>�y��w�c�
���E=�?��sG5�"6R�Ǵ)��j1;��-�<a��<uO[��s�<+�\=�Ƶ<D<�u<V��;�Vm�O�����Dj=�`=꾼���;�h=����=bN"�MY���z�B�$�� 6��z�<姫<��r�K[�<�üPF,=�Ь<'�3��;F�<v�����<C�L���=�:�����;�!��$^=�M=��?=Ȃ�����<��x�E{�<y�=��b��siC=�WJ���j<A��<��=�R}�}��;�༉A�<��U=b�2�[c�=T��q���>��<���{`<��\���	�A� =P4=��:7w&���1=�蘼�k�<�th=%=:�7��9�<rƬ��,=�@���=��#:�Tȼ��;:;���0g=�/�<�]>�(=�S6:�)5��|=:�"�Ƽӭ<�����_��i�����*=s�E�t��<��$�<K*d��L <���*�_��bV���u9�{�<�&�<��D=��:�8�<�mZ�����J=�{�<�-�=��Y=wf�)켗$ �5�T�<�+=��s<h�v<�	ü�?=�<��z�T�$=�4N<��<0��"<���:d�2���{�z�~=����Vk<q~�����<�6�;�=g2�;���X�u=Hx'=��8�O�����Z=�Ut���<�=��5�<�-��[� 3d=�����=�o<� #���	;�u=�OJ=؀#��'��`���d;���. ;�<zr��k�Y����<COD=�*c��O�ń��j�=t��j� ���%�<H,=_w=up=H�=f�=j�"��SK��@�<ƭ<g�*�C$+��8��c�˼F-c<�J�<7�p;�8˼�<p=h��<AɼheW<��6:D=}�{���<�h<ݙ<H1=�kY�@<�.�<x5�<Nc$=�u&=��n�"�&��͞<|�!�<�ü]�W=�;�Q�=p�
�疘<�Mջ �5='�߻�.*=�i
=���޳C�����9l<6���%�e#2��;��!���<PZ�;j�;�� W�����]��H
м�1Y<�L��)E�0u&=�5�<���G��˼�<�ކ<{:��#p�~Ͷ<��O=Y���<{'�<*͕����<)�n����*�r=\���ϼ�(F=�B={�K=Jm`<����/s�e4W;������<k~⹀�<�t���[�$��<���<.��={=-�a�����t@=^{l��O��@1=Y����f=�UH�����sv=�j�<� ���<�k�<�
H={�$��r��LuZ�Ry=/�<�9=1�#<$ <g���+�<���خ�<�8��]�<�q==n.D=|�Y��9K�v��<ub̼���<��E��!��5R�O=ȓ<Pvd=UV�e�%;��<�=�<g?t��&�; T�:V��<�����n<���8��f���ʻ3&�Hƹ<b�:+�<y��A<�r�'E����	��vؼ�l�=L�_���N=�x�[�ļ�7�y�D<i7��<f=�b�<	�<���;���;����xX=NC=M<�-�����?���l�<�`����;Ӊ\�	�:��ɼC�8����*m�<��<w5=��<�;��`Q���<�_;�5�(=O\=���<�y<P�<B�x=HP�<?_-��v�`�<=��ʊN�:=6+A=�Ё�9?�<:2<�~=�ͼ|5�{�"��R=�?�-�̼�7�~��_��[�<�$�Ģ=Vͅ��8H��-=�����cѺi�<�<,:�ҼZ|�<8�7=��|���<MU<��G�=@��;��R^�+�<n����I�~ =)�3=#7`<�6=A�! .�����έ�J�P<l	Q=Z�C�zK���@�;-ˈ<��f��=;>l�v²<Un���w��Zҭ�n�@���k�n���z��;��[��Z=4i���Bp�=�/��	���Z�l)����]���q)���4���7<P��U�;�|=@;A�K�9�ӌ=�'Jf=g�=P`E=|&�<eA���WD��M�<O�`<��;��O<�]7�Z	����<!u���x=���U�=MEO=�2�<�x0=S�<�E=�/ �����.�q��x�S��\�<�8�<j���{�V�����k���ٿ=�^�<x����:�	�H�M�v?;@����uI�
wu�,�"?R�3���;=q���!=��<�R9�*=��=���<_�J=�[Ӽ���<����WK=r�:G(����=^[���0���;+�)=��i={�A=���s�=I��A���HG<�(�D=G/���`���<t�A= y�;Mˢ���i= �A��=M=��=��a���d��J���@=3�;�>�={�Y=��g��9D����;�'V��J���;H���俅=('"=d�J�31H=��ڼlt2���<<��G���1���<�G�����<�H@=��X<1e7�M˧��k��f�k="�Q��
z=R�5=��⼀��<"J<�1�<ۍ<���<�<�U�=�)��c�q�4��;@ռg%�;9-s��=ɻV�<<�A<μB=o[��?=Yh�3�0=uM�m��<�N1=�Ž<�3�;�;|=��<�o�2=�<���oZ���=n��<Ks={d��m�ҼaJ�2ި<]7����J=�ʼ>?J�<N�e�����<�̆�I75<:.]=��Wh1=�J�z��RJ�<f�e���I�F�s<'|�K��<�aB=��A�t�=����v�8=Ëw�=��ǌ=�8��k8�GOz=~�!��jV��V =�q��W	;��a�<�żO��<�8�<�.F����<��*� ���:�<^[��\�;Wq��)�><a��<�H��R���úO�^<T�O{�<�z<weɼ�p=_yg���J=m¯<�[C���v�M��<���:���;1���n�.=�֬<��мW�<r29==2<9�滁�#<���޵D��L���<!y����#=>�C<LJ�<*����;��E=V�;�M�w���V�;��T<t��<��?=�!T�N9��l�LQ�<LaQ���<9�Ӽoּ��q=,��$��4l7����:�*����P�U=Q�� �ṙ�>��*ܻ=0<V�K=_>�FT�:��<��l�Ă=v.��.<����4=�v�;�2��+/@�J�"=vH��u�^����o�p��[~�x�@��]�;=�<�H����P:=CN7=��v��?(<�N�<��X=Ǳ���M�K]	��7��[�H�=����Ŭ�:��n���	=��<�Pj=n��rL�s��<�۱�T=/յ�&'i������k�w7�<��D��D9=Xc��l�;d=��vw�;@o�</��;o^[=�i=����DN�<��g�}8���5�<rc=���<t��<�H���ka=�Em�}6.���`���os=�D��d�̼�a���<�==m%�\�4=��d�gU=`	,�oټ<��e=ֽb=��]:�(=ޠͼ�y=��V=e�w;|/=�o�9uU�m�;���<1�l<�Sμu�x<y	.�&��uE�<e%�s�<D,�<U�лhM�<�*F=&�;3���,i�<D�i=ڥ��&#�;�=\m�<��x=L�j��v?=VA~��{�<"�#�K����<55����� �0��Q�u���Az=���12,���t�nVF=%Fm����<~�6=`-�;#��;8��<&�=-�;��<$7;�n(<m��@y���=S=�d`�gmG��<T=u�g�pZ='�<A%�U!����<�u���I=F>�<Hbm<��
�Ƕ�<n�;�5I� �<<�>=.�<=�t=��%;}`B=F�.<J-T���@=`4j=�v&��0c�S>�;�c=R=S�����@�6�<'Q
�e�=�X������~�;	�=�:��ebq����Ra�<��4�[R=2)�����<ѧ�<
̦�m˪�:9�����zAq�Rc=�k��I�<8�<}S��M`�4�g<\=�n��/J���4�9�<��<NY�<�<0l<�5D��}�/��Ñ�<)��<��ۻ׏��	 �<�o���� <	�����g���=��
=��\<{_=���;Zb�)=Ɵu=S����,;=�w� �-=��Z��~�$��<��<=��+=��P�d�y<�e�*0\���=G�=kf���[=�ɵ�uR�����<�"�⦣���<mDk=nW]=V+
�b�7�bj*={����s^=�x�rCi<�=�H��X#�ۤ!=��q�\=7<Cg���j;����̼��*�J=7y��v\=L���~ҼH�=��;�yX=79N�R�=<���#�=Dc~��4����x{�Q .��ސ�[P��_�<��j<2���<��;�jK:�Y�o��<�4��k ={���Jϼ=:�<.�=�$�<{= �稛���f����ż�]�BQ�<�k���.=�,�<2�<��Y=�=8��<ܥ;+�<��U=>�E�x�"=	=Z>=�U:�0�<����<_
�<�F����:<�`���'�`�<Gb=��/�l�+=(�U�RU��|�W=�Pd<�����'�� .=g�l<]l����:��]=������I=��7=5�����L�|��k��<G&U=g�$��~(�=�0=�i=������3<LR ;��غ����D�oܓ<�א=� =&�<�XQ=8���݉�*��Bl=�0k����<oA+� ȓ<�]��:�b��r=*�<�/���;���<>3=�=�8M�uW&��x,<�[��O�<=��;s��;�v���IAG�"k=��k�c&=V͜��Z�5��|Q<������=��F��~�3�|<g�$�m��u����=9�x�$n=��ϼug��z������[=nr:�]u��%= �O�hN�<��μw�O=Hp�ײ�<_��<�꒼��2=!���9���<��!�C�==α�<�+)=v�໊c�X�=K�=�<�E<�1=��e�8��<%�c��Q^;GR�0%¼�5=�S/�wę<�f#=X���ֶ<!<��<�-ͼT��=�<�YF<u�	���O��<œ�<��Z��R�<x���w��%滾7O��c<��:��=f]]=)H=l��/��<~��=�����Cj�<C��8J9���Z�@����;�?m<!4�Îb�^�=(�b���T<��[<��<��k��}��"J�@r�<x1B�L=X=���<;��<u(�<9uK�}��<��=�!M��>�;�ͻ
 ���ɼ@H7����;r5żZ��<�@��x!��9\<�{ϼs�E<��n=���I=􀃼�j�;��A=�M�<g�I=����ē��<�$��_�#�eċ��Id=�/�=7�<�B��y����c�f=��=$BU�yc��=��==O��n[C���r���^=�һ�{*=�@@��9=Q��<�
\;4�w��P������:E�;=�/���������[�^=u�)=���<�O ����<9?�{�s=:�P=d+�9�=A�<�#=8=m0�<cS	<9�7�q��#�<5Z�<`�8�,�=�UF�"�w<WG3�H��N8��"z=�EQ=�i�2~ �x�;|=�Y�:[�<G�=Y�=��0�<#�ؑv:ٜE;�U�<\��L�=�B�=!nA=�w�]�;�=c��<�p��&��@��yi�<H�
<�2!=9\���̺?I=넊��(o�7���A=���c�_��\�p��ed=D��<�Ӯ;5�O����� ���Ƴ<픣<[A\�󛄼�*����<J^&��<i=��F�"'���	�g=k��:?g�:���`�׼��#�s�;�O����<<]S<NJL=�c���X�"�(�&#����:sT=�6�%.B=��=�����<�"=����%�;Fy"�����_H�4j�<)#<:q�-�ȼ����^�%=��2<V	�;����!��⵼�^W��h��Fr<%o��9���s���
��}I��T=�]7=�Y;=��M=1&��W�����"=%Aݼ=�<�FQ=͓��!y��b��<u�<G&=)��98���<����%=m�[<�o��)K&=Z���?�7�x-<]��<��7<Պ9=��6=�=���a���['C�	�����߼����@<���8��<n�ͼ��<�J�p�@�L��;?ƾ��`h�	͏<�F�zbo;W�<ib<�dN<1��<�����j���Ƽ�H:e���F������j2�ѻ�@H�=K�<?hE<amռOp�,W~��<{qL="�r��㘻G' ����<kV0�i���7��=oI<�=w;�&�;���<�=R<��O��K=C��pTa<�ے<�`=c9Q=��:�x=�T#=��<_��:�.�3���JV<�-=|��;5��Y!=�^'�H��$��;�?=;I{e=�#<�/.�h�+�Z�<�f��:<=��o����;�=�(h�j79��ɟ<=�Z���.=)�x<D�1��=��d��V<��=ɉ�<�����
6����<�N;�hM���<7�=�1�<ةq��7;�L��<��A��v��g��<e��<��)=��x�ګ<S6��~�=��H��ۧ;C.����8=��<:Xe=E߉<�gm����<����%�G=�GR��楹�
;h =�[�=��F=�R�=�t�6���lփ<���<Um'���:�Ċ�<��7��U���r< �=I=�a����<�6�<8��a�@��<�>��r�ׂ�YB�:o�%��`;��(r�<�,=�tW�V%�<�����=��˄�T�� <�;�d"=�B��$�<$�j���<x����<P=��򇬺T�<��:�M��;�>������Y=��<}^���Q�H�P= �
�S�ܼ�UĻ��N=�ɦ���:��k:B�ݼ�t�<��X�Nd��(A�)�X<;=����m9�1�=	���4�<�i໢�O<��ͺ�,[<�p��<=8��<[�<C�{�DU^:�b<�^~���1=�c��z=�'Z�4��<G/~=$� ���d�J��;˗_��~Y<+�/���<�t=��Q���;@l2�1�<�;�k�$n4�a/�;#J<+-=����`<�%=e�G��3�� �9���)�1�����<��
=0�4�ၼO;��Ȳ�9v�ͼ>�^���"=���꠼��<��h=�=��b��t�<�.?=�G�<��<�c���=�`2�MQ�<�AG���0������<a:�u�j��<��3@=��U;�V�<׋���"=0��<`dT<|h5<�g����<�,=,�Ч�;Wy��Ŀ��*�f�R���� �<�tͼ�y�<��0=
�<�aX��r=e�������<khx<�<><��8=?�]=�:��8=^k��%�;�������R����Ir<BN��Ekz��׼�<=l��,hu������h=�G�+�C��U=�[��CJ<񲂼@���7�(:(;�|����;��`;��~�o)=*�Y=2�K���^�?�Ⱥ�d;��I�<��;8?��S������<nO�;�`=��/Y�A�<I9�<�a����<;�D=�r�A�<N��<�8�<Z=�Q��0���V=x~~<W�];"�]={�G=E3�!��<�<!�<rb�=GN���'=wh�ܱǼ֊��kB��9t�V=Ҽ31���'=5�z;=��<7���U=��:=y�D���?=Q漦��<:�5�Q���Ɔ��*Ƽ/��:��"��	�<q^�==��<�,�!_=��l={,�;*\=�Z-��Z���+�V���O_=i��<eH���v�p���N=ɓ�Y�	=`�w̼=���wY�%�0��yN�#٭<���<��h=����bx�<�e��l�;��;�=�k=�X�x#�<��6�(�k"+<'�`�=��|=�V=�/�<�h�<t��f�=�e=�
=8�:Jo����<z��']�Z�<���;�%L��(I=_^�T3<o1���=�;���.Ѽ� L�ȆZ�:�,����<3Zg��d�<��v@�<χ}����<�$<��	�di8=�7˻qB-=u?�;?�g=�=��;����R����<�=)I�x��<��=��!����AR=�9p��N�"|g=�=F�;U�F=OrǼ`�U���@�a&
<�D=Epݼ�gL=�`-���:ٌ�I3j=��<>��*��+��:�<>�=�S�<�Ş�ߡ��C8)�x}�;L�<Q=nz�=�e[=\�<ky����=��C��ِ<��1=+��=ϗ���s&=��R���S��<=Fh���� D|��*���=r`�Q3=��,=/p�=Ũq��H��`��<_�<�SS=������=HGD��`�;p\�<b��:�OI�\]L<��=�QＱN�= 9=wnF=�~��׆(��M=����O"<x ��2bw<�쥼𰣽����D��;9�&=DY�<�Õ��2=J�c�+�<jƍ<b��_ � R�<(r�<�YI=�tM<'�=�UR;�P<���d+/�P]Ǽ=Y�8�<n�G�yQ=���i�;=P�8����!5s=fyؼ�ۼ�l��<�c���?=�:.VS=�z=q���^�=��0�<��B=��E���1��as�=�,Y=�^�Rü=���p��24=)�e�P�4�avo=�*������O=J=�2X�Cx�v�	=��A�|�7=��m=��>�9�6��j��G�<�ټ�|����ؼ�ES�����ap��!	��ۼo��<���
z���~<��ѻ�񟼺Y�<=���5��^%=!'���׼�$4=��d<icL<2����EH<�d=_).�Ď;/k�Gٻ�yb=e�¼�A�<�{������0P��^r����S��z8��ㅽE,�;�.=z~����g��2�=�4��,=a�'�&�g"=�':=�3L=Q )=>�}��=ji=u%˼�W��}s���B�u�	=�ǈ; �F�g��5�;��<H^k���#�^�1��U�{a=l���,��<�>��Α<�b8=oP�x�<re����=��F���<t�4:I�6��d=S��;�$��T<, ɼ;���_XI���!˂=��ۼ�	=m���0�=�Z���A�t@&<CE:*���lڼ���=F%�����Ο�6����Ǽ��C=�`K� IK<�u�=�6��2�i�"x2��9r���_�t����;u=��=�kI<�+=�u=�\K=+�)<^� <��<�l?��*��8A=���;�]��d���=읏�}�U=��0=8�9�� Ǻ^�n=6�P=���;4/=H�>= =�E�Z�<7==DG���[�l�R�H��؂<f\=��eS�W�<D̛<tP�<��K�Y-�<���2�_�E�<��.��Z|����<:v�<X4�<�F��B��"=Ρ<��A=�^J�Zms����.H=gh':ͣ�<]R�B|�<~㼯0���׼~6==�<�su=��/�Q���;��.׼$�Y=G�
���N=Cb��@=`|=� i<�f�:��<5>;\�ٻ|^���<��G��Ba�;��<�:�=�=��w���=��=`L��e��v/�"0Y=�4�=ڒL�&�8=��=��<z~[=\s�R.�7����c=ޕ�=T"ʼڽʻ��<�w �)Xp=�V=̣����<a������\=YW�<Bj޼N�\<{	���:\=�c#�"��:4\D<zc�<^�=|�`=�ڿ<T���9����+=���>��<x���5=�vV�si���=m<醂�U����p�<E=�f�����=�<��*=ݿ~���=����d\�-iA�N�<�ݏ<�nټ8ذ<�w9�|��by�0z��� м�J�T!��Z���};=>�o��N�;
�W�r�`��g=A�R���`=�(��H\=3��=����
ϝ<Tu=6�3=�]�����<}w=OH�<�K��ͯ<��^=,�N��c�<(⟼��r=�X<d��<&��;��$���˄?=��m�HP�2󻘿m��N<m��p=8�D�5������z=�A:=��;�<�<�������<���x�7=U��<�;����<����=tּ��A��,�;!�
<�M=�λ��I:c��������:<��X�G;#����H^��{t=;��+J4��o\=��~��:���;��M=�H=i.�5�{��Yؼȹ<:���;Ow<�eӼ��c���P��W�<��O<W�G�X2��ޭ"=K�v�w=7/=��8=��;'p���D��ʩ<>��`�;Y��<}��B�a�ȼE=�M�A�j��:<�/=�=7w�<V�=T=S�<�5���|���ȼ-�[��R=&	���}=˚�<|*Z�	9=y��<�]=��g��=�=9�<�FC;��R�q��<�<'��9���<遽��?��+)��!��߫�_r�<&1c=n��G�O�����==���S���#��Rc=ӓ.��d��"����L���ic=�<^n���FI���	=LRƼ�7-����٪<h"=A(=x=�&��33�B�g=R�<�;%��
T=��=b�;�d�=*���.�Z��U=/L+=&q
=n���??�wH�fG�la�jx<��=̷�<*n=u��<9�<�i��=N�C=9�+<M�`=���ЈG�E��<&
��V��;z�?���<�i��=���H����U���@#=��;�̟;����I�~8=��I�=��� =%�`
|=t�3=98,=F�<-�M=b�'<�c���`F=>�=�Gؼr><�BK=v@<�χ��e��1�=L����O��ky��E?=�JF<6�b�b�=��A=gx�n�-=kO,=R�=:S���r��N�)S=+4'=�[���+���=>a��'0Ż0��<��5�����r�'�Q��<g�3�=�<�����= D�:pR�<{Jb����ż|��9 /<p_B���Rq�u��<:Rﻖ�P���2<=�(=.+6�F��<��O�kL�Pw���	�4>l���><.�%=Bj�<���=�#
�"����0}=D'�[��<e��<eYż��<
�=�Ւ�Mr=��=���T=�<�Cy����ܿ4=�qa=�t=��<^s:=�=vC��)j;sF��[=X�=���<�hZ�4=`¬<�<�<F�<��ـ<���
@��s�=�n�$�+P�x$�+�9=	 ��<{.�Jr���_��>)�+|Ⱥ�`U���H=��<d�=��2���f��%�&�>���<0I=zo=�I�<ɡ�<�.k�q���=3=	-ƼzL�<+�/=�f��-kq=�oo=��J<�1H��8H<EV=P{�;�1�Ii���K��ȼ�\��Yû�W��Xf3=J�*�I2�+7�<O�p<-�S�l~}�A$5=�TY=J,���/<[q<=Y�<�A=;��<`q?��\V��-?��EM��4��ȼ�]��tB=2�L<�P@=�_=��6=��U��q$��J��� O=}�=���=���<i�<uM=�6�Xy�<��]�<�μd,;��,��}2=pk�<��;��"���iH���/�5�Ǽ�,i�;/�<���<X3�<XO��]E�;���;�̂=�JH=�HA=,�Ҽ��}�����&�1��c=u	v��=+<ÃԼ�Q�;?Z�<��(��$z=�S<u�p��e9=F�S=	0�����j�Q��zA=z�ټ��l=��(<��<�4���2�;�a=��=�p�&=lj=5E��R�;´���=+��;��D��r=e�@:�~���(c99�����=�Vs�<�< @���	<!�<�����@�/�9=�Z��؛���<��<\=��Ƽ؎�<���<}P�<aRa<��Ä��B�<%��;�c=#(�;2C�;�1:�zp¼��;�N�<�rS�N\J�ͻ�5$�;���Pd<y�.)�Bx^���ݼޢ�<{�!=Xb�<�;����<L��<l�*=4�?=0������;���<!;=��<�=Q�~{;t��;!��N=;����S����1(���=�b�<�X���=��E�E���$W�Nr	����<��]=���<��=n��<�����=� ��͗<T�[:�<l�ʼ�̇<.R�<oy*<�׻�[��V_7=W�2<y���)��-5>����<�r=���<�u���<ܾ���=��}��<:�,��B=ĸ�!V���g�<OO���$y<>2B=C�U=�7������=5=;��!<�r�<��.��	_=:%��f�=S��=�;:�ǲ;\k���Q9�9�OYݼq��<"#=`��:sC�k	U��E�<0������;�ޡ��J�usC;����\��"���M=ۘ��O�<��;7�s�Od���S;z�<��;mzE�O>��2oE�/�o��qܺ�e�<�=uI<��c<�{�<���a�0�9��?�Y�w�}�����=�����VB�RS��8���P�?��&=�qK=��}=���2Z�=��!���5;��^=�P����=���5%Z�������n�k�!=!i= d=㽼~�ٺ���<��9u%B�ʿ=w=�<M�<$�9�"�S=�p8�d�3�l��<2��;���<�K��d.<	�0=\+=���B�r�<��˼Eր;Λ��T!�<jtA���=gv8=������<>�	=_�L=W�7=ز�<�1���)=��@<��߼�y��$���夼?.~� �<N�F����<���� ����3</W=�����⬼���;S<?YA���B�@�ܼ�l���<?N!=v7=�*�<if=*=[���x���y�8��<����Q�<�B���5���)N�f�o=�;=^�=vO=N�<2�мD`�y'���p�d9=���6=����u��}<V��;�F�
D-�au&=L���x���<�ygG=~J=ٵ�<���B���T�V-�W��<��<Ky<�D�� 52=���3
��l��<�y���==�!r=R(�(�Q���$=
�9��d=�О�d�D�xI��{S�����=�
=&9=��Ļ��-��=�;�(=o�����<���nl�<z=��<�� =*D<�N�W��<�ȁ<��;����be=��[?�<�aӼ��:@�.=�==�l-<2)�QO<wK�~�5=G8��Z
��c<�����|��,,�=�r<Cs==>a��A����:u��<
#��r�<޼�<IK����ъZ��,��?K
<��H:�84;��̈:k�`�
�V=3W�<�b�<��<���b),=zA�<�=7?�<��1=�T=f1��#�h�0������k�V��,Iл��;E/x��=�<�<4�4<:�˼�_T���G�T�_=w�<,*�<m�=�'=b�$��k�<�\��Z �8A�1�ϼ�rq���D�i=~�}~�<j�=+��<�P{<��𼎥���=�DP<[�9=�,/=�So�SXq=紅=ꅁ��g}�ީ��Z�<�`�<�_�<�-_<Щ=� <�H<V�<�)^�ov��7O;K9��n/�:9̼"B-=�A�;/�B=�
8��=-�<4"f=�9���<����\�������}ܼ:V=D�X���<o�<&��qy.=���iL=z�?������-��2<�P�*$<�����+=3�f=�R=�Q�<�E=]�}=D\�aB�J =	�Y=�}y<���<����;h{<�&+�#?��j:n�=`0F=W�<�f��&4��������>}=�	�:���~W���ɼe^H�Х��SH=.xW�1�:��Ƽ+��<6]<��л�t��"=����ꏼ4�<���;6z����;�ȼvJ����<׀��%6=-_�����^ϻx`[=ۢm=@2p<��=Eg;��+<<���,A=5\=�a4=�9��1?(�~d#��|�=�>����;﫼�*<�=��=��ü���x%n�-���.�<@Al�S�;=�ե��{<=����爽;�=��%=VX=;IC�<����K��GX�<�t;I��<VX2=D���CF�>�e=1�.=M�7=�'&</[<���e���^V=7BD�
�n=ș�<��<S�@=�����k��A2=^l�;�g��=rft=!J#=Iȩ<(�Q��<��N꺻t=�^~�6�=� ��9<�<�SR@����<0��;�\(=����b=ԃ���<!����=D�w�YY�P�¼�Ǝ�0��<>[���ɵ����<]ܷ��dA�7�|��`.=%�kv)�,G�H��8W�<(�@�U<�����rh=޽#=��\����y7c;F�;|J,�	�=�v�<��]�R�#�C=L�=��<\1�;���<�������/��d1<����!]<ˢm=��$=�����O�1�];�P=����N=N��<��1���	�]=),мS�=_e���<=�a�=�2G�I��Z�M<�
l=��	;�G=6�l��
 =Ę��b�.v�5�N=���<�Ҧ���={�:������YŤ<���,�1�<�	�K��<r�\��b�j�<#ly<�dA=x��QR�#��� ���K��W}�3Jü�� =n��Er=���<�7<��	=�W��ʝ;�܁;Yg��bD�<Y��=��5�t��<�pV=��~<�D��t�O�Tؼ.�)��坽4�a<땰<�<��v�S����<3e"���=��N=
Y��kB�����?����Y��A0��K�nGv�oo<��i�߭����!=�Y6=HR��`���=���<Z#=M��; ���h=����;�=���Ӳ����<�ሼ4���gg���<x�g�0=��n��o�<EϼJD�x0�;q�<��
=,=\��<v=[�=���<\d�++���ż<G_��|�{��tm�֭h���<���<���
(C=��<s�
=�'o�Y����f����;w#=>����4�(=>ļO�<���<x�Z��������A��\�<�#�<�v��5=�*�=SD��,�;��|=�ǡ�$'R��4����d/=W͙<����(�<Vd�au���<L"����Ѽ�l��_�;��4<��'�A��`��EJ<����g
�<t�8�pHB�I�]���8<�� <P�麁g�<�`���<�;D4���=.˼*�n;��$�O�6�&=.�<μ�S�^F=C��b:���=/Ul�lb9<�B�<���<��<����=#\<h�<���<�OX<��=�L=,Vg=.��X=ǉ$<�(�b&x<O�"�y^n<�1C�/��L?���eD�,]=?_G�C�i������L= :B�<s�B=�Y�WX�U��<W$μݑ�<%��;<���(='��<�(a<w＋�=�Z~=��N=P�J=i���<^�;�<(�<�?=� ���=��A=1K<Ѿ��Ib=�h:��;ڲp�Ԕ[=�!*�1ûo�.=��g���l��8=8��<�mO=� �ʃ	�F��;�$=D�s����1`�=]�>=A����x��H�<�8=>c�}%z�+�(=v��=8�Q<P-=kv�O*?=镐<%�̻۲:�HCμ~Z�<U����ֺ�iP=��Z=�*;=�?1�0�<<8�;;]y;"�<���;�{= C߼d͆�eg��������e���,\��[�Bt2�ft��.�
=rd=��3��^=�������X��h��*=參�����[����<�����<��S<̑�<N��<sP�<9��<�ml<wwj=˝)=�C>=�=d+�%ȼ�b���<k+i=�?P��'�<]�=�B����,�Ty"=�W�;,6�pn����=����/E;l�P��Z���|���l=Q��<yѼ<��q�X�=w&���;�#��:wӮ<I�=���g�F<����J��n�<� W<ߨ=RxQ�����$c��[-=g�7=j�<Bc=�z�<��@=V^��7Cϼg?q��@�<�ڟ<Sn�������;	{�<�����_���t�i�<�Z!�mz
=g�8=C*���？R�;U�?�Cj޼�E=�NR=يn:3x��շ<��!�p�� �X<�b�<
܋��L���cb��:߼e3:=�%���=�����G�<.�^=ެ}���!=5Y�<�=�;�Z�JMD�#>���$=W�����<�~7=�ﶼ1�Y�#�l=��<�*�<X�s<��I����<¿��d�T�Ͷ<`� ��A)<ŷ�<qC=�nb=h]	����<+'M=2��<|�^=t�Y��̌<��1�&＾P`=_z��F^=c��<�
=	#=�y<5�����;?=�5��c@�/�p�޵�<���-��g�5=�A=)؃��`���k�;em�����;�BT=���<8z=8^Y�?f����e5<Q���6d=)4�<)a@�����|������<�(7������:����<=c���t=�C���c<�gS��y1=%�;3y=�A�<]Y�<��?=2��$Լ>�p�l��'.d�>�=���������<+yZ��I仑����~K��R�9I��%?'=.R���D׻	��;+}�<u���)�4=u��<�]a�#O5=dNļw-�<�no��J��Qռ�G< �ƼS� <��.=>`I=`~J=�ż}�=2p=j�2=�%=*ӄ:��_�T�#�Ag=^��<�ڼۘü09^���L��� =u��t�<�C��
�$�D���<��:������=��_=ʰ<k8�=�u=�;�<?5<@Z�<�[~;@��@E'�/6��yV\�"�=�s<�Aͼ�TF�_v��}_G���J�OKH�bw�<9�o���]�@#=�UȻ�*"=�E=k�4��C��ҝ����<Y���	d��F�c��<]Q��L.=<����~��x��<� 2�%D�;j4���9=�?�.�[=P%�|�����:4����s=Wø: �:=:��;��L=�%�<р���<$u�;�o=&��<��<i�м�l�{Za=�tI<V�B<1u�;��>=��<3pm=0pٺ�[=@�U�=!,=#��<�P]=��W�y)M��w=V�e=9�a=�f��"��g��w�g��<,,G=B�<9+����Z=)@=��=+|ʻ*���[=�D<�T编q�<���!!�Eb<����n��G),���=\(=�}=�M�;�Bd<3�����;�;��;NS���h�b���K�a=9�j=��"=16�<mI����$<vR�<K�=~�u<tri<������<8?=�9p�y�b��;��T=h7���V2<'U=�6G=�e!<�|V<�=�������M�;1!x=70�:8��<MѪ�s���፞�����	K����?8=M�e��h=�^ =K_�42#=x�F=Y�c��+��_�(���K<�8=��=T��<���<�
�<R��;pZ=g��;5��L��<#l*�L��9�AQ��k<������<I�%=�i<��?=�pS�C�2=ܡG��]:<� I�*�T=�M�<_ݓ�2JY�yJ}=�g=�+F���<tF=Տ*�I�S���( ��?��
����U
=�OL�ނ켴����Y�<��<��<�B=�#�+E�<6�'�=᥼�tf�( =��=�����5N$�ù=�|;�-���}�<���S��<��h� �5�'�%���	�Ph<#�&=�3;S� =G�0=D�^����<�p�<M<=�$`�	T�<4�y��x��iƼ��<��M�iqS= c�<��	����Ox�;��<�u�<�t)��x]=0�W�Q�I=� <�N2��py={8���W���=zBݼ���3{e=�Z���=�Un=}=�S������V� ���5<H52=�zT�1�����<�2H�쎼��N��u=���oh��?X��`"< �=ߏ����w���	�=�(Ҽ-ؼݑ�<a���漃1x�NK�<�=�R,=҂Ӽ��V=��{��󫼐Y����G=(�=o��<�d��j�<^�s����>c=���<<=�j���P�{��<��j�4�2�<�ȹK<=펳<�U&�8*=ޚ��e�_�������=�]<6==ir��sۂ=&-d=��0�dc�;�ܙ<.�Y:��������<=��	�M�c=O���2^K��d��Ċ�a�� ��;W?�����<8O<�(]90h�c>�Y�7;�g<DS�����v�i��<t,�ۖ�5�t�m�<���� ��<N6�`�F<m�<��#<�r|<���<�[�;�5�<��{�7Yx�Î�����P'l<�B伨�)����<��B���T��l�x�I=�ި;[�U��ꮼ��1��9�<��F��J¼jb`=B���$�� ��kD���/��D����{(<���8=>Q���ℼ0��,'�:�[=$Uݼ&��<��5�0�-�g�?A�<��<���]
���81��f���H=���u�Ǻs%�����w�����J�.���Ҽ��1�0;>=��^�+曼ɳ��9�"�b��A#=GE�������F��1\�0�8�nq+�`�4�a�>;�;��B�S��<��h %=C<��&<|����#��11�)6޺T�<ДA=7hb� t���D�J�i�pI�C=_�=)��è׼~�?���<!���:������::�	=�3q;ʑ���3��%�<)^e�� S=��ܻ	y=�,ܼ �W���8�t�%=C�/;�L�=����G<'=�{��=6)K=��=Q	d<����4#=t���
�u}q��&�<Z#2=��޼�=t�<��<Yq<�	�	�J=Ѧ=��=�Z�<�O��jû��5</�<�Cͼ"��F*=��<���<t�V=��<�w��𑐻P^~=wչ<�h��/��<�Y���؋�3P=��I�*� =��M;	��E_d<�k=��s<�rO=�s==�	�;�GH<<�D�<����(L �ھT��g�<�;=	$�;Y�$=!�"�x����I=o=S�6��p<��=ՙ����<�2A=�Ta��_�;?�%=�=���IJ���^��k�(��-�<�"=�+�<����w���<��7���1=]r�<�pߺ�-=�B7=�3��sR�wu�=�S�mQ�3��<ɻL�z�ټ��(=��{:�Y�<��кU<�<�,|=T�#=����u��3=�h=~i��cļ�^�!-�;֨�8ꑼ��ļ>��;ni+�^��7��<��N�[1=jK�׃L��Qκ�4=��R=�:=�'>���<<=6��Y\ =��;xs]�i� ;܄Z<�@{<�<n2*=��X<Y���ڸm=���<P�<_�=l՞<���l�w<#+)=�9<;��!=|�Q�U�3�`��J����/=�q¼$�ʼ�c�f�����@/�;�_�<Svּ��&��2�;���<�m�<��+�lCP��w=�4�<��<tl)�T�N;XC<Z�ݼ���� ؕ;.�=<��G=�{$��12=h�Z<�ǹ��V=fM=@��;�w�8-�:�q=X�����/=ؔ2�;�/sR=�Uv�,�����<븟<la�����o.=f��<^l�;����>�;�4_��	��kK�=�Eڼ��+�2���P;�4����%<��緉h<��K�qUݼZl=�F�<�)=�v*��Ҽm=U��;z\�����A��<6ͱ��^D��4h=��=�/9����&����IA�R��<��P=M�<؁	:�T�;�3�<M1�::����=W�	���
�^Z�<Qvb=D$Ⱥ��$���K=��=oƼ/.��8�S<s��Q�"���[;�k�<7�Q=�;R;�+)=�֪<^��������=S���.��`���M���1P���c���S�@Ug��.=9��:�L=n��<k�q���A�7�r��=�����W��!ʼE��<e�e��M='M
=5,�<��^�g�ؼĜ��L�'=�8�<���<�����,=�@�<���_����R�����=�q�����f=l���dcM�<K�fvμh�.�	HR=��O���<�>+=���; :��-�]��<ߛi=}�<�:������v�`=��g�<��M"="Ϲ���ݼT6=�ͼ�v?�}M�;�=^�=|Q��~=§�$ ���n=���LtA=��<�̼аμ�=V�u<�ա;�́����<�m�<�B������=M��<J�@�$8R���� J(=3|n����� ����x�=�`�<+/�hw����X=���<J�<��^��ߴ<�t=�O9�=�g�<��<l�C�V��;�;�=��޼  ��+��<$��<�@o<1��<�橼1ȼ���]�8;�M�V��<�(��ȕ�=��!��Wp��]�<}s,=����]<��A�-s��w�=�+=c2�<��<��7W�N���(����ݻZ:��Yd�����H_�<�㷼��ü�=�����(�S��< ��
���=/� ;�B;�@%������:I`q<[,!�GD�;S�\���;mB=�#8�0�F=�*I���;)��r�$�X��<Y1=��<��@<��<����Mu"��5$=t���x���]5=�Mk=�M2�|c9�LB=�J����;��}�-+���� =�*����<v9 =�Z�U=��-<����ɩ�R1�<|�#�&I�n.�f��<z���G�;�����~��=�x�u�K[���3�;�M����;珸��~5=��<m�U= �h�R��A�Y��@��ȵ׼�6�<0IͺA�L=��4��A[=M��=Q�<�=&�"=l�-�g#I�7'=B�P=pcR=e�r��*�6c?,������ �S^=�ż����D=����W���M��7z[��V�<��֍$�%t=��-=��R<+
��S^�S'=�B�_�=�b��e�(;�n�G��ֈ��{/=�@�<��=A����Լ<|~��s�9=�j=m�=��n�W��#�=���)��<Fm����<[k�<���<o��=oV��*=y<%�=(ɐ;,@#=�N���L��w=��Q=T89=h#�/On��ڶ�^�<�C������c�a=e=,
=g$�=in=�)O=K+Y��M`<"?_<pӞ�H��<T��̯�<�^�<�y��L)=����EA��]1�3�"��_���G�������u�K�Y���U��k2�*�x�K��:���<�!=a�Ż>X�<P�U=f=�p��}�;��J�LƑ= ���n��=��B�;�y��A=a��:�k�;���<	Pb�+l9=���59<�<�*C��x=YR0��X7=7��<��t���3<��<ļ����I=�"�;�,�9�s"=a�Y=�g�<O���t�L<�Z=�J�6pW�N�H��cP���(�f�ߺ�=
�;�~�<JAI��_�ʽ��;_���)�K=�Rn=���<lv����N=#2>������<d���C�P=n۪�Dy�<������i=V�<�r=�b��h7=-\�����J�-���9��<Řy� l}<�]=���<�O <{�=Ñ!��'U=�&�<���<&��uּ,==��<����k|���t�h��<�Z=�=�<}=��<�=����x�=1�=��]<���<L	=�4�<���,4)=->ʼ=c���Q�a襼.�����ȼ\�N=Qs=�W��`w<�.�S�鼙�P=-����,=�q8�v|;��=�lc�83;�	�}�<�{)=LYx<��V={�1<����ʓ��������py����<�������<�_ż�9f=�=��[�.�_�,����\�<�r��V�T�d�<[�X=�D�<Q�r�L@A=` Ӽ�un=!"=�� �S%�<�8=�k:� -���Q�<�d�;~�６1(�>��i=�;V����� ������.=t�ƼA�2��&
�	.�;!؋�>������ܴ^��)w=C���=��� ��5D���<[%�<j�;�~�����0�:۷�<��3��B@�7��<=L�;@U\��<��.=��V����<H=r����x�<�\p��#�<�<�i�kB=_�`<��)��2=�𐼯H=������mF=OP���Z��=��8�b&�����)�B���\=yB<R�</+�<�s�<�������{��U5�������V<��p��X�;yF�� ��ޭ��5c��
B����r=��=�s��#<�ފ����<��<��S<-2=`�N=��I��j�;_����R;���#��y����m<W�i��	f�=�[=�-�coF=��H)�D,�
'�"4�.�=y��<;�=U�"�1r@=+�h��gs��W��Qg<�ჽ��<~�%=�|������F=EQ�ػ7�Quغ�r=�\<K�=9@|=��=��L����qG��+f�k����߼m� �VA���R=��<=?>=�{
=a%3=��1��h)�����=[�*=�O=�Z׼��S�u�<�G�;�-�����F��R=8B=C�'���l���y=�;�<��1�6rr��W��ɯ=;���.O�<f�Լ���H�	=`�$����i��ٷ=�i:���;�6��Aặ�<����%?=ސ=�t1��=/A�;�z�����<�+����;h|F<���r�=k�<��k=�ѿ�3��<%u=��^�|���m*�˭�&] ��vL��x='9R�!X��oኻ�'=<
.����R=<�ڢ�<!ǆ�M�=�Y��<��`<@��;4q	��<�=�׸��<��GKg�6aV��M���<�(�!�k�A����;8t+���ü��D�o�(=�:
�V�W=wFt=ñ�/g ���I<=B<D����+��RW=�$-��x�<�ؼ�!=�D1=��;t�=Iv=�40<:�Y=ͣT��8=�S<�+����<%�W=Pr�y�Y��^J��mQ=��ż���{�u�ba=�lԻ�'��P�����;��B�U7]�@��<!����X��vZ��2@=�?�<�g@=���<��<z��e=�_N�A�9��Ou���<5�&=��¼�{<�=���<��;eY-�ϝ���<d���B	<�Y=��^=�|=O�;=��=sW���R�k=�M�;!�<�EA=�i�UQ���-�;�=�;��q=ZO%=��;�0Q=��<��� =p|s��
�� �<sA߼H�u<��<���<�B�<��#��1*�Z��u�=b�<)�V=+=[^���s�?��<1�-=\�J<�6�<��5�!����?�k�<�!Ȼ�͏<����*���Vh���漤�<X`��U�<h��F��<N�	�K;л�So=��0����	��=�F�cR�� CQ<P"]�E���d�˼�&<�B���▼':o~ʼ�y�<��=&��<��<�+Ӽ6�;��<�W�1Ɣ<�L�<s���E�L�<ZT;3�y�8�b44�gN�ݍ�</*��M@�<�d��17<0ˉ���o��K%���=�D �k�=�N'=�������t�9��|=t����W��������=]
��u��IPK<��3����:�O��<S��,H�lw�9�mz<��� !j=��=�OĻ#Z6=�aE�V�U��_�d�����<��)�agR=��<��l=f8Ѽ�	���<�eǻꋗ<Ylf���<�$�<M�;�u�=��5;9�s�#�;=��.��1 ���;�A� =�N���\���6�e��<��<z���q2�����A���9	�G�.=��j=�	�<f����_=R�Q=Mp����(=��M�ϼ�<���*����)����WRN=�=�=5�<=�B;=�B	��nM��+�$�<wC=��`�W�-<Qv=<�ݠ\�Z�
=>�ػz�:�����a��!ѻu�5�݋`=��
=}��<?�)��t5=?@�ǩ=�a�E�|��<ȗ*=�\�<~ˤ�|�q=�� ��\�8E�<E^���<�*c�z�<���=�i��c<��N��i'=\�<]����d� 2(��,����<=bܼ�z�<���Py/<�G=og=���<7�+��ʼ-�3=�r��<�<�`P��q��X��<|�$��	�<��>�d���=t��:��N<,�T=�*=}����d$<J.��#'/=�/�<�� ��E5�%e<</u;7����X軨�@����<`N=>E�<X� �x<��ǂ����<�k ��+A;v+��ӑ=]R�<EA���<2��0�<�F[=/�d=
�o=s1����)���S�w[�����r�[=`���UW����}=0F=V�<y��<0�<�<;3X=��8=�<��7=��6=�q�K;o��<�i =#G=��c=^�`�>��!�5=2Ph=`b�;#x= �1=w<�l��n�7�R��FR�'�%=BƋ��9��h�;0\=}^������'@��/今CO��埻���͆���#\�&��<�HӼ``=�^H<�o9O(=~��%hȼ�rS�.�缆�=�%6=<=w+�;���<ݟ�<�I�=�ܺ�q$n<�W�\3�;�&~:~1b����Z��;Go\=��<�9$���S�껜�Z=���<}k�NWH=��
�JN1�uP��^Y�FG<�<�_�HQQ���;���+
��L�����=��������<7�:�7%�_�F�#H6���=5��<�V7=D��<N�O===`�=}i<v�P��F9�/�*�=��=sP�!A��l��F�;��f=&лQ�=<Ƽ˨<���;>6k�թ=+SB���9�*���K�cu�U�:=2���$n�A=�۔��$^<�_<����(ϼ����q��;8���u�;)�b�&m����V=*觼�sj�Y3=�4=p=����|�O<���<��n=�V�=�P��-��@Q��=�<� ��
<H�I���<��R<����jg�<c�=
ڳ�n78��*"=7G�5W{��Iz�p�b�t)::�����˟�;��:�=���<\����W����<:�1=�V/=
M=�=�;Д�;�;[=iW=vD1=zN�=ü(^:="+�<��&�n�����<=��<w��?��DE��	s�0�a��-�<]>ʼ�0����<��6��4�<�̦<;�=�d�@=�k-����M�7=՚��!�� �ͻ��<����<�_�<3uu���I=�)n�jD�� ��<C6=hG}=�+��<T������0����b;��;x(�;�X=6�A�C���P[=<����8�#�ּ���.8=��='�޺���<�U@�|?&��x=`@ü��,�(�o�м��@���)��O^=���<�L=�\���Q��da<��a=- [�@F&=���=ݽ�<�\�3�'<L�=�V~<j��P����{=��0=�R-�g�1�=a��rR�+�Ǽ�<�5=^�¼s[���z��H�%=�4�=D�;,-=f5�@� ��'�;)@�:X����N�V��<��F���=�H =��e=;�<��>==/��Ż��"�l<��h=PB���=��廎	�yTA=�ܓ<ީs:eu;��;$M=�Ƽ�V������R<�<5=�<���<C�^�Y�6=��n����<3�;$�<UM��)����<�@=#�ļ��̻�؛<�D<3��<[�=��K�p�M=q��\<~�1;�e8�y45�ZR=�_:\C���h=T��<�ť��X;&�a<v�W=�9���<?��%=���<+�ػC�=�0=�VT���<=R�<F�-�e�<�";;,�;��	�3�}= ˕����;�)=�=��`=���:�r���:	����=~�; e;��i:d9��q=�� =��s��������_<���]����|�$-_�9Kg�D���!D���=�<y�*��ټ��)��2=���<$���'��l<@a=������<��'����m�����Ul�=�Լx＿-,��
=1����,��=xI��0�y�B�:�ʉ�a�*=ݰ��=�<�:�<0"�<���<�km�z�b<߾D<���8�I=1P��ч�@��I���=��ü�@�=X�C=F���z�|<@n���'�<п<ަ,�!���R8�=mڸ�A��;��D=�����e<0��&g=��;:5!�:j�����wS<9>&=��=#���;�>���o�?��X�׼�*��)�;T�=��X=�>+���R�E�����<�9�"���b�<`7���b�<[���p�<.�p�)�>��Z=Sv�9�N\�t�F���E�dV�\~i<9�Y<D <�P=>��&��x=�
�<�� �M2s<�z+�խ/�28"�$��UOp=�f�<��J���Z�R�o=�T�z$�`��<��=�L)<$'��]���Ԓ;A��z-(��组2=��N�[�<��� �ü(
�~�==70�p���ؼ���D>�<��u=�:�<�fB;�8<�]K��<�g���W�<��̼���3t��kJ�<��݆<��#�__q���9�LE�:̈;=L8=v�<0eB=��<����~\P���S�^=g��<W�F?�1������;Љ�4��^\�=`��My+���5=��"���<��B�^C��9��o�=9��;��<O�J��v=._=;����< �μ���?�<��5=w��<��=�<�ڐ=�)�	���&4=��u=Y昽7��<�|��-�<$�m�)?�a�a�f=T/��Ƽ��j=m[s��� =Y�;�&=�!�<��J��M ��uA<��+<��=�L�<+D�<��м{8;lW�=A�ٻ[�;��;��H=�[D�D �<�D�8�2="J.:5y2=�ʼ�O�;���<gX<)h&�eJ�6��m�<D?�*��d�<����P�;������=
�@�U�k�<��<uOA��*<���<W=̊|�Ĩȼ�we��8<	��h�=�m`��Ì�Y0���~=u�,��a�<-��,Z��}h<Y�<�4=>�	�����=t���8Fw�u�7=K�S�������O;D災\�C=7�`=��==8��<!v�^�U��F��M�u=?N��/�<��<!���p��n����
=f��<�>���2=(|Y�i�x���Ի�L;�gh��hT=!80�(z@;��<�ۻ;J�c�a���߷�[y����<�2�x��P(�4��i�P=��&=̺k=F�:=�d=�!<犥���&<�=(���Fs�����?�<���A=���r� �;�m�2=]�ռ��	=����;
=����	=8=�<�9㼟�~<�,W=���<�8d���*��L=<Ş;�� <D�]=�<m���{V�����)=���<�-N<�Bc��$�;3S�;o}[�Ǩ�;��H��sy�}3��=:<!���W@��=^�7<���<�6Y<rQ==�ڼ���<��=�.��c�(��鍼�S�<+\�=�?=h1%=�,�'/=�칣�/��	h��p=���w�5�̮�;0>���J��X�{�<8]��6�@��<�ی<�������=�)�<fsw��C���<��<��;9

�C[�.�黩 ~=.�F���N=����<�º�J�f��!�����;�nQ�UB�<�����Gf<At.�ҡ_;8�������|A< #�=��<�"=e"�<�PT=��6�9��<T8;~xV=���/=�aG<� =ˁ���n=�i=|�@<�[�J7,=@�<1|6=˩L=X�F=m6����z=YP�/�<�0/<��4=�D���j�9�����<,�X< ��<!��<��ފܼ}�0<*	���K��O+���<N|�YB��X�B<_M�:b�ϼ�h��e��t!=8�5��OV�+[��D&=�>��������E�q����a��{�<����r6=m	=��=��Ӽ =��N=$:x�k�I=�!<ʡ>���<Ν��
�׼�������&�4⛼[q����{:��p���ƻ�Q�<����eռv�j=��a�Z�?=�Pʼ��S��PN��5a�7p=�O�<��m���=�S:Py7�;>�<��<$�\��%���$=�䄼��O=
D�G�E=_q����a=&����D=�JF=��B<��P�[�<�<6=Գ<<$�`;��׻�qE��f���;��Ǽ���<F�¼P�8�_?V<x���=�@����<�~=0U�F0���	��,=Z�:��4����<���9"���C=�@�ϧU;QT�<��8�D=y�<�PS��
�<0��5��,!J���<0_@��?��Jי<�_�=&�Z�=3�C��Y{��N!=I@=��P=��&�5(��2x���L�<��l��
ݼ��Z=��0���<=Y��Ԩ=���OHϼ��i=�>f�LBD=�㒼mq=�TP�dP�����׽L��dz�+&=��[�
�ʼb�D�L+<�͆<zļSS\��G]<lOi<�ړ��d�!�<u���螕�ýz�uE���B���FO'�a�=M\��+�\=�<��� B�ٻ-=��< �<,�<X�`�n�;��?��� ��p>=�8�u4?�p���P��ת=D昽�R�<&+�<2H'��+=u�*���7<F�<=�(м��̼��<x5F�&K<"�f����
��i����Pu�Oe=Ba��L|=�t,=��c�s=�<��:����P��X��<|=�nj������=�A@�K�=�AX=�#��#ټ�փ=�c;ۡ�;���<��=�}M����	�9�L;
K���-=/'��*	=,
�;**C�I=B���9��c;�氺<��
�ϻ!�	ļ�Y:�<o&7�x�:j�%=��=���=$�[<�.�4=��׹�Qh�`r�<�;�rL=��={�G��1=����Uü
�<��:�^�;�xL=`�T<5Q=.�0�}�^SJ=f�<M����:<��<]ۈ<�K�<��L���,=����Q��<ʂt=R��4,�"F�<=#ü�h��'=�H��(�e�Fv�<`�<�h<���U��;�.���ܻi��:PŹ<�D���'�V�f�@~J��:Y=YdD<��;�i7��(=$,�<��ڼWӊ<\p��q=�We=k7м�4�<ʍD�\0�<�"=�B�����;��.<��=|�G���>�@4{��˸<��=^�<�e	=�D�<��m=�����*��P�"��-P�G׻(�-=��,<f���s<�P#=�3=�)����r=xL�<^q���s��WN=6��<2M�;�̣������ü;�O=�4	�򷇻�H��'�^�:��!F<��<*��<`������uG�<�-���V;7
F����;����� �Pw����;fF�V9O�M�\<�=����I<����H�ڻS�D�Q+�/p3����<Hc!�3�:=��	�� <�I�<5o��
�5�\=E�"�vܜ��n=�uF<#e<�^���E�<;�/0<�`��f�����.��=C%��ou(<eW�;�N,�W�K=l����+;)U�;�a�<q�g<�;�o����<��IG�1jX=�=?+V=����O��8E����<�FtV=����1���t�u�f<+�<ng:�߃=�3�<�e�;D��ـ�O���T�����R�=4�;4���b-
=V!�J�#=~��<�QR��!����;�Am|=�+��i�;��|P=��o=7��<&��Zv>;��.�s�H��̼4H�L��V��%F�kI3<G�q��7%����:m���m�D���.N�H�ʼ��<�S<�Yg�Dn�<��?=�1<�+E��{��V�L�1@��W�БI�h�e<eԝ<�[�<���:+Z-���M<<2.�:V'����?��(�	��0+=��<�?6<�e߻º:�:���w��;��&����	E��3�<�?=��;k#=��6<��,=�0F=n:=y��=�� �ȹ�4��;��W=�8���@=%=n%K;Vu�=�쉼^Ł��L�;/m�<3�[�7������Y�㼐�<c�^���M�1_~�N���V[��=r��)�<�~�<��mnR=�5;:��<)k�;{�=�z�z����=H̹�~%;�5���!�;�v�;y*=n}?������켇�5�w�;f�<��㼐�0=;��<�s��潼J�=0Iμ��Q����r��>缝����N���<$��<�J=�Һ}T��==�C�lb=�2:=�?����<����:<k7�`�A<�>����=��[=�Ar������<��璘<����sg	<��ؼҩ?=��<��<m$={�<U�C; oc<)5�t�j�+��0����F�M�i=s<�e��2�<:6�;�&<=��[���V=�&@�߃��e����8�]<=�3�����=f�N�����
t=�X�%�m��]=[�I=O��8=�䷻�I��:�����a<˼p�õI<<b�<ܫ�<`P�<���<�d���<�.��v��=���><=���<f��<L��<����=�\�<m��<�]�ʈ�;�G�:=䛼R�㼈��<� �:�k/;�h�����;ą<VWT=�Z/�Y�=�l�;o��<�%`�[� �wb�L���#=���<3肽�^:��-��ã<�?~=֒�<:�$�k%o��&�l
�;)���2=2��y`=�q���;$M=g�d;�8=�_F�Z\f�����б;� h=1<%�t�܄ֺi}��Ԣ� P�S��;&�<1ok���,�4ټv��<vo�XQ޼C��<�b
��5t=�3C�g��;���<�o�A�(=3%�:Ca8;��;[Z��S��<y	��J%����<�[=�Z���=�4=Xx�;�h��R�=�S�<�+J=�p=u�����T;t6�	��r�=A"�=+��;)��<0�_��e�N�2=��=R��<2�d<�7�:�W���<X��<=���=�(��J!F��ۼ���6 (�+=�O�LNP=�D����<\f�rm��?q�7$�p�<Hz�<4,�<i���t���c<L�#�\|���L<��L=NZ<�J�=;,:���Hn��G�!�k=�q1��'4=�=<�;='i�f�Z="]=O�L��Z��I�P���!=�'l=C�T<��ż��f��r=��n<^����@¼
����K�<�����a���c=A=N�Ժ��N=hLr=�ݥ<�t=���<��;r�)R��e�
�P��<�id:��:=?����;��>üx�k�\K=PҼdQ/;!_�<�yw�3}�<��>��N=<t{=�� ��V=��V=L#X�����Td���Ӽ�NR:h@=c�:G�<��r�����$#=��ܻe��]��<�h=ڄ�<�\�<�7�L$=���<�[��E=8߼^����-��Y�k(��G ��HI=s�J��P<:��<�P�<
����
s<�<�&=M��=/a�$�D<]��v=?�'<��9� ������f<�����(�:�oż`aV;&'�<|OD��7<O?=��f�g?=�=WP�<����J�i;��5=�3��O������4� =��»��=�,B�YDe=�<=�>��4�f�L�-&-<�j��Q==B�]=�4=/G�<�{1<��=�Һ�O)���:#7<U�I=^򻼩�����;/�3d�<S(�<��q=24���3��G\�S��IU}<�<�W����7����м�����<���b=fi2�~��:�|����;��~���\;�m�<����;[����#��<����ʻ��r�>�<.����ܼpo��ڝ<n@�;�k~�pC�<�ٛ=��;V>;�)U�qi#=�d=[�ݻ���+�Ѽ�w<ގB=fX@=��;�U=őZ=T�<<�ݼo"�<i�P:�C���_��^:�ѓ���;�ƙ�H{==u���6�G,=�'��>�,��tZ�<����м?H=��]�@Y�3rH=�H�;��=�Iļ	�<�_�<� o�;>�:�[{<��<1+�<+UA�e�'��;=�N6��#,=��<��<�Q�;Y�l��~���EK�T=
=�ڏ<�����?�9��+��㹻L6��=�=�AZ�VY#=��=��{<o���
�s���
��v'�)��<M^�;��<�n�<�7=у=efb=�
i=!��<�w�<X�Ѽ����-�=Ɂx�Y�>="��<�&=4>�;w����B�<��"���<5*=l^D<r=��Kc=�V�
�{<�7�����혺<���<���<t`!=�C�=��l������=q���c<:�ڼG�4��(=K����<�.����i��g�<�Ǥ��cD�~X����;�2�ѯ{<�nм�=��S=$k^<� �<��S���^����-��;$㖽����)<�J#����<�I#<K/1={m�����=����@�2�.���q�5�<��<��8��	R<b�Z=�L�<�S`�g�<=�sv�T�z=����V�5=q�%��Թ<&|o��1=�*�.�H=�I��� �!Q>=/�d��=��q<��ƻby5��"�<�=\CJ<q�C��CB��#�{]�<�?:=�45���'=(Q���ޏ�,��;N& ��:�97�<�����F�4� �Vxn���ry'���һR�4=U�}�U	���\e<i�l<�v=���T�Ϲ�X�>=M��=`��=n�/�S=�H=�a����<7?�<��&�x\3=���;h*�<��,�;W��O�<�
�;��!���L=r��<���<+%�f_�<J�?�!�p<�[C���*=�V�<wG�<��;�2Z8<aԓ�瑮�$΅��<��<��8��=3/�;أ�����Ѽ�!��a<v1/=�
=�	<�>�i�=����p=��*�4���=U�._�<,��=bQ=�?X<�6�<�y��
�^=�� =��W�е�2���bü i1����<N�=�l�<h�=�yM=���=,�I,=��=W|�#[h=��p���K<in0���E=��H<q|ڼ��(=L��믥���v��ȑ=�@��S<�һb��=f;�<0Î=H|�<n�K�����e<��m<&(�LV��1 Y��:b��a4��@6=`��<��m��C9�i"<|��<�d߼T�J�?.=��L��"=�=���U*=Q���,<�N>�ҕl=S�л�e"�]o�<�~<P �<��/��g�;r����i���,�o��x����v=.]ź��'=U���j��x��<t�{=�B5��=U_+=LV[;��w��\V<k�S= !=ъ�<+vs<�䅼�/J=|4J<�~�*�*��=��W��$Ҽ�ʼԝj=�B�Q#d��TL<ģ��q��<��:=���:��*��J=]+=Bo��a=�d.�V�<�f^<��V=�����V=y���U�$|�<����8��5|<��1��`9�5�<�OK�\%�<&S��G�K�g��ݽ<�v�;�� �||'= �~<�.����=!/�<"z���|�?�-���=��<q�}<��N�S�<���?+���"ּla���4���' =k�*�e�^��]�s�=2�#=P�c<�=�4=B	��{�H�b��<Z�{<��<�W��,&���ջ�yY���|���,�� �<Zl��RK�I�;�#�9��*��Z.��� �XK;355=��:e�-<2�=8=K�d��=�֔<���<�l=ʢ=��T�s7Q�*>�e�ۼ�f=�7��C��,m��H:��ܘ����<5��<]4`=i.G=W:;��)=<���g7�K�<=�s�<�ӓ;.��!=�4r<�=�<j\�C[�<��=�N��O+����v�E=�����<#C����/�jo�=�(��=���r�<N׎=�]��8+=߆�;,E�;���<)W=������(����~�r=�o�;75�JX<3R�<��/�X��<"B=��#=~��<:�=1����<�6�ЅW<���2�����=�=x�@UM=��T�V�=���1	H�|���J��;j;�M]���� ���<5��<�D� <<����U7�<��A=xْ<)���|�;*a�=���A3=s��;�CK=���+���G���L�<�μ�>:j?��Z����<�� ��O������5�œv���i=��a=��=3��f[��D�;�t4=6��:d==�1F�)*9��D=԰E<Q�?;��<3FP=iS����b0��r��3����I�;��=<j$}=d�=�%��6�F��<��$=I�<�o=R���k�d��`�;9Z�<�Q=�?M�C�	�b�|=�H��
�H���H#��W�=�_�=}��1����;���:�P�8O=��Q=깩���M<�cF<�k,�[�=��V�K��=�Ů��{*=k`�#�����I��]6=��o=�l���ɼ��,=��;V'�UA={=�I=�gA��?E=+xc���)��e�;��?=`�ͼ2,.��>�j,=|�D=/_=��=��K=��6��47��J.=���A
=�u����==��-�.��;PX��m>=h�,<z��퓑<��༖�4�cwּ�c=i�f<U��<H2��}�<�N~�YĴ����J��<�6&� Ps<�`���$<XS�4s��g�<\��������<�D=\
=i�*=@�<� <�y�<��޻��<�C=��|=׃(=G�[=���^�e=�W�<wI0�B�=�w==�Ớ��13�?&��z��6�
=�7�����B%<�߼�*9=���;3�4��;��})?�E%#=�A�<�Ud��C�F�<>a�<ҿ�qzp=E��_���vH�<���;'>�-:=��K��yT���<+�F=��<n��b���i����<�_�<X���p��B(<y9��=��=;����^bj<=����S<�)	�A���C���&=��,�,�<E�_;1����qw=//=?!W=��U����:R��})��%[���E=��e��f1���$�G��@Lc=��.)�<����ۓ�<
H"��L����*=�3]����;�뻃�4<�=F��:U~=6�.=��/Q'�#����+�U�V=UQ�ʟH=@s1=

G=��X�XP)=W@f=Y�S=N�=���ϻ��L��;���/�'���"<�_=&,&=አ=g��j	=��u�S��<i{�g�1ܤ<�U�a�K=@�&<�8�<��<̲���M=� ,��@/;	�&�C~{=@$������k��Eż����������L��<MMJ<�C=�R�< �=��8��<�ּ�~;�~�?=�C�������<��|<1�Y�!Jh���A�TAݼSKɺ/M<8�.�B�;t���&�#�<��(��<����wQ=��g=?�<g��<��@=�&�M9�=L�=����Ξ<��;=��X���������<�pм���M�E�/$�<wl�<ށ� ����V�2�"��{��^CD=
�<���<H��<�mH=�E�<P�F��s.�H={j��S��<Vw�<��=��<�} =���<�M�<��=�Y��J=yG=^�ȼ��;�k<FF�N9=f�97,W<C1�<g��<J�^�k��s5�;�7�<�l�<�e����<�RS=yȰ��|a�Z�L=�J<;4�=��';���<,f����=O�<��<�=N�r!@�5�9�ш<_��< Q=�*<����%F=qݼ�<I|:<Y���,�O=ߌC��?��L=l5�<�����J<=`�<��L��x���_=c�=�hR<SS=+)=W���0�<�o��\ϋ<��J��S=��;_#=^W�.���	=����՚�Oo?<��C=
W�<[5��uA=�d���T)=C��<.0}<�ͼ!���;�G|��/=1��<�L�-oo;}�W��Dl���<��H�9�6�oL��[&=�#=������'�6�;S#@��k�x��y����==D�������Z���_���e=x#J=0�=kDa=8�W�:�%�(�x�p����Nj=��A=�Eջ�q!�^�4<�)H=K!<uK���<{�A��2L�'�0�8I�sO�<Y�L=Sk=��>�`���ٍ<�P[=+�=I?�C�.�"3��
�;J<=,Q*���D���"=۪�:�j�}��<Y��<ӡ=�=Px�<�5j�I=z��<e=��<ƥͼ��)=��#=1��<�'(��Rּ�)��_<���+�U=�� ��T��;�o��!@=E���B=9Q��r5<��<vl<��{<�����+a=�4B=��<� �;Yhg=�7�:ͩ:�E<��Y�<i?-��<ڻD9�I��"K�R.8��s	=������;'[;�w<[K3=�C/<Xx��LL;e�!=YzP=�p����9��ET�^Pl;{�S�<��<�d<0�������6=��뺱޼H^żc]=�I�<��{�s�!=ʹ)��W�<���;� U=�m}�<�b=����)=I:�έn=u���$=�����S��<`��.༬Q�1<6e����T<�$��W�˼���j"=�Qb��~n<��q=�H$�=�ϼ|�h=r-=�\�<���<�נ;eK,=[)��?y��Q�I�="�弱����X<=�!�+�k�ޓ��6�V=lp�<:I��-g����\K.���6�݈_=D�$;D��/�=7,M=)6:=t=���7=q��;�/Z���J=U�<�k��[]=��,��#��<{\=�Yټ1�)��v=r?�:y��j�z<P,"��;o=��=r�q<�D=r,T��ڶ<fF=k�I�\]�<��=�7켍;c#<��~�e#8�����4=���<�=L)<��h=��I=���f:һLl<d�G=��<���E�z��b����"=�D?�OD�<�7=Yg=�Ng��T:!�=/��8=������]�v�;bG�\B�<#��; ���R��<�y�;2S�<�T���:��[Ƽ���,N�<D�<$c�<�< Ӈ��ֻ�8��9�㼖�|�kt<Ŏ<l @=n��:&�=�ɼ�Mu��h6=!a��;=|��<WqƼ����v�R��<�o�:(=���(�u���Ѽ�J=дʻ�;Y=��W�1.���<��5����b�j=��]<~�=@N����W����<�J"<3-<]bk=��"<�KӼ�K=h��c�*���w�����ϼ3�<��s�����g���J=�ZR=���<��"<��d=�d�<�EU=�s�<��a�Z���K�t:N��<���<$r=�\���`�����W�:�1�<J$�	�A=��%<�`�Ѐp<�=�K�<��<�\�
��<΢߼�ZQ��=_#׺r�X<vb��^_�<w�<>}�[.W=���<��;��-����<�hr=�y����{=V伡�F<Ri=�i�=	����^dʻ�U�k2�<l7=5�M=u���f���C=��I�>{�WԐ=e�<��a<��û.W��D ��=T=�E^��=Ά����N�
�<� �9�6 =?)-�`?�B�<N��p�
=�|V�V���0�ϼ�r����
=��~<��ݼ.�<V�$=�����J�M��J�j=�X;�t-"�T���=d�����q�NIs=ȁG<��_���y��<2.��E��<��!:! @��)<��!��0=�?-=#�J�/��Q�$=�'�V��F�9�x@=���<)4�	�X� �G��t��`��dD=h���n���W=TrY�R�;��{<5y�=�Pn�GC���m��yz)���?�U��;�Od=?j:=/�9���<��E�k���k߻a�p=� =n�꼲^Z=�P_��gx<H�<�q�<b�<,d���1�>l}��U�<���v%��M�(=��Ƽcw�<��<��x<��=_����bD��a�;FU,��'.��� <:Q=��ͼ7�q��{|:�!�c��*��<�e�<k�5=��o��b�<��&=}<o�=9Ιd��Ce=�<�7=����"B���꼠��<�Ѻ��@=e��<\�%="9T�E�=��R=��ļ&z-=MH|=-X�)�L<�LD<4 $=
S�;W��=��7={�i<����Xf=~Rż�eS��-b=�7=\��"�XC�=e�a=wz�<����-�<�U����	�B�<Iüh����dH=��ƺ�&�;YST=+)�cs�;�?=��9�\=d{����n�m�>=N��<�?\��2;�Ì�<�2����1"<ŕ-;��'<ܧ��\T�*�C�23���粼�R�⍲<>�1=�<�	=����� <��F�ֹ��������;=�X=�1�'7�<&A�<<��l�=(=A�;��D=̾ �50P�k�2<�P=�&2<��M�����o�_�=I@;_¦��JB�E.=�/�P�����*=��X���)=��{�7=!"&=�:�o�������<[�;<k���m���{g���;<�	��J�j�	1=�A���: Մ=�5=�L޼��g=8�<(����]�I���jO�l1D=���x�[<�i�lUw��c<�cX=�k.<�����pj�D�F��4<|v�����,X�T4��b���^=E���A��<E =� (=�����⻨݊��1=�X��l=��<(F6=qy��ݍ�<�f�<;)=��<=~=;]�;D��<w8�<�DJ�#3�Jg=��t;��켈�y<�<��E����ݼ��1�&R�=[>=�(ݼ c���{��!�P�}���?����!=��f��[��<�V=�rS�hbļ��R�Ѩ=*�=bË<�=1=<b[�?��<�Դ<��	=$:��%�!=k�O=�Y�<�E%=0�h=b��8����yd�xb���E�2�.���9:�1=m�o�[%h=�K�ъ�=�ْ=�v<[�Ǽ�0���"R���ü6XU=����&X�Q��-3��?h=Un)�+UX���<�|�;�.9���<0����<C�<���;1��3�<�Dr=��N=�=�<Y�(�X�j�
%��s2=6�q����<;ʻ��X=N�=׬�<��V���=�`�Me<�m����y��K	=�|<�f{<��1<%W;�Lj��:��(�=ٚ�;�3<��;qy'�'[��`D=ȿ`<�����pm=��S=\�ʼ��<;Mj;��J=�BX=M�̼�����	=:=/���bϱ9�v�	�>=D>;�b����}k��P �=d@j;���<R_?=� �s��<��B���;�RT���1��60��`<ax7����8�G�H���� �;��$�s%%��>t;"2=F���b.-�0���,4���Z��E?���+=;%/�~A��l<�O��,�=����S�<�=��w�r��<˾��}`E=?>�� c=޻?�����x<��=!�F��D�<�Ah���=�+6�վ�<�����޼�ӆ<��;Z�+��t�<��1�8�;�����;z�����h�+��D�<� �<^ǯ��K=.MA=�F@=�f��;T�;�N˼K�>��wY<���=8S�;��˻��;FsJ���f���O=_9�<BK<hѼ�h���:=�T����^�}F�=+���ɵ�C�󼠐�<*=�Ly�n/���=�������5=�ڻ�x9!=���G!��<E=!�K�i �<z��<���;�A߼�c=ij�C@�7�t-�<I�e=�o<��0>�"<���K=��A�oH���<��=��\�����2��A�3:�p*���;
��2�#��D)=��;=�Oü��
�ʎ<�B�;k/`=�ۻ����#������P�Y��/��-?�`!C=='=�6�W���O���;��׼�S,N�7h�����<���<׭=�"��<T��2?=D�D=�eX�r�U�d��X��<OxP�=|�;����:2��!�ؗ8�";��;|�߼a"���	<����J]<:�l���<��+;<1z-<D����3���a=��j=�ڎ<.�=^Ф����NpF=��<�=(;^E�S��:5���O��<�N8���<�A�<��=K0u���L��H;=Q��<Kߕ�+��P��������<��=ײU���׺�p=$��-�x<�oG�8���Á���c�����{pe=Cg��]#���Z�Y8��Of���0$<�ہ����<(¹��S=)�>��.���Ϣ��{=�!<v�:1)H;��ɼw伙�"�4��<Ql�<���;d�C�[H1=b��EXr;>�;n��<n\t=��c=1�/�Y,ż�C��v��j�9�6�<�����<J=�<�~���n�R!<��Yܼt�*<e�� �U��G9�X�<Ssq<a�)<mY[�ێ�l��<�1ϼ[uλ�{K=es�<QRJ=A/�:؃��e�0V�<�ܳ<\����$��C;�Zg;dS=�ޅ�Hh�<����H=}�\;�EӼ�k��B���4��|�<�>�;�Y3���߻��̼���/
=n���pj:T��<%�=����7��;���%�*���R��L��/�����<xe�<*��=��<�;'�׼�]#=U��6�;��\=��h�m��;�X�<o�V=�?�<mw�5�`:BK=�6��'�<ꤱ<��{��]�|��;/Y1�8��	�x�7�#<
�x�9mJ�ً<	�m�{	=�Ph=e$��
Ѱ�\j�<G|9��7��@�<8�(��H�A5�<����2�j�\z	�]α<�x��/T�I�_�2=k�a=�?k�@˸<�Z�z<�������<Ȟ3�H�>=s�=��=)�x=4Z<�H��ʀ�2n�;��=�ϼ7ּ\`������	��BKe=&�=U�JU2�!�==���;s�=�z�<NP<�1$=�F=5�<��<���Dzn�{L�<�eT�tB=a$�<),6==
���v��)=�[��,_Y�w�G�q3$=�#=K��j��<;K�<_1:������<'���]=���<�Uӻ��~=��z�ˆ�<�=n%���[��i��Η{=
{߼�R=��0�lQ2�u�6��"5�Ju����;��2��k�4N=2��;]���QF���A=Ð;��=�@;��E� �;RX#�Dҿ���ܼ&/R�P=�����9���E=�V?<)^$=;�L=��&�ve꼹1�x0=�s�<��j�,=x�=�"���g����J9Y�:���<�8B�'�λC,�<Jmһ��<�\�<en�=-(��3f=�Q�;c#?<]ʻ۫B�RR�<����d;�=��x=��A=[�K��ZE�-���d.m<� ��M�:	=�L��4�/�3�=6W�H�O�9?p=%�0��<_��<}���}~���5�_��<�>�
࿼#�ἸI�RtJ=fs;O���H7�\UX����n�d��?<��E=`|&�ke8<�R�<�\T<̦Z�z?b�@."��웼�м�N�� <��żRb9=�I�t4��T���kp=�0&=48Q=�=�<�\�<�	=@�	����<*{^;=��	�}&�;�~-�>!T=a����*�H�=�/<��
=�7�<:E��ėL<%��<�kP�t+����;��D=1]=6��K==mNe=��=^G�<o��<�#,<�'=ku'=��*<���<�ջ)�<���<�)�
�;6C�<Mzݼ$2=t;,=q�W������n3��L=�)#�Z���J{���ἒ�8���F��B@=WS��9�*=�����T>�/*3=�?P<�2Z�qR=�Mj=[0= QZ�M�&��n=Q�P� ���\�;H׿<�t��7�<��ܼ򊣼��T�f���)�9�@.=�����E��5�����Ve�s�s�x+=���^����;��"<W=Aω���w����<�D5<��C��_1=+������
d� 6<��O����̼�N;Je�>k=��ּ֬�<r�
��:�?�Q<Og��@��:�c =ɫ�=��\��[=OM���F�&A=���t���!c���3�,=�\=��=O+]��="�4��g8��-:��#�t=�6<HH�<4�<lT�;J������\���fK=Tü�:��Z�/�<2- �J�< r+<�ek=�cP=�"�<�ꁼ�0��� _=Y�I=ӥ�;���v�=�����{���@=��9���<���C��<������<��V;$���A=9:=����]I�w׈��ۻalt<ꤻ;�@��hv��.&=KO�ƙ6���*��_�<�lܼ�g�[�<~]���#��sּ�x��W�<V���9��<D�1�r;�I=sv=r�<��j=��)=b}��w_=���{����d;Da"=�wt<*=(��g���>�;�漳\;w#�4��:�u��'jA���!/<f�-=�0C�H�<�LU<D�v���=�W�hdE=�J1===�ü��eUT�*Jh�Z1=�A�V�_���(<�����j;��<K���Յ<��<�[ <y�1�YZ����<w�3�s2ɼL��<y�)�{��<�x�9L}���=�Ё���<\��<�ϼ�?=��;�W�V�<ոb�V����p �����;<��c<�J�;kZl<�4R�Ԙܼ-eJ�JF:<1�<��/�"�^�.�<Nh[�5x�4����=G�,�&�x�
�`�<[>=�[��g+���(;\�����<gK=�]ͺ&����-=xr��y���`=B�F� [A���i�@��<�8z=F�h<�y�s��i
�<�e��5��Į=������L�q��ī�;ْ ���k�=l��;�<H=� =�X�|�|=l��<PzT�;�[z	;26Q�E;�ܑ �Ϛ<[�<�G��O��l=8�=r�<��=��y=}@B���/=�Tm���=��<���<@;+(����s= ?�o|3=�� =j��<2���� ���w<VR=K�(=���<P�w<휑����<$�Һ�]=:)6<V)��vż��:����}+g=בp�y�<�D<'���;=��3��/O��Gj�����w�e��P=쁼�����w��խ<�=��=2�W<��_<���X�o��Ed=��E���8���=�&�v<�� ��{d<yP�<�]��~L=\ `���k<�7�=�ٻ,�<��ʀ;�49�h9Z�u��LR���6�<���d������-�C����R�<���~3��� �]I3��z0���=V�=8�bZ<d�=zܫ;�"4=o����P��n�ȼg1<:n'n���z�q�K������6�F�:=)��<^�E�t4�;�
=�������Cu��� �n��:�6=�4�<�ټ� �<�h�{P���`�(]P�|��5໲%8��8���"����e=YgZ�Tn��ݴ4=n��<��R<,d�<��;b���ջ~�|<��Z=�*ջnc�L� =��<���;�����E=(�;td�g���=�:��<�d;��P/=$0��@=�4˼�5��iͼ����0t�=�=p,�<l���9<�ad��u�<u���μ�;�<�"{=$"ռ�a=)~����<��̼\�e=��g��~R=�L=ъQ�1�=�DS=�몼�#ϻ|_��q*!=.dZ��h*=g����D�Z@��e$
�+d3��!�Rz`=t�<IS�<��»�4_�?A;�g��Q��<���<K��kBE�
5��U�!�#M<��=�5=D3�=��*<c��<VA��_��$ <����M=��6;��;
]����A�nSj�\��[�F�d�y�Fz�Q =D=b�@�!�0=��g��p�l�c=]v'= ���Y=W�����<���</��ƈƼ��	=3�l�?%=<��A=�e���G��^5�x�Y=����Q��PV<���<�%`=����p��:�ܲ���=�-�Q|�\����y�dOn��~�;�?=�k^=��;|=�_"�9c>=DwX�i�<�vܻ�81=i�=�;�;�)ʻ��.�i5�;&�<g���ؓ��:E�VdO��=#��O��<�jY�~�=6կ;چ��e����a�<=�����x;�ݯ<"�K���y=�<! ��YH=Ò���T�<1�W�.KF9
�>=�Q�<��^�[�c�E�-��-�< 0K�����@�#�M�N��<�E�|`H����<(L�X*�H���-�̼';s�3��6<2�<�T��䵼���V<3��<�<���_�=���;͙̼"����c=԰3�n�9=eI�:�'��p�Q=tU ���U���<���
B�<ό��͉e���;�~w���ϼ%��R�?=*�=�a�ʜ���+=P�=�OO�/v���CT�S?i���C=6K=P�<�����=�`=Ph5=�B�(d=l?g�o{h<��=�cb<:��<AeS���l;�Լ���o{��<فd�� =-�h<��=����!%����;C�A=�/p=��(���g�{�,�[� =�ɇ�z�<���ao����F�ݳX�t='ֻ�L �s�<i�����R��p�Os�=�V��GL]���1<��R=R�I<G
�<�[X=i�<�=��=���<j��<J��<�ӄ<�S�<�
@=��[���a<%92<��=��G=�D�w(U��<�`Q:�tƼ�>o�^&I�r�=aRC<�h3=�1=M��e�����$���޼R�`��=��=d^K�U��e�*�m�B�e�<�;a���<�`�;3QҼ�<�9�]�;��A�?ؼMv9=��d������D=�"=ߵ˼&H.=
.{=��*������v=���=�MǼ�7N<�I�;�K�<�p$=gG���;L,u�F�=�L�<�=Y�.�s�Լ�^��i=���<~�3���s�4*� vl=9�=�G���<0�f=Un=_�=�� �
�.=E7�/Ԉ=UJ4�� =�A;�gǼ9`@=�3,�$G��aL6��7��X�=�H���,F�8JD=���<��<�뵼o0�<WJO=��9�2=�t�l�<�z	<b�P=��P=���<ey����<��%�R����X/=O��<�����-!������;*�<�V	�a;=����<�2��,Z�:��F�n@�<�p=���wՒ="�=6a2��Uh=��=@	;�y}�:np=Z,�<M�T=/��U�̼x�Z;�8=��%;:K�<Rc����<U=�Y-=��p���ۼ?O;=\R<�2��_�;���<��C=]>����=t�U����QiO=�Z�<�96<=�=��C=&$=�R=;���;��N���ռ�S;X���k^o<�=�<"�üi�ټ����;1�������0=4<�l��=<i��#���B���f�B=Q�=K�� �t=�`7���������ܼX��<��P�6����
�������\=5y=]����C&=�mx=	v�폃���6=#��E�	=�%?��顼F
=���<�Ƭ���<_�=`E�|-M=[�s�-s��:=p�L=�3���7���<�u��,�m�^�ຣ�&�O℻Q8a�F��<�u"�B�=�掽�Eo=ã�ao[<� �����L���+=H֪��b�j�=��;���0�!=��C=�c�K�R�7�່���֑�<z�C�A�C=F�<�{�n2��.�����<�4ż��<�~�<]0�8R���[���	��b��y���R����g��#��-4�o�M;��8�S�<��<h��L�;�=(���:-��<��=�J��;5��P=�W-=ո����!<+D�;u�<��>;�CB<�h5=�SB=�̚���7�s` ��4P=�r{<��='Ω�*��<���I�,=��;<��f�fʼ�i���ͼ"��<Ú�=/�p��|켣YQ=�u=�Ͻ;Bao�d�Z�p�;��=�v9�?H=ANϼi��<���qX�}�<�T$��	F���j:¸~=����J�{E%<�錼Sj����,=E$�<��&=e�����}�r��=��u=�
м7���U��h��<���<�i�cBP<rϜ<4�`= -�<�(5�}p
�X���,=��	���g��<�t;�Ι�4�A��Z�<���;�BC�J�$��\��#��;�6�;�S=��@�&=4�K���<��-�K�L=u�T=&��!�μk�.��+�G�,=0��<3Y�<�N��dԼ���>�2��O��QR=&�I=�~��=dT=l����d�U�4�^�><[�^����O8���$����<b�n;�>���Y=�ʹ�;�<a�]�^�=�;8�&h<�8a=���;�Z=G�<h��<A=�6�s�*�Տļ{C=w��<@�����\:�8!�q�;a�Z=K�ۼ�w,=���<�2J�N6 =ə�<�Ɲ<*�?�)=໴gD:o�@��xIջܻ������d[�<{#F��$����A<�����4<�����<�F7��n=�C��j�<vt=�K�<.е9X[��H=��&:K��{�;\8�S�L=�t*;In0<�0ڼ<�=5��<��>���9=|����x��<��<��1�;�Q���<�(\;���uӈ<�r�̡=�҉<:0���~��&��<^�n=ܵ<P���b��w�����V˼���;�s�˜�������W=�z�=��q��ʦ;���;�:;ye<�_-�b6 ��o����!;��C�0pԼ�*E����X�f;N�	<�; ��<��F=��<(r�2^=�D�5=wVQ�l��<�8 ���T=�j<rۘ���<ɮ,=��B������S=;J����`"��_K�j��@X=kX�̕�<��2����;fr=�=��<�G��hJ<��w<	g�y�H=�$=�+=��:�,�����~���+�ߑ[<h�������YX=yC�[s���W<��<=Q�9��/�:�<�+���ϻ_�8�[���������j=�<�J=a8�sQ%�Nv�<�B=���<b3�X3�<5nC=�i=`�R���X�a=�a5�D&"�ر=ޑ"=�x���6�#�����8=�"�<�^���<����T�!���ɻ.��<��̼�N%=
�`�m.�:����UZ�;�>=�y	�%��=g���DF��~X�Jǁ;	 ���!=�Ka=�qu<�V����<�q<��&�DzB�d����F��t�7=��\=�p��s�;��
<� T<YA=�b<�x;;g߼�y���\=xI`�X攼jB�<�S�h`˼Q@<�� =�_{=���<~Ȟ<�x�}�<[{���=3�<�`�����<aW�����wP�R���	��(%S=�&j=��<���'5����r�<Op��!>�9k=�K@=���9��w���'���Q�
D]<i,<�^\<0��;��<���<��^< ��<�<�=2ڹ\u���O/��?�a�'=����w�
<��J<T��<�['����<Y�������;�kn���<�A[���0��j <ꦼ����E=��?�=�bP=mt�uu,�5�׼d��O��}�7<r<�H
�9�１DN=�Y�NX�<���)���%��\��/'=�l��J���T<n�)�����1<Į��:"�<~˷:A�E=�2<07<�=�T�8��<�X<4$=�2��� =���N"+�]�{���s��`|<�T`;;S����==r���In<Cp-�t�=�iR����;ê:�^Q[=�3��h={8=��V=�_Q���*=�q �UEI�Xzʼo�<\&�J�9�L��</?R=�p���ޥ;��6�q�"�)o8��}����S��d���&�4޼u;�<��߼���Ш>=�yS��ݚ��sY�
�D�T"N�uW<��%+��]t�1��Ma��a0;�0=�k�$��:ZSs=�ȣ<D�N=(��<�+};�&J��lP=��<��n��;�tb=�;k��Z�0(:=P�P=�zl=J��X���p��<�/�l���"��1p=��Ǽ�)=����zq�����E����=8h�^��<�w=v�=�"�<z#��~<hl6=�\^<[c�;(�<K��<��<���<������;~�Y�jO=��G�m��<|�;�!X<��#=� Z����G���*;[�@�[���	/��m��]=˦��qu�F=�;|<�Ƽ�.����*���z��j0=��:@n���@<��������4�[����KX���6=$/;�J�:�S�,�6<�h7��3�<n}=}�m�<xav=�;�@i`<�<��&=0"���=<�|_;2��0ʰ<��.=0�n<�=X=��P<q?�9O�
<^�@� r�}(<J����2�'`T=��
=�=�^�l�=��<v6^��L4=XGW�{R���<GS7�!�;�n�<�߼?Td��$2�8��=Ay�<��2=+��<��6=�$�*�<�y{<�[K�{�J=�<Q� ��\�<�lo�����0�l���=�=%=�4=��(=Ɛ߼�j=\$������cd�}�<H�;��=F�T��u���k=�P��]�:<r�s=o�]�0>��!/!=� �e�:|u��D���&<A�<�
=�=�$$��r=�&=�$��T����<s/�<��<=[X�<(�<u$Y��*�<�=r��2�o��E�����*;���I=>2�<�ѯ<��܃��5d��Kr�hc.��%"������mX�	�W=8ZE="ƅ����<M6��Œ2�G���=�_�d�<�xg�:t�=՟��X9�Ĭ9��H�<$=�^=�}O;M!��a)<K~!�5���~7!�o�=%�
������M=��z�Z<�,��|��/?6������J�[�=qN!=d����;�TD���;��-=�>6=H���u�y=��G�D���4��,=��n=dO��?=>�<�\f�W�6�!�y<�8�;��=�}^��I�<\��5s=�9�t�k��<���%n9<�X1=�BN=ó=�J=d8=�{�<Q����bf��;p�;��M���2���=�@�=/�Y�@������L�L#=��g=�۫<���<�=A9׼UT=N�����=��=����PT=kF=:��{<=}�XD=��һ�=��,���l=�@<�T=Ҽ�ռ5�=9u�<�|4�m�x�\�:nV���2�°��?S=N�=Һ�<@�q<�A=J����#�<AϚ�{�j��ڼ<G�f=?�����G���;�#�<�d��L"=lr�֨<=jK=���/ּ��n���;�/�^��h=E,=okb=��<S��=A^��ǚ�m���ļ �;�U=��Y��}D�X1�-2��	,='��<z2��η�b2�����,H���@<��];�����d���=�C{=&=�
|;fF��	%�<@�
=�^��s�:�\�=��2=��$�X�^=9;;�Bc=�|ļ'�<]=Ī1=N���0��j���8k���<��5=�U�<9[�8F)�qI:=·A��}�<�r��s�R���^<K�<W�=�?ؼ� ~=����i֣<�!`<�ʼ$,;=q{�����<W������<�f=#�N=}�(=�GA��V:�6��=�:<w`�<%��<�1O=� �澴<}��D�0=󼱼ɒ���¼>��<jv�I:=�<�<�#��!7�;-�Y�����ؼfg=��K�p�-;}�#=��<���<(~���P�>�,=�\j�>��<W#=Ń���DB�����m=���u��<�x�;�}i��?;= )��.�<,˲�-�T���Z���H=��{�(�E=$}׼�ۖ���<Ł;��^&=�;�OM=ϐ���f�}�H�#�Z��1W�yg�����&D��4�<�<N���<=	=X�<_�l=6�3=�6����:�(�=:j=
��;pEE�#�<�*�<͐j���#��_O<��=ZF����F;�FV��L=�#$=uЀ=vD=�3=:e���߷<�V=�q=��м��=�һYV�<o���'�V�<�J�<��0=�//��+\�qۼJx=c�
�M0$�� ;�dN=9�һv�<��J�gl=ʃ�<�P=1�$=e����~�=���Q�<�'=`�:�K�<5�<P�2���=x�M�4��=ȳ�w'W=J�����<1�K=�h@<8/��=�ѣ<&�J��G�<g��<[��<Q0=Rس:�>�;�q�ֺ����g��6�<"Y�<�c��^���<P�y�g�|�Y=\mȼ��8=�,��T�X�2��+��\�7�^t=����������<��=)#�<�q.�\8=6^<;P6=��;�!�����<R��7i|"��e<[����q���K��<�<=�h1=|�<޵¼{��I����ԼȖ<��b=�3��u=_��.^�<���:_݂��XV=�s#����<,)�<>��w=�ʼ�~���U(��l,=hM��"=��)9A2+<M��4�<;p�P�	=R
!;��Y��#?=J�����*z��)�Q;�qy=X�-�;=�Y����o=���<w�;�(=))v< �l�>�O=���:񓓹n8�<�!�?z��.�E�N��!�\�(=+��;�5;Y�<X�B=/:�E�=�F����o;(=�<"R:�i.��NG���@=	ʼr�ۼ[O�<N=�@�<���Ux�=���;G=-s�<���<_�
�j�D��hp<�rb<�0���8�`��<�P=<?�D=�¼4矼0�D=�h��l(���^�_"�<L<���@�<'�:��"��,���b���#��ռS��AS)=���p#����7JH����E=�v6��'=��޼%2=�Az;<,�<0ȁ=�f(=�K�?v�<Ä�;�E��T<8Ĭ�nm�(-�;��@<DA���s8<W�>=aq/=��X<)R=�>�<%z�6=�<���@����=K�;�p ���=˧��� <ȫ��&7��z\=R:�<��z�S��ҀüDEZ����<_�7=���<��	�}�t<V^=%H<Zc=A%H��\#���<:�O�����n1'��X=ш\=TO��
�k3����1� ��ɼ^`!<�jC��3��� ���E��s=��C=��;�!<��I���^=�B��g�H=�EO=��+�!v<���<|Ch�]U�����1
S<(=�����Η�T��W0=-�:�����h�<��,=����z=2q9=����<΂[=y]�=o��<��$��������o�;��q<*+��,~���ּ�S#�X��p���&<7(6= I�X�
=�!=g�<��<�,=���<��N=b�ȼX�n����΍���<2��A�C=��<��6=����9s<���=5E��eb=簾�K!S����<�<�<u�j<�H<"�˼�.�;u�ֻ]Oi��ǀ�T�+����;}�2���8��9�<ۓ�=3:o<mht�@��<��:�������i���W;��<�'=�JA�	�#=j@=z�<YS;��6�DRc=#��8��A=�j�0���ʺ1=Ј!=N�=��i<��N=�FѼ>ZE=+(.=exϼ[Ө<�^�Q@=ި���X�"T|<G�c<i+ۻ�;�����<,�=[n=Q�.=AQ�<�P=��.=,ӟ�J,>=)j<�9J�<$l=�|L<�X=�-=x@��A^�_��<�j�<� ��9= 8C�PJ���n=@�g=+}�;�L=���ȉa��ߢ<@w�<CS!��-2��6�<w=���Af�@P]�a_)<�_ünLü�U ��ڻw���V"�ʸ0=� d;#q=�/;��5�3���idD=Ql�<t��<�ץ;��,=��:��$����;j����<��=���<��4�<}/<5�6=�;�e<2v޼N^W���뼽t��w�<��j<��i��;�<e�Ӻ���:։�<��K�;�	��3�<I�=sZ<~�L=�s���%-�عq=�f�<��<��O��>b=�ko�` ��M4�z�<h��<��u=b_=]v��V4C���b�	t�
�޻�;�<)�|<Xv����><؆�;���<��v���)=t�	<o𞹞v��$;ntQ=��<t˶���@��Q���h8��%"=�_
��.�4�J���1]��~=��h<�@= �N�a=�82=��8�vա�&W�<ʇ����E<�E?=Ǵ�;�F��=��\<LS3<� ��_(���(;oC�S'�W�U=��<�%)�xs\��cP��c��y=�F��Zc3=��E�I=e�<��ѼVwV����ƶ ���p�Ϫ;�¼r 5=�o<Y?�<�O>��6���o��%����1=G{<��<�C�����:'ȼX}��L��`ԻX�+<��f���<���U<��\��2+���N=����9��<g=y��;�aм�'���P=�N�]��;{l!=_�=%r <��~�턇�ﮔ<	�[=:'��������=+�<=�=弊#�<n�<(}����F=(��jS7��դ�,�v�{��J-�������P�v�D�1Q�<�y�<P�<�2��ױ$�G(����"=}R:=O�=4
Q<y�4�b�==Y�"��M/��ɼ0���ź��h�y�}<d�<�p6��٩��ޏ<��<�y�<I
=QM2=�K�<�*Y����<�i��<���vs=^�>=�|Y�!@���?<M�<C#�<��q=�3�%�f��;֐|=��� ,i�\�<����D��<D��/��;0-<tȃ�G�M=e���WS;��9=���<�_"= "�<�x�� ��<�J��9�?�S�$=��=d�=F�I=�@=�.���T���7б<W>��7��:��r=��=ߟ?=�°<�6�O\=ء�;~���� ��u�<eLD��g=��<�g�z=�\F=.�=�=B�N=;�$�\�=#]=�js<��<V�Z=�u<��O�F�?��X�i�o<m�=�*Q��7<zO�:em�������C�e�:	���hЊ;b�h���<�T9:��3=�
����T=��-<�e:=@�0��0��\;=8�m<�/�<RE$:#��:�N=��{0P�rɧ<��\=4�����j�=eIC=(>�<��9� �˘a��xn=��S= X=
[@�����N������d�͔�����D�3=���<"K�ܹp=�u��c��b=f�<Q=B\�<�,ɼ~��;��+=�s�H5-���;4J,���`=RF�E�Z����<�[�؎��;���?=�W=���=C�<nm�ݙX�*�==���7�=�a�I��<M~J=K�9=1u�#�[=a�H=���;�»���A�=0=���kO$�:�+=ه��\����a���<�˼<K8)�.P�<[qY� ŗ�qI�J����F=���<<��p�;��:�9�]�e�1L������^c<�|[=[�;|�N�;$="�t��=p�,<lO=^D=rO뻌��)��<��T��E+=t�/=�z$=�Zc=�v����_B��ME�ٱ[=��'=I�v�U�9=\�B��=�4�<�Zy�?!=����g�EW��;<��;0&�<�[ =�b8���u=��
=��=7��<���<L���/�Լ��=͇��6i�Dl��syV�^��<i`�]�=-�=|8/=y�	<��<�^W=�4<u,�,�=!c�;�oμ/�;�޼��=�s��hfY�k��<�2#<K�����b=%k����;��><ǘ�;|i*<�C�<��(�L��;4�<*=Q=�6=ݹмE�T�5|����<9�<Ƈ=�N�<�K߼�ɼ�ý���=�Vx;��Y�h�}��<56B=O{�;;ʾ���0=��;��E<#�K<"�<��x���I�<�"U������I�<8Rw���)�3��ٖ� �e:QV9��%=x��}yE=��g-0=~��<��<��<�t��:ۼ5����<m`~�	��=~�*�a�:�\5=�8I=R�6=�qE<��J=�'º 4=�Ky=�a���c��}�w;Ս=|�м	�"����<�j�Xe=�3��JL�u�:�nm���=���<�
�;��q;���<QՕ��㻼҃F�Tw=\A=�7K="A����;���<-�+�O�&���<y����lm=+����l��ۑ<g��{j���T=��;5�d=V�A=�F��*�j�><~̳�0K�l}�<�~A�w��==�8�<�=� �<�a�<��J�Z=3t��H��-;�`��g� �%�T^���<�A�v�9c7=�7�LY&���_=­1�8�����X��<9���sM�C{I=RR�<�F��Μ���I=�jʼ�><{_=;%��*=\<��~=ץi<�;�FڼC�_=ћ�<D����=z\���ݸk�����R=�K}<��=1��<z���P;�@���S=����@���2�N�d=������1��>=A�d�f�u=�.ֺ2�=�࠻��O=����&S����l�X�8=ts"=����P8�F37=��H��䪼[�r=x�*=�;����h�2�\C��5(�<�~w<���?����W=��<���-�b�O��8��ĘA�`��;���<v�=�J���_=�oK�B�E<��&�uN���t=�R�<�a�<��ۼyDN�(�<�O��Z׼ŘM�	��<)O1=�VJ���üTl=��|�=��e;���<�-�<�B8��'=
K=�s,=3��<ͳ)={��<ଏ=&r��/L=�4=Gv<f�<L��T�<ə��&�=����<��<�n[=�=|3Լ _T=�?=ځ&=4P�b��9�\o���d<s�]����<(�^�<Z�=U�<=�[1���<�)��e=~��1�s=:=k�O=]T='֖=� =�;�S�3�r#�<����xK=6wH=���Q�`=D� <;�I���,�<���]e�����g뻶S<*��<#�_5=��=Ne<i��<oJ<y��<O��0�>�ky��Sn�"l�<�o�<Eq�G[[=��;)�z��fy����<e����G	=���a���Q,=�
a=�lI=2EO�?z���{<x[<�*��	�h=��=ͺüE)�<x+=^��=(8=�t����c���H�(�vٳ�c�`��)Ҽ�u�<ѿ/=��H�7d <&\�<w=�=���5b�Z,�<�s�;;Gϼ�I[�B�=-?;���5����Ҽ<BQ=&2Y�0���AD=��=9\=�P�<UJ@<D��<d�{;Ow�<Y���7l=w;V��:	���-��Z<��x���x�:e�:;e��<?-��E�<�<�l���������&!<%>=�W;�3s<����oc��F��ӝ;,��;�Dc�5͸<��w=wU]��l=�5�:/�Z�)�=&�˼��!=�E-<GJ_=��W������X=/_ϼ��7=� ];�=�����&�<��-=�!=�<hf"���=���<���;d�m��O=���<�=%�F=�Da=��=.4�<A�;<�(�������N0<0i�;�X�]�%�X;o��g�<�&=1ń=!������Š<��g��7���>��!������=���m=;='%@<�y(=�GH=uO=�)=��$=��=ЀS��-���麴�5=����Uy��E��_�:���ɼI�n�;�����2��U|=�ټ���<�P�;��L='��ܼ <��]=����7=o$ȼ�4ἂ~ټ����z�.2�_�]=�7��AG��S:�J��
n=C=��_��uӼ�R�;�$�<�A.�z����ټq����������rŻ���<nim�3Ki=��<�
�;��=�o�����)"��|3=z��W$S:
`�<�ǈ=EG<�=<{.=>�X��֊9��R�Zo��&TL��^3<��<��#�c�s=\��<�Ԛ��T=�}���+=�Qq<�M=���<����`+I��=ے?�N�X=��A=p�C==6�:$�I3� �6�S=��$�C�Y;e�5����H�d���:<2�w=2S%<@A=1
�@qG��N�;����9iA=gϨ�����F=z�4<^
F�1�<�[�=*�;x6�<��Z=���<H�{=d�����;#=��\�����<q�~�FF�r%2�Y��<Dp���\���b<(��QY<Ê����<U��<���?L���:�e=OE�<.P<�=�A;q&=:wW�[�<�c���O���;L��;᪂����=����}��<}�c�=\�>�s?;a��)����;���~���k7=&�;o�<7�X�9g޼O���M"���A<�vP=��;������<p�H=��I��5
=�V6=CY�<�U[=v�;<��b�\�C���^=(?=9?���[<b�����M6c=�2�:�䃽L��<�7=?�-<�E;J'�WbI����<:繼|�L<���p/$�qp�;Cb�XMK<�V�<��������7=c��:6�<��T�,=��s���(=����a�r��@=��x��ڼ�҈����<��&<oG-=�ָ���<}��@@�Ql�<�^�g����<[��Pt=a�<�Z�y!�<��<��%�����v�<��\�s8=��,<8A�<+ _�'����t�<���<ȉ��b��G��:�|��z,�ܶ�<�p����2�»B.����p��ѺJy�<��<=�d;�oQ=�V��,��C�= PJ<��';�Շ��?�<M�.�/b��<)I<�C|�e�໮l=�T�;�8�:s�i��A� �=a�G=��B=)�5=��L�)��<�ϊ<��?=ґ��
c����p<�}��)�B��4��eN���t���<6�9�N�l�!2V�RjF=oZ=�lT='Z0�ӗ3=�Հ9_)<��<�i
=h�x��D<=۽��X��<��X=W,<������u�V�=3�]=�h���4ļpO;��N==}.9�a/��UP�^Y
��
i�L|�<�R�w�=�+</��;οN��_U�;��<�a��+=?>�<r�
=�:����<=j=v;�����??=`��<���<�X�K�T=o/��,�Un��x�u<��=e�_�'=~�<�������;���RX\<M�<.��s�;�t$�!Bs<E�m��5��v�<��$=p��L?6���M=���q�����n�:�<=�!�<<�(=�	�����<�/=_�<T�_=.�=�4lD�92^:-�Q���(<���<�<�=�[�{�����;�"=�=�U�=+�'=�͑<����p�<��¹�ڕ<%�ѻE+�� �SM!����<;�<�.�<ʉN��>�:芼��s��Ĳ<�[
�hqQ�=�4=��<B�z��) <�Oo��N(=X2��9�=�
̻��<�����
���'�5��~�޼��_�q&=F����^Ƽh0E=�?}=��?=�c���_<��<.�=B��-2=-a�<-ͼ
 =��=xc�<��<���<�<%�^"�<Ǧ	����������<��Z�RE�<Z��#eZ�p���K	���z��;b��<�@Y�U�(<ՠ��miѻ-�P��H�tb����� �o�B��<m��<�L.�㿞;�X=��j�D�� `,=���<p�<�jT���7<Q=v=IM=�"�<�v/9�p#=�%����e=I�=V��3;=�Tc;��#���@<��;�cb�R��<�|��ٻ2:��@<�$�<���qx�<q�;��&�w$��.��X4��AX=X =i�X�;�m�<��A=��P<�C$=��ůC��D<���<��Żv<�~!C=��<� �
�y�٦F;SB<�;��+8(�� �<k� ;�c=d�;F�@����V��k&��L��b=�����<��`=��� �ho����=�!=��ļ�Co=`�$=�B�˃==Ⱦ;|�&�?=KB����M:��=-�
=򫼮6��Լi��<N\��Y΀����:�W �� ���+<�t��8q=(tv=���$ۼj[3=I�U<=��М=sX�<�4	�-���8�<�9�+�=�:����]l�6��<�-q=R��;��Q=���<��X=��/=nc^;E��<9�P<<�ܼe�A� CV<e\=�1Q=W+Q���鼇�+�q�)�_V�<���['=���:kխ���W=]�B��=�,��j8��=�<�}�G8�Z��.4�F�;}v9<Ɛ@=Q��<�'ʼ�N�<��5�ÔJ�h88���L<�L��<̀D���p��~�{�*:���z^���=2Y<I�3=�Jb=+<<� �=�uS����=�T��@�C�����*`�H<Hy�<<;Y=�=�Ga<^�<�"h��<;&�<W�<�M=�����o���'=t]��q2=�L=@�����]�p�;�<�^�<���[�ͼ�' ��� ��=w� �]�V�����������/d<�� ��:*=)tм����,m�< bջ�+<'�z=��f<�4�=392��p�<���ɑ=�����V=���A�<�6��%�����W�]��f��ƬT=k��~t�}պ�L�<��b���'{=�w=v-�aQ�7kݼ^Ci=ܨ?�"�j;�+�:�M�Юw<��=l�?�M���>?���>=��+��g�<5�H�}�X=�m�<���u:��=<�<��6� ҹb�[� �E���<��j=K�A�$��=�!=���<B|�<B��=�g�<�7��wd=�߅<$��<���<��*<� ����<$��<Ԃ=>=9�p����<��=]f\<L�����=u��]̔��
�<���<��9��μ�7=R\=�� <��\X=_TI�B���ۼg�/����<�X�D�J��<z��xȏ��%�<�<����[=�z=\8�=��<��#��D����=��+=:��=^��<~��<�=h�=�f;EK�;���<h#U��O�H�Y���?7L<�	��~+=3�~=�U����F;ߴF�>N"=�|�<.��hC��ゼ^�<uJ�����N����a�M����缇�Z= :9����a!��x<�<|��s��gSW=��M=�<%�[��/�<��:���K<��;����!���r�kT�ޔ$<<G<�������T?���D�E	3=��%=���<YZC=��b�TX=~*K<��=�Q8�������k��kN���廼~�=�t�s��<�T:��^=VW=� )���9=Z:�6���&3q<����"0d�s�=3_���O=�Tl��Q-�w$���<�.缌��<_>�<J=�5�3'�9��=R,�:�N7=��=���<	x�<F�$��R=kS=���@˺��<	��5H���j;�����0��l���q���O�=�N8���;��;��мgT��n�S���<:�U��P2���	���ϼjQ�w=�<$gԼ��*��[==P* ���<'��$廼UC �˹<9��8O#���T=>i*=~� �dx��4���#�=y�U:�W =�}-���6���
=��\=�`=�=Jy�;��p��*���'��wR�_ݺ%��ؓ<
򼈜=�At<��<3M�<� ;�4p?���X�� ���� 4��7�;��S1����<�T=����;���i(�<(�>=��,=��:�J��ot<a+�<95��1=�!=����wM=�Z<x�=��|=�U��&��)��F�r��O	�߇*=�q޼�V�<���ګ��0}�=�E���� ��C��<׷Z=�u$<�}z�4e�c͆;(�s=�XG=�j��9vb�PJ�:s��:���<��g�µP=kCj���@��<,;���Ek�<Xo߻߶�<����q1�<$���6	= mc<�
����(�|�<4�S��Ӿ�ʭs����Q;d�#=,��f#������[�;��<�q<�X�<W��<�^=H�N�Aռ3\�<h�J=��L<zϼx�#���
�]<�=mXr=^�ݼLN�;�u����<��û���<�x!<�Q��+fq�UW�~-=��Ȼ�AN���=�$-�`��;zP��|�cR�:�|U=��F=�0';6�,=�dq=hM�T�Q=;��<~�;�ih� p����M�E�<�z�<��<�*��ٴ'<��*=i�ͻ�y��Z=f|m�p�4;_�;��4���'=1 7�W/,<K̎����y�Ҟ�g����=Xʣ<��m��AD<�~^=���< �:�p�#�XX�<{"<Ė8���l��A��J<\��*��J"������$K����U�P=q�;Υ<ÑQ;"n_��,�<Z;s?=&A���1={��;I�Q<��D�6�|�.����*=�;�F�L�@��Yw$=�7�<ņ@="<˼��1��c���ZX�C�p)=�=�y:r�7e�<��:��<���:UH;������8;)g�<��O���N�?�x�'t<n����p� ��"�:q#��oE=��%��hg�xڳ��=M�W=��'=&�x��y�<����E�W:j.|�~��;`&<�Sѻ��=�:����Z�y�ۖ��,c=J�%<ių���<����	=E,�<�0=S�;3
�<�=�:���� ��w�<�jc�0��<��:=ݿ�<�w�����j��.m�;��ʼ}�M/�8�k�L�^�%��<�Hi=�՜;�.<�!=�u�<��:�N��x�=�ӻ�&����k=�#o<��_;�+���=ǅһ��^��q�����:"GǼ�=��L=�Z�P3(�'���M<�L�^���[����<ň��L7���<6��<P�����8=#+���T�MG=���w�g=*%&������;�Am<���<�ڒ���=��<�GK=��<����tμ� n=�wV=��c��B�<M�S=���<m�5�=[��<8l=�x���
<�N.��v��)��i;�<H�-��Bh< ���x�������UP�E�(=��<�8=Y1��&����<�e�u�q���=`�<\�h�g����<G�=�d;�59�<�T=�*�5iG��2��<~��f=��S�^=��%����<#��<+#�:2���R<r�=�I�<�=��A=�o�$W;ĆY=2~#����<\���Ƌ<��R�(u=��;'4J=7��;� ���%=�O,���9�-��:Ƽ��@�'G�
<��S�m'�v���	���=E�k=Iψ;�i=�)U=�u�<�*Y<�r��`��;�����/�ڐ��E����)>=m��<�s���޻<|����ĺ��#���,=���<`���1�<��>=ƤZ=3��9�|7��Q,=� =�?<�*{���l=�8�C� =j�G�*:��\�=�<=����ed'��5<ԩe;�cs�/�ۼyW7=^-=I�G=�cJ=��=��{=�E�=?�Y�l6�==&�<�����<3���E=Sр;+X��3�+�L<Lё<�Hk<�$(�?6Y�Yuk=��=�=P*=��7<�
$�F��2r<�G= �c=�qx=Qu=�gj�ʆ���l>�����޻�鿼�?r��I�l����3<�d�<cD6<�x���M�s������<�M=���<�Kw�u�C:���AF��Ã<#�Ҽ�("�E���<���<�p�<X�9�(� ��F��To_��V�<��C��Q����|=rh&=Pɼ��N�l�<a�'���V=2�*��/P�2P��k�<(�c;��F=m����;��&���==GB=-==�f�;Y�=` ��:w2�"�{��ɼ��"A��M��8��P�n��8<�ݔ<q!м�<}�=�e=Ѓ�<�D/=h����<�f#�_I�<:��;�4ǼHK<(+=qú�i�<�J?�-�==��8=vs<��R:���Z
�
<m��==����=��W�8P =��&=9zH<9F򼣜��l=DҔ<%,l�<X��<�Y=[�O=Ԉ߼��i�W�=��3;|��<c�7���e=aꥼ���JzF���������_�<2NB�9���8 Ѽ#"����==1\��%�;W_��;<=��+:6<cL�;����W����`��+�F�����0<;�ȻZ�F��k-�(�����/�{<�S\<�*"=��(��y};�==�5���"�<�&=�E<~	�E�<�-=�;=;�p����C=�<�j;�aѼh<��
=�<��<�E9�Z��<���u)���k=G�c�W�F;z� <ͪ=��F<���<��j��*�<���z􂼈��B9=�|�9%i=I=[�c�K��Z�5�-=>;�{}�<�ʄ:4r5=�=�H�FÖ��g��R:;X�	�_�\=h1]�l5<��.=��b=�$=�o=��ż�g�R�; Ӄ�C��^=o���U_��N�� A�B8��M\:�p�<�[W�� 2<L�g����<��=Ҫ8�l���6C=x6��z_<	X<�pἍ�?��=n=69�����9=�$*=;;=BT��n.=��7�ޠ[�GW�7$�=����b=:F�;�=$H���Z��<�;[<�Һ��u$�U�=W�M=`"=@ʇ�c��<�<�j�<�1=�+���; $<�K�:$ڻ��1="�<���<��j���������PA��=�=v�v=RG<*��<��:�	�ټknT=qż}�5�gqS��Qi�6g��L����k;tX=�f=�hb=����>���=��缿��<b>:�m=���<�4��Q��5q�V�ܼ)8(�G����~W=�18=h�Ƽ�ɻ��"=%<�ӱ��-=��8=�	z<��<�c��� =�!��^�<�5��9��<�=�y�mM�;j�5�Sp=��1=�j����=;�C�PҼ�m=���ֳ���"�P%=2W���q�<rb=V�E<���<n�W<.!=%3���ey��II�ÄҼ.̼Jɂ�mϷ���;=[�<���<ޕ��R��u����_�C=m�_=�d�n)�<[GZ=��"�Ay =��<҃���Y=��l=��<-�O�m��]#=��S=�e�������<R��vS=�V��*�L���<�5H<t;b����N�U=����7=��м
��<�]��r��ed�~q3=�B��~8�p[;��>=�?ܼ/��
Ԙ=~7�<@#�<���w�<�Op��*=�}�<"��<c�v��l;�x�Z;)�:�C�м$l<1�?=��m<w�=Gמ���}�PM�<V�t=I= <b���<HaA=ͫU=}�Ӻ�"�<�{=ʜҺ��<F=�=�cf�E2N=e�f<�.;=^º�`�g�*�;��
;\�/���=��=��<��<�<�F�F�4=}1W�SՖ����:kϻ��񼹙���\�<l���өA�d4��[=��g���<1�C���)�,�_=�P�;,���J=1��=��A<}�K9e@09��;=='�[9�y+<��9�b���<Z�<z.I=���x�|��.e�����w1<� A<�C�f�=��;hԖ����<L��<�?U�������<���JԻ�	��բз��ep =O����껴5�<N�Q=|�������s����O�-=.<�<�����>=L5�57�;��˼����6=����_�@O;R¼�Q�[�	=0�?=�iB�Q�x���=�)�<#kM<	v��:d���[=��c3+�pG���P���9=[��;b�l�y�*=��⼷S߼�����O��]!�Ijn=��`�Ǣ�<�|����'=�M=�yA<)��<�Kb;_:=�l2�d�<�@E�-��8���< 
���i����<K�h���༸_V<x+ἓs꼶��<���<��w��QB=ؓ|=[�к��;t?<%|=�!��������u��)�<
ӈ<GUC��%��*[;/�=�Zw=ϡ�<��<(J>�H�)���ۻ7�W�M�{���n�~�5�ֿ���<�;�:w��=o,3�:����+���A=!�
<3����<��I�<�f=�฼�>�v�<0@��:K��p���n�3 ���Q<[9ּN<�E����ZC�<��6<͜�<�[8��L�<LK��Bo�Ƚ}<�.!�9�=�Q<fD���+<\�=��<��7=�^9��S=O�O��n"=w�<]��=�ha=�&j�R��'���=$9Z���u��-;���<Da<�����-�A���/����<����.��=����ϩ`��#3�^[��5�<a�Igm<�K1;yz0�۰9�¤<��<W���D��:q=��l�Kf%=��l�C� =I���#<��d��@(�Cgh<D��<"T?=Sc=��E����<%��Դ9=���LA�<�z<mU<=Wm�8�*�<rD<�Ή��<�<��#���:�<\"�%DQ<���.�:��m=+l��)k�<��=�ł<�o)<���<ϪG<Y�%�*y9=��M�͈)=��������|=6�N�D5==��|�"��C�<u?������M�"��Β�>o=y8'=�߅��N��( �͓L�7�<4�4��%�;"�=7Q0��u��d;ټpdc��J���f˼r^'�BJg<�1��?+�l�@��)��B���<s��<�.=ʔ
�į���< TX<�'�<��-=�e�<��l���E�������E=?�<mWa=7<h���Y���<��%���=�?=��<��<qV=fB��<�U�`��=��N=>��<vJ���Q��ȥ<yn<�)���0��������-W����V��)Ce=P�[�Л2=�<�_=�8��w=b�g�=א�f��m�,�O�Q=휻^倽fߓ��	=��s��x����Y��E�Qd�Gwz���<#�]�|c]='�$<�bͼY��<�]<zWJ=iO<,/D�X��<�� =�%���!��F=�<�9��̼�����[=~�"���Y��ߚ<�˼�Y��4���rT��r!=�=�R���<&�<�΋<��<2�</����~=IV��e�Z0�;P����L?=^�I=8K=.^<�q�W=��<��;Hc<�Q�;�)=o֪<�P</�D�BQA=�`�|/�'��<
�_�MQ�<�������i-����/b0=*e
<Y�����<JM�e�<P�=�� ;
M���m���J�Y������<|�Z=E�T<��q<�+�k�ʼ�R�<(�=B=Q*=c<ͽE���6=�O���8=���<ռ��rO=����w=Ov�'��u�%�\���A=�ո<~U.;�Ԉ=��{<`2���~�o�6�<�S=��;ei�;E�U��<d��<�fƼ�lw�N��O0K��\��oV�2B�<r7<�����<�S��]����E��Z���F��Sػx����'<��='�/=Z���S2�߁$��ES=��1<����� �uA�E�<�qv=4v*=�H=�ټ�W�<�ʛ<P��]���P��3����<^�g<�X%��o=Y�Ѽ~$-=D�$=uv?<�ȧ;�"Q�?͐�`"��ݼ�Sb<�E��n�;�B�5'<��=��H=ˑ0<���<�Ih=cw=��sQ�37�:�sD��
�TTҼ�1=ۖ8=!�_��_�� <���9rl�����<zZ��J"� pc��HR���0�d<Q�]�]�E�V�R=�#+��Ԃ���< �r=�0<=��=�<-��_=�I����e�Y;�<�<��g=�5���S=������5��;���<�Y'��#�<��I=��ZI <���Lh-=��(����<��l<ƹ�<s����D�<K�C<�
����<�p=�=���ZA<�:����[<�AQ�������=��g��-�<p�|;6E=�bغ@�$��z2=�-X=�	y=��=�>�l�@�����1<��<ė�<h��<��/=�	v<�)<�=�<��V��e���P=�e�<m�M����H�k��<*d=�xB���<
�1=݊��S�ԼLL�}�8=�e��Ϛ�	�;�:�DoN�CL���:���,=@�=��-�ɿ��0@�Z�m���1<�P�<h��<*����3�-��<������܁���r�����Ļ&�A�/�����k�;�y+�,��@����g �B�b=���T�79p/�3>=�
o�o6=ַ
�W���=�;zeM=�ǻz1O=��T=��g=��<�T�CZ�<1��_�<��4<>��K�λ_��;�)���L���;�Z!=tc��[=.H�=���%q��;�<��`<V8v�Һ1;�)��Z���?\��s>=5K�;�~C;N��<��</x)��s;�%Z==r_=��:=+k�!�����[:̼w�h,�e":AT9=q;�W��<cE�����ךZ=j�}'��o{�<�==` H�ǁ��9|�4����S?=۟=�|@!��_=z�<�V=(�n��˺co�;�
=�Y��ݼ<F�i=D4�<7w�<��S;Y���6�eB�<�<K7�`�:<舠<@�?)�:-���=n�<�M�'?�ч���n#���(��ࣻw�]:��H=��<��6=l{�;j��m\B<�Y�<r�w���=�}�<m�Ӽ������h���i�e=T��<�ӻ'�1=��;Hi�<}ѭ�W�ܼ�z�<�H��x��FD"�g��<3����jA=B�l=gMȻ���<�$��e��^m��J�,�@���X\�� ����;�Ǡ;n��<pe��'���ֻh%h������s
�I�ɼD�����XK�Ċ���?��X��X�p=�����k�'):Xu�=�=�<9�(���`��=�ș�Ѥ<��C=�%=p�=�&��軹�P���: ��p=۰k<��}<�u�t�a<��\=cD��KD����;�Q=��o=�O�cA�<x�<�7�<h�T<7����Pۼ@�!=ت��\=
�B=U�=Mл���3M<�RR�/5�]�X�-��:!C;=����;b���=����8W<���<GC��w嫼��I�<�==<n�2P'=;�=A�I�t�;�+7<�v�<�3�����V�<��U=�,=D�<���8��c�&;B<����$���Ty=wp�<#u	�ۖ�<O�L�Ѽtd(�C�H<��'�O��IH=�,,��i�"���n��G�<C�w=n ?���<^�	=a@X����~�<�A�\%���f����"=vC=��<�ĺ�=		z<l��<�r�<��A���;�g���h��D=&=e=]C�x�]=�?N=���<"�;n���������4��;�F��������<�=�G <��?< �q&=I=�eI�P�4;�I=k�&=27��Lt��W*,��=��<�� �����c=��F��8T=Z�`�mU��w�X���B=u�`��Q@=
�Y<�5�⚌�
8�6ae=X�	<mf=��H=8j�;��E����������;W	(<��^�����=&�<bR�����kK"=�*<�=G=X�?�����\���+��kD�0wػ�Wۼi-=�Ԡ;����ŋ��+�6f��j�#�j1�b!�Y�>=|@غ�[#�h�ļ�.�<\.=�������; �U=	� �u�M=а�<�V�<��<�$2<�*���;K��=q��ިT=Ԥ7=�
��x��� R<��>x�nxռ�������U�:����<=_6��@��X�T==�*<g;ӻc� =
��<��wA=��<��.=����Y����=Y�<��<��ݻ��A=h:��,='+W<��k=�+=Ia =��@=8�ڻ�mf=��+���D&=Z�;����<+��<;Y�<�x=S���8B�lZ����;�,�:��ɼ��<�Lk<8�<=��_��P~�tC�G��<U�z��:8����
�	<y�y:�zɼ�;�j�z��<�T;6h��fvz�����0�<��ݻ����K���<�A;I<ọot��R?<.B�ڕ&�*u=��<��;pU���#=��<�w��z���n+=�3�<������<�>���ռ�a�<W�@��7�%���zn�@���%����Z��E^<�H�<E�Y=B7�y�T=��y�;�&<��3=�N-<Z۹��众e��F�<_�����;j��<(i4�"�u=�P�BP<D�J����+a�<����"f�-'k��@�0�;ڏ�<L�=}<��([�ȼ�<��\�.�ߢS�i�K=�"g<��<FI<��N��;��;���:�=X�r{U=T����,�<�@���e9=`N�:S��=��c=��aA9=�A<���;T="�5��}Ȼ�Cb=�a=�<X?=��5�4���=2�!=���<��<��^=���<�Ҽ�T��H�XaG=�P7�'=H�<�k�<����5=�� =�?=���<Sdr�w�R�S(;��ڼ�=oa<<�<%�<OZ���*�/�<wn#����;d������;b���f='r�{�����$��bv= B=*=Do������K<���kp�V�	=�N�y�
=M</=��;��< >=�'�<-�ɻ�g�S@�<��U<�D���Ӓ;Q���(7���<v�BK=�k�<T3���]=b���;Og=,� =]��<#ٙ<��==��W<K`h�a%<�Tμ�#�
A.=�K�z<�ڻ��<���;�5=`i������D:=|��X=O_=�&�����<�l�����jh=��@�3=y�2���_=A�;��=T��Bǘ<sQ��6�����<�C�<����z	�?�P�� =�����+=�<��=NB
�˔~��X<��ܼ�X=�Jd=�I�^�!=�]N��_E=+B�<2{�7�)=Q+�9l��;B!W<�f�<�CY<G�2=���ǡ�<^�=���-�<��U������ �s�)<�5�[�t=.1�a,#=-#-=�m��p�<s7�<�jۼƪ5�(��<��/�r|�<�k<4?�<�TO��A��$=%��<mY���v/��e�<�I�<��<�X�;��=��Y<'���&�Uj�<��ú$U1�b� ;*���-�<��p<0��<
%=��F��8=�f>��u�����=��Ǽp =��J�)��(�<@��X�9�L@��vE=��%r\�����3^���h=�33���N���<_p?=��+=�����0L=���<�X���&�1��<�r2<��k ��"�<5+�� �<-�V< �< GI<�}���U=ŋU=$�<��UW��EҼ�Af=̂,=�;=�wں[����=��:�k�8S�<u�=![�;̧/=_�;���#�O=�+<5�M�*��<�ѳ�j�f;ۍ�<��90����ۼʯd=��Y=W�s=��<�i<���;z�^=T��<�٘= �<�~ ����������Y<��'<SL!�u�});�a�<٤b=��0,�h<���B��5ݯ<~�<���������^�Ҟz� �$<�F���>��򼡛m<B4�<�-��<%=��&�*W=�<N~=��:���n�R&==w���;�\<+4=p$=	l=�h��Ɔ(��͚���<�2ռO���92<c7�����<�Ц��@Ƽ�(9%12��p��5�>�H8*=RNa=����o<���NO'�J�'�o=��8��R���t ='
�<v��q����J��+�ڼ�c���E;*�8���]=�Q==r�;-Q��<<#�鼢)�<j0�;�E�	2=sK�:^��~��v�=�Ň;:W̼m=�饽s��<105�����HU���s���<�:��+:WY=��M��a�~�<��>=���P�<NeD=�R��=m��*�ü2�k=��_�$��<�1=���<�f��b3�����"x����U<:a����{<K�=lK<[��<P�_=�QW��b =*�5�4
\��3=�5�;RU��_�:�E�<nYO=���<rb=��m=L!'�=f=�}�<� ļ���=��ɼMq�nX̼���<����L=���<ƮU��E7����!�,���Y=�e��Տ�=��<�Hz�a�f���<>�߻Vet=x�4�����7Y<t�=�3����<̓�<�4=E���D~�����Ȳ��{1=ّ޼��"=�*s��f��w�<�a=�>˼��K��t�-�.=�
�W6=/���θr�\A�<g
%��X*�=�=��n
ټb�;&�z<����-�:�Q��%��;�'� �B=�&=/>)=&L&<�{ټ��5=\	=��=�����=�Ԣ�}���	/=��[�HMQ=�?<��#�l=s��=M=G�O=�S��b#��8=Shn<.����;���k�p��<�r�<B��<7����"�<�t�<�:��$;�D=ri��ҹ�<��k��P��%{�0�<����#f��P=InK;��<r]B=��0�9��
=�JP��z8����;}xM=�lȼ8��9Q�l<~=�Q��:����~��<�p�o �=�<<�F=_�<7����ev�e�/��	=��l<��K9t�:;��<��H��6��_�1~)�)6?�ߙ.�����C`�u=��!��i�����(B��!�;�<��=k�Ƽ�n�3	&=5.A���:<���<$�5=!�Ǽ_��<&k8=[i?=�Z��%���ἴ�@=C��a����<e���=W���=H=gcH�Iᴼ�D��=l����5�2�?�����w��;�\�����;ԭ������%�< ��<WGS=��3=��J�\�<���<@D�@`e��@���g��Fļ�;��>�G�b��<}< =ְx�}�=�P=%+��m	�:�<;o���N��=���D'U=��,��#�<�!B�&^=A퀺�r=c�:Ş�;��T�q	�<[��<]Ӻ�fW�aѓ�O����/6���K��_g�Y <=P��*�z=�2Z<ٛ&=��K<݀�&��<�)�޴<jټr��<^��=-Yl<�_]�*�5=�bP=n놼n�F����<�,��G�<x<&��/=r�4��#���ɼ�]f��P�:�~���]=�:��_�=�҂<9�y;h�ؠؼҵ�<�w[���P{��I��<�%�F0�<���Q�(����<����!����)���%=�w#=mF?���ҼDOڼ&�-�=
*=�P�<�9�<|�"=��0�!�c��D<={��>*,=4A�i�=��I�Au���ȿ����tn����'=<�c��&�<B�b����<�L:��]=�^���D�P=��=~��Һ��A�*�M�xM�<�w�F��<߅=��=W����`��=.����Y�H��<��f�a�����H-�=/&һ����\��<r���T��:+<�{^��b�<W�<\�<
]d�.;�W>;��W=pg|=ޛ?�_�#={�A=��<�}&=��K="X[��c�<.�=��==I<�C�:O�X��̝�xr=�z���<��޼��"��H����aOҼ]�_=�]3��=���XǼ�q;���!^ݼ��T�AA���d=��%
W�q�F�r1(�9B��DT�$v�<��-=�1�<��4<�M߼��R=/�]�.= �c=ȣ����&�2@��3/�+z4��`���0�ūf�)Ѿ<�T�������qi:Ex"=�{=yq<eƗ<oQ�����c=��<9�k�(kͻk�Ҽ��=r_�<n�?<-���3�w<P��i���=�8��� ��,F<�q�;��=Òr���K<��;[�����;�9?�`ϩ;+B\���C���<I<��+�ws�tn6=�Γ��1.����<�z=���<ߓQ=.C�<�]�<���=���;�4�<�¼�5V��';�P��I5�<���<8'?<��<T�a�4t���>��n+
=
�=��=�)�=�ॼ�[o��7�<����x�Ǽ�k;G(8�E���Vk<u��<w�=�m=���<i�V=�뇼
��(r=��N=����,���:��6<��G=j�T<
�A=B��<+ڼ$�,��Q�<�_b���Qg��^=W�j:��<*��}i�'�^��඼�c��y�_y=�G�/P���q�¢<. ����<i�<\�<�P �׊i��g�	2���S�S�@�b<s@�=���;��d�2�O�+��A�<�%�!98�*=t� �~qJ=U�T��`�������*�����1;�W"��֧;p,��=��Z��j�<��<&D=i�<�SRT=^t�Qۻ��;&�n=�C�;��#���漵C�ls��ꆟ;���<�R9�`��<bd;���<��=В�<�ܻ��=}�=M�6=�B=<��<�%�<�Z����<g�3�Y<��z�(��$�c�C;W5=�4���<�V�<K_=b�8=��[<�EH���n���O�tF�o��Hn0<���s��g(=��<�?�<�c\=��;y�=����?<���<�L[���<c�g��HI���G=�6\=�_���j=�b ���;���<U��<�/��V��k��O<����������!�=��<B�Ļ�e���t׼� �F==���;4<I�4-�����|���Ez�>Z/�'��<9��<
�T=��L�����;,Q�<G.F���7���B���R<��h=��F=�쪼��rl��w0O=<$��5D�i;���Һ�1�!6���_=��=V&���6��c=�)=�1��=.����=oD<�~e��F=�1�<`y;=Y�=�fל<e�N�8��������	��=Ws@�k�#=��m=�/�<��	="g=����O<w?=�%�j�4���	=n���E�ȼ��ڼ��0<�-m�@��g�:#�p=Ť�Eh����1�k!�<���;<D=7x�<�5��Mz�$�U�;���_�5���|�DL���Ӏ=*��;a�#��97=�^=p�e�2M=&�=,j�"�.<]으%;�;�k.=�!����p�&=]K��1��ޘ���b�w>&=�ؼ/ؼ*Ť�:ZL=,=����;�}�&H?=�J=�ę��{e��b~���[=}{�~�񻟗i�v$=S�w<�g)����E��:�\X����<k���ʟ<3�_=3W�4r��r��=Oȼ��`<�K&�̽	��0=_M=��;���#����]BJ9���<�j�C�;�}c�����r(�0i��AW?����u1�P;]�=��<�(��X!��1�عA��=Rm=�_Q;��G�{���i�<��b=�=R�i=@S=d�=hȮ��i�<!�$;&ċ��� �Ua>�.��<A׺����id��=��<f��Y!"=�{�h¼��;�d��[u������P�a=�k<�:���<V���R�_���N�\�J i<��=[=ݼ1J1=5����W�<����F�ҼF;h=fV=�=�_������Z�ܺ�s<��ü�R븠Ž<��<p�;��
�������ټ��м�: =`����A�gҎ�NG����8={e��A��´<���Ă#=/=�<ގ�`;B=`r����7=A$`=�V�;���d��<s��<��<T�<[Ԇ=B�=.�g2k��Fo<��<��;��#=��;=�n�&�
=|1�;K�=�3<����-�=w;=��R�?=��m�?���_<į�ϗӼO��k=&]z=�+����,;�f����T���a�0�P�i�=[P\��@=8�K<��[=�ˀ=��=6W;76}=4w��C�M���<�PD=��	����<s���^_��i�<oU�<̼�Ό�m/;��/<u[=��7�c����x��!��+���g�:=��<p-���h=��+=tj���L=&]�=pE��?'�'C���3�n�żlr$��W[�(;;=%߻� �Ҭ �a�I<3��;��
<O�˼��j=J�o<kz�9$���X�<1
g�"������<#�;gD��\����=�i�;��<��ü�5��mfO��㠼����*l<�v�<�4=&rx<w���1V<�+:^�T=�s5���=s���i�<<�9�[.M���<Ub�������<8{Y=�7�<^��<��='��8$��<s�k�-=9c>=���<))�����`F_<�A��JI��Ԅ=S�O�h�
:H�K��<�;5��]�<[��<��^:Z=�����`�ů�_�4=SM&=�;=�����%�Tނ����fF=�˯<��=��<ml���[8S<6B�<Ѫ<�^�<Ϲ��k���i*����g$t��;ML����<��=��9�	d���-�q
T=�����k�&~b��.���n=�H�<��=C���B����<��:��<MQ��D�:q��;p�R�I�{�X��<�E=�e�l���O�<{:� �n=W��]3���[��D��Hw<����s��=p��:��%���}���7=��=m�?�� 6�2)ļ�+��!?=Z�M���G=�U��K���Z	=�+=v���h���<��<��=N����OƼO�����!��ļS�8����B��<u�q=�[�;^���!��Nc<����/Y�4R��>=�{�<�=&��<[�� aE��P&=G������O;��%�;�E�sr�<*�=E:�<x��<�¼��1�i�;\�����~����;c4=F.'<G������k�<p�=]���������5��{�����p�=��;&��<�.=��;=�G�<��o�l=Y��;�k==�D=s3�d�d��<��?=ƼL��@*=�IM����L�Z�Rl���e�I����k5�r7л�򍼃�=��;�P�$=@�=U����6=�=Fq���=URk���t�V<q���-S={|�=Yܤ<�f=�.$�9U���JV=Po�<���;Q,R=B�S�?�����4B=o�<o	=q�=��^<�켇z�<3h�<ǘ	��`u=�<ݫ�<�u=c��5�%=!�,=���AX��yּ?^<L�[�RK�<�*ֻ����$��i%�SK�<T_�bQ��"{�M�f<�9���U��pf<�����Dd<��=�^�P�=&�^=|�5�"$�+���_^=�G=�|6�1Wݼ�	W�|ꭻ4��;��-�$6�;��<b+P���=���;����(s��0;����)�<f�V��o=�?�;�T�����좻<�Dm<2�<�O��%$==u�����	/=�&�H=�B
�O�&=EA�;�y༓��<J��<��;*�E=h��.�9=y��;����{<�$�:&=��j��>=*��{ș<"���"�<n#��zc��QP<aI=ᳮ<�畻(/==>=!X)=:�<x�-����S}�;�4��ƪ<»�6T����;��=��X<5(ݺj�~<ǿ��e;=��>��EN=i�8�==]�%�3�!<Xֆ� ѡ<[�K���D�2-V��By��<��Q�����Ѯ�2zJ�2�!=Md�}"��r�9�ܼ��<��o�r�u=N����k;��=~�c�*m����<[��?�;��<e!=vR=��-�(��\��t�<䌍<-�r��F�<��뼼TU�O�
��*��<�"0<8�:�!�<�2=ۥJ��TI=�fT<�r'���=�D'�^�<����2�5=�-=��=�~(����<~�\9�>&=B�v=_�����X<v�>�|�>=2A=���<�J#<Z�K��:-��5��u�?������z�[i��v��<1$S��PF=#+;���;��
�1E<�fS=m�e=�i=�\�<
eL=[6�tb<�Ց�m˓�;cɼ|$��c��˴2�G�7��H<;Q�;~���gK��x˼��<��O�"&R<��/=�gU=n|�	�1<��λ+�6��BT=z��?=�t#�``�<ѶA=�v�<b弪y%����PNo���'��5�;�m�<����&<'	�<�7��$Z��g�*�u=��Ȼ=B�<V�%<w�m=Vs!�C�4�eeu�!&t<1�#w ;�i$=�!:Q�?��
(��!1=�=U���%��
���<I�H=-X{�K�f=�=5<�಼:�$��o��Լw^�;O:t=�_H=,:��NEG=� C�J� �ڸ����;J��K�[���!���[u^������F8<����<+�<}z���y<{[I�
��<��M���C���=P��D�������,����M���Y=�6=�a�<p�<Nt=�@-;�	;���򁤼��&<�<w�h;��*�M��렼��鼴Ee�h��;I#=�v��ǫ:z�)�ɋo��pQ�Z�<�x���L��';�^��>���+/������K�mʝ;YL=P1o=/t=�ߡ��`p����;Mq<��;��<��=惊�D@S=��=8,=!t'=b����3=�F5�_�ټ1t�;��(��0�<|� ��O�;,�=�?�<6�D�lμBhD<�+�<�_�<{H>���<eHs���<�_뼖� =��V�ot�^)=�%)���<�i9=c+f�E]D���L^�C<<�g=r:��d;bg��5�;�E�;B��;-X��#`���
=�F��� =�3�<�z�<ݻ༽���w�;A-4�!���6=R���ȥ*<�P|<5ν�c�f���6μ��	�u82���K�PJ�m�Ѽ�Z�<��e;��I��g���<+�|��Ѧ:ud]��L��n�.�1�=r���r�<���%ݑ�Ȃx=H*9=�<μ1�M�Osf=_p¼� #��,=F�2=��=e�"=��m<�*=ZV\<*�I<��g=��X��:*=������H68��G<f"���|W���[=6��o�<�#=&��8(`�Oռ��P�9��<�a��)���N���5&�#��;��d<=��f��A��ﭼ�>'����88�Q=�����R���U��x�<�nV=#�\�d�=��;%��� <�48��$Y=���:9��^�Z==!=ZyI=�JA��0�}�d�<q􁽚MM=�T%<=7:�f<IS��Hg���8=�t����"=|:ļ	����<��|�U2�<���B�=��{<FO�=1�<��=?��<ˡJ���=��=f�<X�U�]R�B8�)b<��X=��=��&��H*< !/���<A���Oݳ<���;�NL���2��J=`���ϼ<͛�;��\����<#&˼bG�;��+=�_�<���}���@4�S������RJ �e������Tg��*�<J�ܼ7/@����<F<񫒼�@=�s#�s��6�+��Д;�1�<�'�=��N��`=�:C�=qH=����K=@�0�3i���F<ٳ<x�<�	>=?�9�ZB����<X8��'= y���#=��e�:_I�<� �<�w?=KiU�=�
��p�<~�R�}d=.�;�n;����<(�\��j��0��)̼������j��V=Z&�<Ȅ��0��'�����!�u.=��<ܤ<c<=\�o_�<���<<Q :<�~�]!�+;,�%ڐ�`�P<<~=Y�:y��<��|<M�V�.��	�;���<>�u�Ra�<�$������޿s<��<�c3<���G�O=  �ox; ��<��)=�{I=ɮĺzf�<!�\��$=Nj'�LO�}�< ܀��#C��o=�d�)���@����a}�<_��;�����˃�}�5�NS�$�q��c<����:u��̍�8=��¼�H7=��A<[����[=*1;�u����	=-x���^=��k=��a=�9��1	��C<������=���{��<�s�;�@=!��?�s=f��;v-o;�����i�\ȡ=�K[<�I���=�<�)=�vC=�#����<.C׼��E<:���Ѽ�R#�-.u=JR�;*<��f��Tr�=��@=��Y�㸼�O��X�#=
��^��*(�V�P;����1;�G�(�� =����UK�h��<(
�g]�<��=;���6�#��EM���r�a��4��i�B;d*=!�;+}����&���;���=d�{<�$=f{����׼`r�<��e=�78��t]=�U=��ռV.I=7� ��qҼ�F��˫=к�<bT����0���W<p�u�^US<� ���M����]q={�=��'�H�=����Z-�m����=��@=����%�R�$�ʼb���sL��;(;���Y�<$ ="i�<�¼�����D��C�a*���<� :��S9�:u��<=Y��[0�Z�ԼT�5=��<���<�,?=�#=Yo=�F�q�<���w_-<�aB��*�<T&H=��U=��W=��<����߶<�h�;��j=� �<������=�vFC=�$<��i�%��=��T=���<Ѯz�Poh=	�X��+�!OE�*�f�X5���+O�c��<QLT���K���
���ӥk=(qY�z�+=Sk��ܞ<H����<����O�8=�7 =X�������	�<��-��v��I��������h=��=�;=��8��<=�?|<ŋ���*��+��rI=z���ho�k<T=���h����G�1���e<��<���xq�ڵ�<h�F�0|4<\"a��n���8=y���L��(�yқ<|f;�`M�/�b�+I�<�~	�V��w�>;맃�Lc<�;_���n=�"4�X���M=Yj<"�P:8�ѝV��DG<	�2=��!=i���� ��H5��x��,�[���C;���`Q��b�<*�"=~H�<+a⼞/0�!e�^�><�\ ���=��F;^�*���-��c�<;<�G/=��Dȯ�n�=F$&=z�����~V�����$=t*4=�^¼"�;G)����=D.=T=���<k-=n1=��=訠<�tW�j� �j���P.�����<q�޼��=��<��;=w�;<�{=oj
=�N�<�鯼��i���<:&���w�j�(�S��<Ss�;�C=����C��S0o=�	=�[(�]=AC+�I��pDs=����<��&��e�<*jI<���;>����j��U���-�<���<�r/���0���غiס���Ҽ��%=s��<$v=9�7=[��<[��<g�$�1=�/*�����D�������[�����<�k_=ׯ5�;��qn=����D=�N���7�bČ�7�g<!���(�~=W`�<Ap�<��<2=1=��K�U㳼�J�D=��f����{n=Qv��T=��;��P=V�7����k+�����Q�<P{���m=����\��<�8U���c=���<�}����;��/�Gj3�=�*����{w.���%�]�����Ñ�=P�8=�T=�I�<G��<dwd=z�P=y�;y�=�=U=�^�:J�2�p����t���I��m�P<9�^������M�����<USV=3Y<-�i���?=?V=kȒ=��;� �{Yy�80�<��<wB���r]>=���3�L=��8��}<O�2p�=7�<�@�7ꕼ婼|(�<��*=����vP�J�<�:��5�%�S�O#�^n<�h::&����<h~���.�c�s��!}��_�:������٠��g�:�f/(���t;^t�;�t$=�k�9�IҺY�=g2b��!ѻ$��iΈ:Μ%=+�,<�ʼ~_��Y+ݼS�*<���<��=׿:��yE��o� � �0g}�L���q���V��>��i�</�=��"=q�����<������<��q=�ff�$�=ա<�n6��T0�|�ü[�*���,���3=�?_����<���^�m�e=O�<=T=`�r�>��ؔ<=m׽;x��<
-=ފ��@J�J?<o�
�����0=1�<'g=(\���Ƽ*�����;����D�<:�t<�Cμ;Y"�@Ռ����hh��7:�,#*�M�Y<G���1_<��~;��߼e�=P��<u�Tg=�<��_'��2;�<G��<�ǻ'ʼ�<.��m5=77@=�=�<g=��ռ�Ϙ<X� =|Uȼ��y�<ɐ-��̎�*޼"AN=���<E�V;�!�<�.=_(H�!b=.�=f<���,��}^���7�K�<��0Z���<]�z��(��LD�������;�;��=�F=P���#�<�����;�%|<d�����`�<��<�O=p����+=��x=���<��<� �=���;;����A����<�au��s�<��M��=;���I���-��kR���'=�==��={���ܼ�z�b��NI�*6G<@;=�G;2��<K��<��<��#�W�=}65��c�<M�j=#Q�����u�޻�<��V=/���eO�<kC*�߻�<���u�g=��t=��S�e\=��<i�<�<b��=����<
�?=�J�<-s���u��5�;𺺼FmC=�g��N.=i���/�K�G��䉝<�@��<��g�_����n��#�ޚ=���<"F<��V=R=z��m[A����<#!3=�3M<�ꁼߋ��I��^:��x;�	�<I��;�@M��z��(��;�l���"�<+�=���<t72����<���<�ʶ<_�_�+	���u=�_�ݿ��3ļvo��	]������X����<�:����$ي���R=��;}�U=�0�<��q�5Ҽxj^<yn0=p�m�0��ItM=�נ<�T7=10�
Q=�9==Ɉ�;�W��Z����i�Z�S����Z��C���z�<pkb=d�%��H�=�Ɇ<�� ��j������9=�@T=%�=sR
�l�9=��9=#}�<�6��1�iPG<�}c=ª�br��pc����;#�_=�pJ=T�}=�����ռ-2N��ܺ< 9μG+�߄I�ڹI<q��i�<�q�<��=������"����(<61t=W��9ŌQ;dy�;	�����<�@&��׻"�<׳׼�X=�9��	p<1�S=��7=A�O=�醼�r˻?���ǎ(����<� �;1�=��<}~\<�J���=N=sg4<�V�9Q�P��<����	�;�s��=�;GV��"=���7��<�r{<���<��<���<m�O=<�?�	�S�G􈻌�l�^����'=��ü1CX=	Ѽ���Fxd�Ʌ��:x���	��G=���<tY�<�x"�.������.��<�R=i���]�=X7==�^Լ��e=�N�;��w<�Z{<"�W�'�N=N��=�&����:�y��x��n�<@H� 3,=����i;ͼ@a<n�>;H�7�;�F�;��=�Q"=��K=�C����F=g2�<l��3 /��<y���3̼f�����<�F=$Ǩ�i�7<���=�n㼃+��=����,�F�D�2W"=b��ܒs�Y�<=6�T�:,@�����P��:R�K�u=¢��$r�;O갼���<�0�~<�<|}=�z�<��!}�<�6��:_=t\]=��<�c�Hk�<�X���>����q�,��p=�5����.�=R #����T[<.�6�	�V=?O^=� ���]<�^����=t�H=U"=�Jռ��Ҽ��<��5���3=�(�<�W�;nř�ե4=Ż<�"��,L�<��Q=�QL;�_�C����y=a�����Á����,=F�V�:��=S =�0^�6v�	^=ςK=�D=+�Լ~T����E�$�=��;(�@���m�%3�;&��_��Ȕ<</8�^P	��!�<a�==�_B=/Ѹ��ŭ���:�}�=�Q�<�=�!��g���,;94���=�"�nԻ�a�<(�+=H��<T��{�	=��~<��c��;hE=rG^=/�JH]:�>��Źd=��G<�Y���m���p��E���]f=]��<���<�s]��=��ͼ��N���q��B>��*<�JS����,%=���<�,���~<�R����_�$;��_=+N���,�<��Y=���<�����K�8i���=׳���~�t��TR�g�4��2<��;z��<��]=yo������&�<A�����< W)�eF�<s-=W-�<X����B:�H-=���<�5=�~�;��=�v�;�0��;���Yp��������_V��:��g(x�>L�<a?�<�T��XK�t�=E����v��R4=o�!=��sF���#�+��=VU�<1(=*"S=�H�=o�)���=����<��=�#<�5�<�6����'=��%�?�h�F$�E/��!�f'= �O<&��<F=�;[5#�[��R��<eƼ ����X��Su<��ʼ����Ƽ�[-�}��<Gx=��!����D�l�^񽻖��<fv<\�:pA��
=���<���<�����;S=+�+�ߥ���QM=��=f�8��jl��3���ڛ��x�<��)�F�GY�<-K��M�I����8Ļ�я���9�*w���A=��	�(��]�#��������J=%���Fs$��b���D=��h�<U��[q�<��Ｆ'=_��<��[=�E?=տ��м�`r����
+�<�\I=.'=�!�;�e���Z�ys�g؁���.<-·<UU��I�1#�<�=Q��;
�O���3;� =ч��7z��� =�U�<��*=���*=w�N<
�x�K�=>�;�?�T�7=qp��Ocx<Et��we-��.=r�=��i����l=DE�<l.K=ؓN���!��F=�(��ļ�/͇�1m<db��Otݼ�o=\K=7��<]�3=$��<��N=ը��|��
a=Z�c��K=�;�<yd˻)}==��>�u>3���U�<@�x=�8�@���=��k=����.=.f��ソ��<ȗ�<f�������A���_R�P�Z=kE=�쑼h.�x��<hi-�ib<)����TZ�;\
���P<��;w1m<��<)��<�aO=H�s�ў�Sg=��/��B�8Ru=�`��d�����.*=��=�@>�2�S<�&�9�����<0E;=g����<����NM��P(��HY���8�	��;X�S�f/���ä<�*�v�E�Z��<��<nV4��7��=��)=)�̼S.��\�<I4����<��B=Z�;=QZ��ӵ�;�7	<8�!�0���m*=�?=|�V<0������º;�c=�2V����<}W��ۼlx~�.�Լ�����z���@�9N�<��6��!��\"���<���;��P�5Ԅ<
O�L�`�S2���~��֞�<8���u< b|<#��9�5����<^�<�=��.�!��;�#.�<Z�/�A<�a,��-�<��<���/�l�!W��s3=��7=�|��v🻭�<����Q���[�>�<�Q�<�d�����)^�<��<�4@;`�=�2��D<x�=��<��'r˹�O|�K g��c�в��j=��S��<L�l�x�'�4'���=ǘ#=��@=�P�=�<��V�-$�ҹQ��#�~Mf�~��<>�e���=�,�<�]<��=|�J<��B=w=�<��v��-5=�Uj<V�N��3��<r�i~ּ�������~p-<�;6�*=�Vo�F���s�~f;P�N��2�ʼ�P"<h�^�M�����=˺2��L��.o=/A<vp�NPK=o.�e���<��=9��S|~=�u\��׼~U�;�g���<��<�W?;� =Sz��k�<�얼�O=�M5���=��=�	b��P<�<�y�=~S�<Ĝm��	м.������P���f2=�1�V7=k�=��
���U�0F@��>���`=<����м(���!��!}8=%O<=�\d��"=b·� �5�"��;n��<Ag��;���ȕ������r.�@�5=cI�_BI=�����Zn�N�<]c!��t弢�<�_R��Ә�o�-=C��<�q�B0+�2��<s��P��=ݼ2&��y˭��ق=7���R�<�-=�q���/��zk=�C�e"���O��,|V��t<<z	S=`��<�B���#b=�u8��0:���p<B��H�/=4��<cl��š!<�+<y)<Td;<}�;4v�hD8�pq=nJ��	��掙�$8I���ļ�>��~��}�=����[�<�h�����Q�F�X�H��x
�3��u��&\�<8�-=8��r8���d=�ur��F�Pe<�t=u�<ak7=]P2��C=�&3<0肻[�;����o.G=W��<��9��<��J�F�;=���<�@�<,p��p#=v�$��Zj�|�;�,+���Q=��b�v<�㼄wR�X=9�
�=�R�<g�	���<E�n<2�R�%���k2=� =fG=�Au=�����Z�<ƁG��U}���=���2QT=!;�� u9�������<�u\���B��U�V�^��"]^<�U�<�v<�L�s[5<;�R<�fa���<��i=;b�<�a��n�<��;���ۻ��5=�K�<�����<[$&=��m���D=SV=�4c�i���<��8	;�sĻ��=�<x=[����0=�Y<,g��;s�=���wCM����<�]^�L��/�%������<6���=�RA�⣋;�Щ��+�u_]=�I��mL���D��@j=���<^�<!�:��
;� 缝B�<!�G<��;c�<���=d�=<�k`�}-3<���<��;w�8;��.��u3=V��Z�e@T=��-=���<��!��UZ�fc��s��݆�����:�A�B᝼�꼤�=Q`,=y�
=�EK=��<�ƫ;���;�)m=X������;�#��<Q�t�}6�;aw�<}_��a��<3=�F'�:<���=��+�Nؚ<]i�<��\���y�`u�<�8��a�#�
=�>̼�2=`�<[�&���<�כ�BD=U�G���(=Z8���F<	=����/�3?=8�<l�<%�/�hu7<���<�\ǼA�#�lt���F=]�'�4��;�3$<l��Q佼L�F�)�����<g�˼��Y�$=g�+=����u��<x(=Ln
�}Ƌ��i"=�E=t�a=�5=�<V;a��0~c<\� �����M��V�<��-=ƇＥf�<�7=)E��?z<I�n����;\�]�)�/=�F�<#�y;YK2�H�&�K@:��.n<�j2�?ko��z����-=қ=9�e�ii���=�H'�UI�Ø�E!r��*V=̴=pT�<��;͓���l�<8�c�T4P��s!<����T�$=�֚���;\�=�N��A�<��>=ƌ`=��q<��<�vͼ�ʂ=�6=l�.�ǂ)=ox�']=:�
=�4�<��	��
���;��o=,ż�#��Y6=K#W=Tf�<����=��&O�<03��~|!<ĳ��$=�.=�v�`=�������<�֑<#�T=cA<�*�C=xP���?��m;=K���W�X=;����z�<�]2���<V�;͗�;�q�z|<Xo]� ߽:g���V4k=��������P=wi����D@=ءk�n_ż�R4�$vS=uf�;W�;k�m���a=1c<�E��p4���]=�i�moQ=�=4<3��<N�ݼV�8=�g;ˣ�pH�z`�8U���<�����:=���):+��E�~!�b�漿�-������ɦ<�/���[=��;�xM�����5*�*��<�T	=��*=��u<��=;��r��|;��� ��żj��<��a�mQ�F8�[H����;�U2����;=�����R�<�����	[<���v~���>����<Wf��E�	=SD�<�(�����d�SB|=��;�^?�z?�"��X��;Y�y��O��;�=���<%�6�b��<�X=�D�v7w<�.%�-�;���<W�Y<�/ۻL�-|�&m	�'r6� 1���t����Y<��8�����	��ʘ<eLK�tU�:��@��b�<[�ϻ=X�<Ƚ���u=wt�nO�ǔd=���]�\=L==��FT��ׂ�r�<u��H��D=gS�w�}<P��<�_`=}�=���<d�J���d�6���o8=l�<�5=u�?=k��pӣ<f�@�5~�<�n�<�Yy=`W
=�s�<N2��_IS�Q.����V���<�\W�<QE?=f�<��k'Z;^�����.=I;���<"c����\=����/�<3�_=զ[<Q=�@=�;X�:y=9v��3>=՟�;��i=q��LC$=ͦO=S[&�Uw��������<I:F�ۼ	��Æ=�5p=��9��4�)���u�
=�6@�)�C���>=1�In=�v@�w�K=%G=��~<sK�<F�[�3l�<������6��*=���wg,=�:�JX=9<=�3�<*L%=�	�<����ԗ<��4=D�|�V��<�K8;z�4�^�f=���>=?���r���I)<-�k��1�<3{�<X�Լ(��<J��<�%%����~P<$/�0閻��;�1�<�#g�U���Fd=��4�5S��GrJ=�y��x�^=&�<a:v=�L-<%��<�Ѻ��-��-=s�c]=��%=A�=V"9<ӥ�<߰�<r��S=k���(X;EL�;��<�6= lX�����=J��n,=�:=�6]=d���<=�;n@�#Yϻ1GԻ���<,(�O�C�
��<�<�袼?��<>3�AX�
=h:ؼ�˴�J��o�?�4=	�&;�=��＼��<���M"�<�jg=�ɮ:����$-=�$0��T�<cE�<t��<8"�<��&=�=�	<�M�c���S<�E�?�)¼/]Z<F��B�Z����C���B�3������&�f�]��p�;�FZ�q�;��T�9�<�K1���<�^D�b�<Kۼc4=��<�o�<�$%=
�"=f"�&�!<�;������H=�1 =�8=/��<_�'=-�:DQ_��¼�)�K�ü��U=Ȓ\�2=KN=7d(=d�T�%�>�=���0�������_a3�J��߽<�B�<�����V�*�4�(a=����݂<��<�R-=;¯[=��W�=>�<�]x���=�@;�5��qc+�ԭ�YϺ;vEQ��$=
���C��<�{=�A={�=.=#E#=;AY=�%�>ܼ�l0�=���s2g=!4I�,3=��I���;w���S&�.��{�K�K=V2�<�$�<|�;M��i��0��;�\Q=�a�`��<в/����<e:�;,k��I����o���(��I)����<�i����M=�O�:G�9�n����!=�u=�ּ4��<�U=6=�$��@��W\<��O=]=:�<�K<�<u?���B0)��ּ��@=밼�=��c=�
<<�Tg�`�{�9J=I���v���+.������n��9�༔�>��h=Q���C��<�<�ڻջ˼�,�<����5�j�����t"ʼ�����Υ;:��<��;r�K=�"����<+�>=a�*=�aB=�4=�Jû`*��l�F=�,N<\�&����;�����<d�I=s7��P��i�8=2�q� K�� �"=[�v�f��I#=EH6���8=Z>��\<�"��Gl</R�q�@���}���<3�;=��a���=d�^=}����Լk�<Y!]=��O=��T<A�=�Ky;�;J�H!���9��mA�
%�<N�<%�<�� �G۾<�x=:�C���6=�=�xu�~�Y�j��<�+8�@�J�i&�)Y<VB=�	x7��%O=遼�Ȕ���ռ�P=���<,�_����<X$�.YA�W�4�SF*="ﰻH��j6=�=�&��=y.����;��=�==��<G�$��� �#O�<�h��<^=ِ�ge=%��<�]=���!4i�g��<'t�<iZ-���=�4��I�9jl��2=bpo�,O�<n:+��D3<��3�S�<<գ<X�<k�z�%�f��,��<�<lqW�.ߧ�Y
d=N\���'=)h<��<���<�f��������<�V� ��=�%m�<��;O1f���S=E/C=��%<��ד<��=��	����.:�v�_�M :���ݼ��<Btռ�k=���;��R=�W�<��<�L=�_�J=��ػ�I=��?=�<��j�:�{��<0��_�<i����>��"C����<?6=��u�<�d�z0üI)�<>	=��.=@*m;�X�������{$�a%���
��;�E�介J=qP2=?�<��h:s@=�F� �;�9n
;#C��J7=�ao=�<hN�Z��� ����!=a15���<{?�6���8�<@��<��=:>��%�6�X<�N�9�^�D�<������<U�J=R�`]v<XJ:���$�<Z��ZP"<�3<�rF=���I3=6K=��6;��.�Z:)4U=�YX��o�S�<a�ټ��<��<E��<8j鼸N:���	EZ�#m�q�k�މ��W�:�֬��N��</�3=����b�*�N=��(<,�/P����D<$f<
=��r=�L��O�=����>�<bl�;%�m:�h}<�a=�~j������<�[�����=޼{���<��U=Rpk=j� =��=?�</���/��^:��a=̫=�ü�c|�_�<�����!�j��<V��< �=��&<@C0�k=����ܼ~=��hXC��A=�<M�=�5�*O}�9Y��G =��-���:��V;���S�g=Lj�S'�<Bj����E��,3=j�=(�r��<�?��l�<�"�!9�2�"�L==���<�e�<�5�/�ݺ;�]�>)k=\�_=��?���k����:4�J�{���J=3l2��B$��><��pM��Dټ \���F=�M2<�|�<��7��s=��=�)#=<'�0�B�'8����<\�h<*AG��E�� >|=\��<����Y�<�&=��B=��;<����O*����<�$�< s-�)8=�ʼ�'�:뼼P���#_=&
y<!XL=2}����<B���Q<���)�$;��=n�_�<3���7<΃�V��;�c�<x�����:H�g=�m��=eU=��=��H=�7#��[	=�g&���==_}y=�M=���<ȜE=j{��}]�;����<Ǵ�<�@=��Ƽٽ&�`7�^�ۼR=o��r��<�d=�$�CG�;Fs�<h=a�μ������<�w�$�ܺx�E:�>]�%'=" ���=��E;+�
�n��<���Э�d�,=��G=�}�=w��7s��c`���=��<;��;吼���<�q�$�T�YR»O+)��x�<�B>=�*=N��<�c�]b7=	:�t�<�
=eC����U=�3�t�!�lc-=���<��S=�/��������<��A�w"):<Z/;U%	��u�T+�I�<4׈<�·�YL����;e\���S=��e���=c<z�f=��<T'��ъ4=��6�*�X���˼� 4���/���G=��]�X��?��{G=�&=��;��=>�2�e^;�6P=�\�<t$��T/�bY{��,�=fʁ�M�k�/�<�
=4J4=|��<�I-��y�:��;��=д�,�={?����:�8=�����0�ހR=.�񼍫1�C��>��#0=.�D�>[;1�F=��n=5?-=dtV<5�<�ӵ�-�<)��<��A=W�Q=p�Q�ϴ���V;�Y˼oQj<����m��W�<�D��4=<�</�2=FJ��N=L��z�<<�?<��)����=e�T=Vc�og=Xu�;�r=�=Z����:����LN鼷�7�>n4=Sq�<��ܼI�!<�ZU�2D&=��:���*<j�
�b=XU¼-��<�7 �5,=�p�;^�����{�=�����Ŕ�yK�<m���Hr������tH7�"h�(�<C0)= 2K�EX=�A�C.�W=l�p�J���J��<��\���:{I�ɨ[��.;!a�c`)�6#<�!���_=,�z=Utc<�i$=p/ѼӒ�<�/=ȟ��,<�5��@��<N=�Եڻo"F���J��F�h�9����<9д;�V���=o��<��>�F�^���I�m
R�V=ݟ{�&�����l��� :g�! <�q�<���,L;n����R�\����<���O��%x���_=�a�:j�μ��<=Al=�%�<`*�=�"�<cN=0�%�D�b;+X��m�.�<vH6=*'-��9�ͅ��=*e��<�@3�̈́μ�lm=v�0��q=@�����?��o5�P(N����;�D�Np���(����Z�<�+Y�M�S=۰�::�P�=��;[߼4�<]Z/=?I7�{�(�Y��<���:,q#<�S��9�<�3=
�S���;/�>��F��O�;0����~{�Y�D<��N=�Ｆ��<C3K�9=k�@��@m=�k���X;6��Mi,���V=�/o=��`�<����@���@��|���o��G=1�����;�I��pɧ<�=�9Ҽ�"=��W���$�H�Ǽ�|��jz�;6�+=�,6�	<�`E=� =!̃<�<=�Md=څS��<cPI<�,><���;;Uɻc�$�h(�;��W���]<�#���J=��~=���g�7��:������D[=p�_<����廄W��Qi<�.�;$�<=d�<A������U*=��"�M�ż�G�<�珺��/�i-=�P*<{&w�2��<#�==W*�2���e<��?=�s2���<!2���Ἶ���'i�<!ꁼ8G4=L�=��5���]�%1ƼWZ�<�.�;5��K�ۼd���� a����<�X�<�<��j/ =�Z'�%�D�і���\\;Q�;Z�Y��J<�),��5&<���y=U�*<�S����<PL�<<h?��2=uY4;�h=G�R<]m+����;
1=�!)����<{�O������.��'6�^0�a���i1�<��}Y�={,�o2����<]�{=�rû_�绡1��fć�D]'=�e&����ƤݼGkK��=T�;�;�@!��Z��To��)�J����<,�ͼ�$=m���|=�T�@&^=k�?����|A�<Q=�۟�<���������i<\û�/9�w>����Z<��=��NE �+So�x��:܇=V��Xlڼ��k���
=��K=�V=�#=h���#�-��=h��6Y����̼�+;<7���<
�Z�#���Y\�������6=��,<4AU�Z���P̼h�=�|/��:�E.�W���&= �4���m�ǀ=T=�L	����;H�=%<O;C=*@o��Z<4qO=F�����.�r�z>=L=����5���\o=!OZ�f�<'g���r=�B�Y<�M�<��k=U# <����[=JTj�G�0�<���RN<��G=Z�==�eM�7	_�r�>��Y���r=Хx��9k��=x$4=�z
<K�=� &��r2��c���P=����r�!��g�v���e<���<b�(<�r������| = �<��k=��6�>���F����<��s�O�;S���H=і��Es�<� �<�yF����<��2�pwc=J�8�ۍ�A2�t�����!=] ��+�j=�9,=�mQ�<��<e��<�=��/���J�<�����7��.=o	'��;=ά�=�Ḽ��.=#�j���.��((��ϼl�m�)O=�A=���;��b+<ӪJ<��߼��w�e;%g����=��=]�o=������7���N�	;��`=��<�;�9�=�
o<���<?[<�6I=:�<%A�ePe����@M�<u�Q�/#=H�����!��@X=A�ü��L�t{ �y<����G=oz����@�l��<ڡ��z\�<̶ܼ�A=3=��=���<u}=��Z=�J��J<�=x��DR��N(��H��=L���Z�,2<X92��AQ<;돆�d�=#e��g�;!�S��	�D�ۼ��-=�-=�_b=�O���:w=\'��D �M�k<~�ɺ�|ؼy��ޤʻ̰�=����L%��=��,����<�O�k�4=ְ5=e���Cd;g��<���<!F�k����8=��?�=-
��c�<Ռ�;��N=%��<���[�$=:�!�N莼T.s=N�<K�n����]�8=i�����d<t��<׏��6�<h�?<cx�;;_�;d�����F��=g��ݯ<lt���ͼ]��;�-D=�b���=�=��=��<���<6
w�K�B��b�u�}<�ד<��c:^p�=�CP=F[���=�H��y&�<C�ռ]*/=�uL��W=;�(��>ż'ϒ=��=���(��O.;[+<=�sv<J�7=��l;e ����;�x�<� ��)�W=�
��J,j��Xļ��<K�k�	]��L�@�m�I;�D��4�Ǽh��<9�ټ�G=�^� �����!�h��<`n�����,���{m�8[��V<��~���=jࢼ�=��G=�/�����4�=����锻�h���ą<n���$;&�R=|��<��� =�n	���m��a�<��<b����� ��<m7�<�!��pT<��<.<i<̱���:�Ř<� Ǽ��?�&�����=<;��4^���=�J�Y=h���T<J
S�j�;�=?�~�P=�M&=���<�<M��<�%�ǂ���j�)�<
0[=��<y#�<��=^-<J$e��K���püfAR<N^��L���n�)=��:����wd;b�e��t�<A�ʻ�/;;��R���)�Cw���<���<c=����%=w8���p_�������Ҥ;Z�m=�<?��XH=ͥ<.L=(�<]u=F�i�L=VP����<�=gt;�ȳ<����/��<��:�_���d�;dT�0�<��<����U��/��<�Z=����=�C�<�kgX�ZL�<�%2=�?�;������de��	�<=d��<0�<
��0�V=(Ha�S31�G;	;�k�<�;q��;"S�<���;ڎ�[)�:T.=���<��r���#=�\����<�f����<�K����C'�� �<U(W=���<��a�{�=L�Z=�ʿ<�+_7�[_<���^Zo�\@ͼ��v���2=�� =Q��<X:<޼��������c���e;=�W�@=ζ��C�<�O�����V=(={�[<��R=<	�	U<_-���f��H��	�.=���<���<-4=���<0	�s=��c=��J��D�<�� =�@;��<9+��.g�AG��[چ=>7=)��<b�#6�f�9����==����z�=�2���==-#-<�f�q,�?���d=pp=s=�.=��\��"l:i(���ͦ<�%��$�E=|��;�H=�6�1z�<H����.���<��H����B8�{8�<��2�� H�I��`҅�ОR=�I���(�<�;�Y�<I���X=_UR�i���|t><�E���W�1�*=>M3��A�<xS<
���;�`����B���"���^�`�H=V��1ļ��;:�;a��p<�L;�n=��K=(BS��_������F )�;�����<_)�<��L<����Z:�C�t�����	�8=���U��P�\��9
9[vC���1�<�^�e<���<~)�;;��<nB���=�9i�;qOK�|]<�*�<��L��0E��6����<-Î�lM ��'q=�w�;2y�<��<_ȼF�V�r;7=���<H���Yt<��T#����<L��<<v�<EH����= �t�fּ:��<�򃻬�'�@=�m#=�`��V��;-�A�c
��-9�<��F��<�[?������&;(r�<B������Y������\��t�<Q����I��Hb��w=��F;�-�<���"=��=�ZT=7�<�� =u�<��(��q�<�"X<�?&=+J��BӀ=d*b�Ь.<1S��Y�K�U�=��<Q[)=5Q<a�K=���7{ռ�v0�-�=�V���e����<w�
��:�;�f�<jc=b�=�B�<h�=\Tؼ;F,�1P��_�@��i(�>}=
'O��y��}dP=y��<dMX=��=�[	=>(�U��<�SF�Ռ�<D�=�5\��^�x�<C�ƺ.i��$=��ռ`��<i�=O����~W=�1=,�J��N�g�w;M1�X=��^�*=_�+���R��}��EY��l<$,�\'��i�D;�oG�} �;X�3<�9=q9��<䚣<aNB=h1�uI�� H��k<�҇=.�<�܄��ME��딼�<�I��4�{�ֽ��U=�R:=����ʼw�<#��<�V��<�OA��uT<�i�<��<�A=��<�+��{�	���=�ә�W�ԻM�B�hn�V��@�������=�!X=��[��`�������!�d��d�<R��<�Ƽj�򻍡d��a=0=�!�<{�=��!��|'�[<}	=G�K=����.�!��(D;R
�:Ql1��-	<,‼f��<T�1(U;�/׺�?=��S����|�<Mb�zuH=K��<�8=��G�y�<�q�<	�<Q��<���?q��ux=;Eq<;�ݼ
�<�2=�ͼ�]h��ع�)=f*=:U7=�d-��LT;����Nm={!�=.6K�)0;~kt;,�-�z=�<K�_��5N=�';���<+zo=�1=&���$�}��/a��w�,^=��=֐H��W�Ԙ��{&��=D�<�hѼ-��;MJ��^<�ߕ�I��<�[��'�H�4�I��<�8D<m�.=ꇼ3�0�FR�<�s<�B�PY=�T���h�</�ǼԲ+<n�:=w(k�3c4��_&=!�<��=Q�i�7�><��;�-�u��<�ᠼ��;��<��=��m�
�=t�F��㼞=�]!�#;R��xԼ���<���:2k��W=��L=����r<��ś< a�X�H��9=MAм���<�YO=L4���Լ7t�������:0� �d��Դ&=-���I𹼗��<I	=����`q�A��<�x=�}˼�*=��=���<�h=o�_=VY�염Κ�< �&�3�/��!�-Z><�,=��;g�Y=m�ͼ�޼�S�<Q�={���:^^�-=��׼�=g��<��<��.���<WJ|�S���LT-=�eF��j��:��2y==�dO�ǧ��@!=~x˺��캱�<~GM�6��<K��;x�\�YJ`�jGK�::͊ͼ��.=Y�"�=^�e=��=쳍�\��<�2H�;����Ü<� =#w仁��<7�=�V�<7b=*�뺳�J=��=(�m=�/=їN�8��<�!0��L�;4һ<��<A�=��7<"޻:�h=�K};��U�I�<t�`=��:<+s��`0�<�N&�t~�<��H��k�<D����q=�%Ի6�ڑ����<��d=�uR��rż�t=��a��j�;:�7�Dn���6=�H=�v���;)=tOY=f�/=����H�R������=��#9�(��⯊="�T*�;-)���ỤKX<��<��ϼ6����<� ��p��q4ۺ�JW��:?�.輖���߼*�w�$��<��B=զ�$<Ѡ?=�ȥ���ɼ�?��Z�n�< a,;�Kº��<�*��z�ۻ.�Q=7t�=�^����<t��A��q��;H<�=Ҽ%���Q;�c�;���Ft�<t���e�=W3<utw��)��v��K�&��I�m3=����s�<}�+=�5O=9C���Y��
6��;-=jW=|Q�gi{�8mo<K��<��<4J��EV��z=B=���-���hi=��n��8���<Y�<9���A�� �[�V<!d�;w�<3�^�L���bX����F��#�<�=����[���<�Kټ��+�_<Ta�<����m�;�i=\ =Űۼ��z�\�=UCy<\�9��E�;��{=ʹ���p#����;���	�M��7"�%�?�b���w3=tǼ k����E6=9P=�G���9����<��f���OF��0�<�e���)=n=I=��,;F(�v���U��<'����ڏ;ww�}�?�2����5*<�"���̼��%=+�ͼ�;=�*=�[-�!�<F���Q�B4��8�=�	�<gJ��n=~�:��v�:Wt=���<&~C���y��;c<7��3弪3��O�<Z�<�W8�����5=u�:>!�l�<�U?<`�ؼs��<�=G"�<��7=lKh;;=c�u���ټ�=�V�gZ���V�n�v�^�e���B�jQ=�[�=�����3=~�-�M�;!T��<���<V*w=�T����#�S=��酼���gg�4��<�>��q�<%=�e^�R<�<��<6�<���\8�X��{%=2#���k=0KB��U%=�Z���j�<�-�=#�,��p��M�K=(�+�;]�����<��=��sż�%D�\Eļ�Fu;H�:=&Ku=�ʼ>���/k��Kɻ�1���=|��5y1�l��<��*�𞦼�6�&D=_T9=	�s=�AH=�px<G{��a=�b�;b$򺠿m�8"�� H;eC�.@W=u <�e�#�=R=b���$�����=���<dj=���&�s�z��<��$��@h���@=���<}�X�^vI=��`=WJ�<�x�;
c�<�=K7D=��0�sU����<��:3�>=�=F�_���(�u=-�:�B����9l�Y=������0={9F<���<�u=�.�<<L�<(Gj�Dd̼���<@���` =.���/<�C���J�Q����Zj���O=��鼥+/=�,��;&�-�	)W<4m��ɡ;Z��ƨ��'�<�q-<�dK=��	� �&�;r8=�O=�)�<������=���^-v��L>=3S�3�[<�6;�\��L����;�0��P��<�_�<��߲�$9A<%2Q<�k@���H=x-q=�`=E�"=j����{�;�(�;���<f���v=9NW=��R�Fʻڍ<�g4=��ż�H���<S}�	��"9�<*�K<��R�;=�t�=�2q<+Rq��s=চ����;�.F=Q��<�('=.H��a���:<0�U<�S3=G3%=��ff.=��<��'�ǋ�<˒��ǩ=�u��~c�w&�#����fG�<$�\=lһШ[�/O��3ˈ��<D=ٓ����<7}N��V���(<MJ���+���M=|�<nB}=�1��]�o�9��"�<"qf�n#�ނ
���<%c@=R���|��;�J�<U�Z�=�<B1�<5��c7�V�<v_6��Z<�K���-�<�*������I=��M=@o��% �`��%x���)=nN=��[�RW<�}�"�E�5�F�;;�=�+<��-=Li�3� =��:��7�K��<L���`�Y������!?���=��n=\m<=�?���=��9�<zr�<ʬ�Xu���`�<H���GA�i�Z��D��8<p���`*�M�����<�B]�yc�;3 �1_<=��<�>�<=��r=��M����Z%����틙<�N�<L1��z����0=�e�<�G=i�0=ʀ��S�%����<i���X�=cT����߼c�{���0�f+���P]=�����DF���<	�$��OӺ���<Q=if�;�8꼿��<�B<8q?��R����;;�<4\5��ݼ����T�<>����1�2�<����<�<��O=j�m��%�2������j!=��<���,R����<�9���h޼j~��2�����<=��Z������|�I��<�4�;Đ==QZ=����\�:���-�yL�F䞼�����}>��;={!Ƽh�F<�rE���}:4
V=zȝ�k�<{+���ŵ<�>�C3<y�<�	M���M�c)�=�e��� =�Or;N0c�R��<���e<���:%��;�c��e=�[�vLR�L`1=�Tl�&�����w=�j�;/E���<�%�/"�;	tE=�JE=lr�<�}_<�l�ǹ=���9'�[��;�
7=�{�<%����]=L۲�A[><� �m'*<�u ��l>= <�����/u=BI@=��:���:������<Y�ܼ�=��9�xJ��>��l=i7�]��<]V+�	�M��	�:�U~=G6���a<�j%�)a5����JI<��ڼA�ټ�����)=`�I��g��w��w��So[�+�;<���XK����<- �*�@=8�?�9��<��޼����K��<E�^��"��ʹ�<�~����=O�^��lü�Xu=U�6=k�3=���<��J�999��@=}~3�NE=�<�[==�?M=gӅ<�=A���廼��U=5�����=-4��ZrZ��ڜ;�o��4=�zC=I�<�U\<��<8��ω�<-/���-#�T>�<Pb�=[C0�h��K1 =V�ټ�7�������ϡ��=hH��:="=]C�4�ּ����w�;�}�<��=�9�q2�;\L=�"-<��H<�֋;V���?o<0� =�$)=�#�<[�	�̶>�CUU<�� <:�@�+�;�.���6=6ܗ<��'�1)���=�%8��'�<i��:�컼�WT=�	��&W5=�2I�����tQ�^f0=���<�y=��N�.El=j<'��)�~
+=���<�7��e�l<��U=!iD:"(��eK;�M:���_��"Q=F+L����d�4>`<�Ή�昅=�M�;��W�����O<Z�L��*<������=��/=�$h����<��;=ӡ=4=W#��ꍼ�J�;��.<AI���B=yO��!�Q=�Ue��<��� >=�-F�R��=-�D�L�=�4V�A%=�0�<N��<h�i��<yӊ��Dt<!ἀ�]��/<��W��Y��9����*Y�F�:����Ո;���';��T��O=_
�쬊��-���^����l�=۔M=��R;R+�<���<B��CiS��
����n��X�7��U��!��;&�G��wW=��'=@w>=B�Q�8dP<���:vZ���O�;u�<X\N<�6�:C��}��H�<�����+�!�T����;T���Jɼ�-=x!�:�%���=��<��=T��"C=���<��5=3��<b��␃=|�w=����:e=Q�<|�<.y9=�'>�G@���w�t��I<w�����L=r�_�=Sh��w�<��X�@<мE���U\�t�z����۰�<�9=��!=��ϼ�ާ;����dn��N��A�84�ڝ&��$J�y�>=��*��\s=���<��=�)��b�<#ɼ��p=�h�<`�S<�쾻���E+�<�g=�Ly</j'=�Ï�ox�TG)=Q-�;8�Ѽ�g<-�z�5�Y�YHj�&31������0�<�ռż�b��o=Uu��6Z��>�;�	i=�*�$�&���<I6$=��><~�=m;�<��{<ǐ��!&��/S=��4+
<y*}<�nd����<�C<�~#=��μ�<����)<ɿ��Z,輐�,=��	=��<�=�$u<�Rû@K��|=�0`�OZ=����z����<8=Z$��4�<v�<��*�6����`��J#.=�&�:b#�䊼����t�?�˦-<i2a=� �KT
=_<f��?G<&�Լ�LC�ڐ����w
������Ia�߶D�]�|�Wd
����D�<�w���<\��;hn��͉K��:.��ջ���<�0���S���z=���<&���#���v< m��%t����һ�<�o��<kO��=P�M�׼�U�%�,=���<�Ȃ����<�*�K��;s�*=��=`���AU��ؕx�o���F�ؼ����(q ��D$=,D;�Xa����;��4=���<S�<�t5<�"=��6/��e=�"�<�u��И<��ż+p��
���<m�,��^-�"�%=v���<W�K�=f��<�j�)O����@�<�߼��2=tY<�鳼yo��=���<;#N���d=��*��+���o<9�=����k�;�l?��_U=��������=� <��x<U3�8b=��ռ��=Ĥ�:}`�;ᚮ;?��<NtI�h�V<H<����<m��<�J$=[F=�w��G<Z=l
�=��8<�-�=�x�=+bP�kw9���_=�K��v����><20=H+�;���uш<2��O�<�kL=y:��m!H<o�a�%�<�
G=5�l���c=�v�<�Hm��$<�x0=YES�ǿ�<�PC=��=��D���=���w��Rb<�m�;b#�<�nv<�NJ=z੼iCq������u<��s��u�<�İ<Gu�w@�dc=���?�>��<�9����<�^�,܊<D��<���<*g=��/�bN�<�z;��!�"=-)�:����g=f�#����Xb�=�KB�,Ȍ�� E�E��<�0�<a�.��N��dm	���;�8$�~$�< ��<�»G )����;�0X�ȡ0=	����={����OG<�.=]=	=�Y=N�+=���a�����U�;lLF<Om�<��>��pG�Wi/�)��<"��~�׼my=ɩ�b?=2
�<p��;�ȝ;В���Zy��:�3==o`�p3 �6n
�O���^E��@�|��C����=
#	<\�4�1T�h7�Iz.=�,���a"�#��<��<0��<^�����<���/�A�*i ��=y
�2�$�ѯ;�g:<�>z=�j�=��ѻ�(�<�)}<��F<��=��߼ưt�-��������e<'��<�㌼�@�=�<�!ż�m�=@�\=pc&<�*8=>0��ME����S�n�%��;h�F��)�;�*[=�)=�;�=�kl<	�.�;(J�<�SY����;��Uz<̓��K4�=8{����n��P���`R��=�A��K�w<�Zڼ!��<�F�.L�<�''�n&]=�.=��ջw3B=w[Z=��=�v��%$4��E�<R����$��u=Z$�� <Ks[�!b�;9na��Q��	����k���X;)��<g3=�g=��Ƽ�㧼�e=�̼�@:=kF�<m���$H= ��=�bH��:� ���-:�r�=IR=�l�<��;`qU���/=%Ҕ����<H߼�]��n6���e:c���-}���OeH=6�ռ��<N6=�#�j
�<�x�����L\<����-%�9~U=ҧt=�W��JʼBA]=@��ل;���;��=���=`�q��I�>� =���:qL}=H�X�&��<�3=A�R��*h�K�#=�=.=^-�;�3�;R�	=]U��$�	��Z��ه����<}U���⼘Y5=��L<ŵ�s�/=$��<(,b=ltF=��+�s�^��sj=d��;چ���0<��]=�gS�⯅=p��q�H=.=�1��|2=4�=ǻ���>��^g�<��s�W�M�»�H/����2S��븻ȫ=� ����(=V�<~t<e�O=!�=��G=�
=w��=��Y�+�O=��*=��<��<lꕼ7�8=N�=�A=Rj<=�"5��.�!�.=C��o��<[v=(�����<C�o;���<0&(=�T� �9;�L�=��W�0�+=c#a���Ҽ�䃽�2���(,�?n=Վ<�=ϩ鼆�*Í;�?=��E��g��b=�g�=�z�;�YB��;>;[�="+=̽w<�E1������=ɃA=��<��ғ���=���)�#��ټ̎e���=�qq=�&C�m^(<=��;=��=}J(=''�mn�\�� �<yl5<s����>��
=��R��=���<,U=�>Ƽ���4!=��=��<�H���=v��XrA=Au>�C��}d�<�N.�]��<Q�=
}�� "{<x�=��1={����h������:;�
�;X�M��ڡ<�w�i��ׄ�@m޼�[=�rA��{M���;q=�EQ�d�*���=��-L=Ps�ܺ<c�<��j���^k=��=�=TcU���P=^f���m\���=�G���K�z���0_�CN;ަ!=�{<U�=�\����_<|	h���x��yU�&�=��e=��=�H�⠢��}�<Vt="� ���A��@�=��a����%R���=k5ݻmΩ���5�{�d��fٺ+n<��=��<f_<?�����<vyY=�"�D���Ҽ뼇=#�=<��<��=��n�*=~�I���;R�t�8����=�؀<�t���F���F=Rӫ<7�==rPh=�=�<�/=ַ���;�wE�<�༮���eG=���氇���#���R=����y;�P�5�;�k)�gY:��<F�<i�G=$�~���<��<�$<�����=���;&׿;0=#!�<鄼�r=d�,�9��<(F@��w=J���4=�{P���_�_�Y����;옑<��<x�;�����[6�� <��2=�{�=��:�QT=q�`=L:伌5�=b��ݩ��Ҽ)7a�u����Y= F=o����&�����ʁ<&4ڻ;��<����2��mV=�N���˼�R=�4V�H����j.��nK=�;���7=�]�S�<-~k��<&<=�~@=B�x=>�H�4��<��9�P�<֠��a f:�d��(�<��;�܁=֬��` =kJ=K)�<�\`=:�X=��K<�1һȉ<�I=I�麆��YZC��)�Pma���ټ��L��m�<�<�.A�\��Qm=��=h"�;<��<�#<�9)=���<4�<��;=�q��IuQ�P��;�B�iM�<*%����==�o>�VV=v�Z�AF;إG��
.=�U�<�US��pE=H`N=m�Q<�>=PU$��	)��T���%��a<>�;��z^�L��<^4��&��<��<��
��:S=��_=��]=k��P��k�=��ۼV�r=t)=���<};�!��{�J=%W��{�<pP6=k�<Ż$P2=��&=�l=�&��1�V=�I,�u���I=+���Lm<c&�r�V=�f3���l]=:Fx=��R�|-�<�=��\�[n=��8��;=��<K"T�q�������9�<d�R =���k��f�;te:=p_�<��h�Ag=[O�?z�<Ns=�F���3��2߼��	l=�nl<`3���5Q=��I=?�N=�@�<t}����<}IN���;�fa��+�<|߶<��4�6��B�S��!	��� =�v^=��p���<4�$����<�B=/]	�:ͱ<栗�A
>��៻מy=W�[=��ټ��<�=�<u�ӼQ�;�ӵ<X�躺Z��
q\�d�@�"_�<�0��)����#�$
�6?e����`ؼ�&�<��A���u=�v=��z$������G~Ӽ^�Q�%��<�{��91�I湻�~�;��N��_��=N+=��=dx����l�ڻ�������
���l=:�U�I)2�M)%;K�򼬒U<-���A=�������q3=�M�n���m���0�@�=�)=���ɀk=O�
���G=��o=#���jD�8��;Zw��}�żf�X����<��>�S$i���g���r����@<7�e=�6<�o�����y��$�
�x�V=S={�<�I�<������<=�@�l��]�b�i<������a���V=N�(<��{��V<��=G����<�o=�Z�"�!�#�L��,����M</[�=��=��Ƽ�"B��d�'0�<\�=���O�W=�Ub��[P�h�)=���<��:=�����e��0f�أ�<rFU=�2Y;�<=	��<�=�h�f��qϼB>;Կ�Ф�<=�<�o=��V�J��<��)�5=��s=�&p=��ϼ&<�N�=��8=��#=	�����U=בt<�=��h�[��<2�<��=�	ϼ`�]���2;�Y)�X�T�L��V<���XG�<���8F��JD�3�=��=�D������8'���K����=CH=!e���@�F�<�CK�p�U�m��/�M�1%�<�<��/Y=��q=<��<�&=y�r��^�������N�{78=� M��.�`Z��f�.=4���[���O:Y�R��O�=�s���P=2��Fk�)��<����8�<��D�wt;��k=�9=lT�����$��_߼�2<��<^v���%=��=ٱü�)=�aE��߻�Y=J�><�g��]I�6��<$D���e�rO;��<
-<�*�<�]�=C��;P_��ϐ\=_��ώż2�<=��7=X[�e)=�Q=&�����a\Ƽ��;"l�g���J����l�<��$�����3=#�;�t�<v�)=y�Ἄw]�VR<��;�i=+5I�	��l�;
x7��	,�@�p=Y�<��;���<�Y�R������Ш����:�=ӴP<��8�HKC;oA,��D�t~�:���;��պ޼��;�S�گ�<|�˼Rd8���=h��^B|�`Q��ރ�=��缜�f�ZWj�*d�� �<e�;<�	���SW�^�K�O�8�AZ���<�^�<��ü�I=�>=��F=k�ļ���<����s=��������f��f
�ut<��D�����I�p��U��
��v�\�k7��ۿ�<��`��Q��^�=���'�����,�w�ﻂ2����V�l-���`-;��S�}6�;=��=MŻ:���� ���'=Y��0T���$=U�=��<<�ؼ�x;:�u�<7��<뵼��=�3�"�B=�G<i��2=��D=�'E��. =?^�L��<I��<.A(��m������I����<i��b�U���q=j��IlF�2A�'�����8:}������o=���<-��_>#��Y��:Ӗ����P�]�� BG���*<�,
<aǼ�r��$=�����<E�=/�/��R=���r8����E=��\=$�M��g�<Z��;>��<��1��}���=��=��s;s3�?Xl�?`=��9<]x���R=��9��Q�'Uq�Qi	=b*=���d�un�=��K=n�<��B<��P���=(v�;�D=2�5�@z<�{r=n�<C��:m=ΖE��z~<��=��<��P=6�=�F����3<�I������`n��)�<Lx�a�<��ݼb����A�('�<�9;��D=��4=Ι��=9�;�޼;�1=.�=�T��|s;�=V�C=��A=CȐ<VY+�<?�}{r:
)a�8x����i;=�5?=k�"��bػ/�<��P��'J�0촼k�<�J��p2�|��<,=��)��&˅=����#7<f�E=fkJ=�8=.+f<*q�<�w�;r�A=SIC���j<�9�<��\���1�'=���;�r$=�у��K���i=���ap?�?kN<r� =�@�<)��<� ��ub=�N׼{k4�&����W�S�<^�a�W�<�<��FK=����%�<*�;;�IY=�3=1��=«,�	��<����!=h=�n#��8ּQ}����9�2=��;���<�'=m(3=$A=��H=L�?=-=ʎ)=�8�^�<�2"=vL�f��<�����O�t��<�(�
v=� =�`�<e�9���R�Z�Z<�GH��a��['w=�*�<�ކ�,$�<��e=V�;F�d� {�<V���CB.��hE���=�0�'�<��a=������ae�W���J�h8�e�R���޼��F�)O�%};]��<��t��[�H�;�0�;�����+�V[Q����<�<�1@��ɼToP�!L��6�<'h<��6�����4��d�;�76� FF�~*�<D�c;��������\��Ll<R	3��6=4d�<X�=�(�<d��<�M�<�zs=�t[���)=����"�<��B�'�<�����R�{�B��dQ��yF��j=�J:=�GJ��)�i}�<�G��H�Yп���7;�j�k�=�a��X� ���4=��?�����yw����f���=n�ۼ�L�-���>��5�;�����ﺌ� =g(;���<�)�<��*?�<�;g��u��e^�Ja���>=-=���c�<���5d�3�M���h�gdI�"�,=~Z�<�ab=F��QM<=��y9\�*�0s���<�!A;��;G�:=܃��������<T�Y=����<(��<�dL=��ƼOy(=��X����aB=?A�2e���į<+�;��;=�]	�6I�<H�`�F*���a =xv)�����B��N���'�<X�8�{�e�=��� I�u�A�E�=pn$��v�L=��������׿༿���%��<lG.�;�_��u��5"<�$�� ���=@A=8�;����Ȓ!�f��<0"�<�k��_?� m�<���<��w�~oʼ�V{�)<_����A=��h��ռ�]�<��0=��P=vI��ﭼ�=S����;�b�<$Q����=��.S=*uǼ/};=P�$=ӸE�<�$�^�z��|�<��7=>�g<�59���7��u2��+;�0�!=vGq=Q�c�� �u�μ fZ��`V=�-=��"=��5_ =���D�8���'����(4<h�<C���AҼ��=ilR=��M��B=�@=9���*r�:@�=uY=��N��)�<=��Y=�}~�$)�u��<���3�<=��;Z�*��t2<�C=A4����r�=6�i��5&=�E���<��[=�¼�-l��=]�;#��gﻘ�;��SD<�$=�@�;�.Z=�p	��2y=fD�<��-����whM=.1��
�^����J���;9��p<�U�G�&�.p�=s<�I��t=lu�;���d�-=r�4<�;=�lɼ�7�<q$�=�5�ֺ��9�=��q=�Uf=.(=�%�<iJ<�=nނ<�0�;�KU��'��Nh�`g/<��&=��=Lu=>�!�\��;^WI�Qq&�
c=�+_=�tS="N����޼AV��;�ӼGp�<,-=�<ŴT=��;���%��&~=�D�����
�<t�U���
=+yn=�'=;�=��c=F��=#H��V`�,!R���%=E~����%���3ۏ�
z�;ϳd�w�4=|�>=�_o�����w�<�9/�	�B=g.=�Uq�V
��\�=�H��]W=Y7���=�b�<�I;���<���<��@=�R�:��:2��Ώ4���3=��b�<��<W+ �G�3�CM�<���<��x<�J'=�Y���+ȼ]��e�<��ɼG�,�UǕ:kݽ�t��K�<t�L�z٦<������@��i�<߹E<R#>=��H�6�m�ݶ=N85��1	��e��'ɏ<���<�Q=�
`=Wn�8\-�����p���=%���{�<�G=���<Ô�<Wu���M;5�#�����=��v=D�==���D;�ռ-���<3^8=P�_=��@��e=�VY<���%Ul�P'e=�:i=�D�A���(�[��s뼥Ur=b�+=��:!�;�A���.S���T�j(<��*<꽫�'��?<ҵ<�?���JI��c=|��;Lv=<� �<p[���(���<�3�@�[Hk=�	��V=iF��%G�����}<a3���1���n�G�9=	�0�y�V�P���B=�� <��1��;��:98��E��FT<���"߼��=�����b����~�3=��%�.=�^U�m<����e���V���<-���,�>��~�=��=�b�<���	 �F\ =4�G�i,��x�<�\=�����<�	> �9U=�ד<E�"=0B=צ���^ּ��=^�=�@=�<���.�;�������t�� N=�s<$�H�9V[=p	=&�:(c��j2=\�<$�c=jm�<Ⱦ�:�^ۼ]	#��l�:,�P<�� �8�=Z{�	釽d�S=J.��� ���?���=���<��Z=W�]=�c\��yk=���<�-��x3���_=�\=���<�%���������<S5ۼ�wV<�x�<��=�`(=S�X�FM=���
Z<�����w;i��;�}�<����hR=�z��2<p�};cF<nZ<������<��]<��*=���<��ӹk�;y�Td$��K%=�p�;�S=)�I=��<_����M2=.�ɼ�F=ȪM�W�;Ro�:��;%�=E%=�8����<2TƼn����^<��=�h3��ͼG==��'�HL!� ��<�=�G�<�Q�j�/��[;�*|�`ye�-�<�S���`u=��@���y�=D놼Mߢ�IbY��m�L�:=g�S=�ͪ<~:���t��_'�+��;����ͼ׉#=y9 <|#=���<�׆�.�9���<!�ϻ�!?�S��V�:��F��9-<u��9o`��4ٺ�o�<�ZZ��Z���`�禩��8=8�e=?<=Jl;��<%j=�f�=�(���*�,�Ӽ�v�;���<�h:�� <�p�ҿ����<�����=��ʼ�����@=&��"�p�Z�X=��2�hp=��q�<c�=L3<�;{�!=���ܘ�Ѱc�5x�<>�=��b=��E�n���L1=�[���=��=�{��^F5�=qݻ d<޳2=� <g ����ؼK�/;�A7<flR=�N�l�k��)[=@M=��j�����x<�5�;0����>�̘�<�Q�Lw�h,�<@ш<!��<�d���v=�0@�̴������£�<��<��<��R��i=������e=O�����<�3=2�f�6=}�<��><:ݼ�=���<�l���V=s$Z<�ʼ�jxZ=o<4=��"#�핐�oz�<C���Ѽ�)=zJ��)/���I=��a�w4�<0^�<桹�~#ּ��>��{�<(^2�5*�<���<�rG�Ekܼ��5;S�:��@N�3������R)��޹;��λ%��0�<o��;g�+���b=Uh=��<b�!="+�<+h=X�M� ���E�<�{;�8=�s�<E��<[E��&�źU5�eѻa'.����<��(=1�N<���.�<�(��B=u�<�h]��=�P��t�<\i=Rx"����]d&<N�<I��!��d�<�W��=� �<�n�<����my����A�t`	�ʔ@=|$����l=��=8��.B0�Aoy<����'MQ=�u ����<&U�<���<�Y�<��$=����MD��N=m_��jP=��<>r�;�)�<�w���;�+5=�aB<g,=�=�	=�k=ߍ�<�͹<^iƼ��[��0�!�&'-�]�:A�ټd�<�S=����z�5�_<{����<g�(� =���<�x=eE��jx/=TJ=�\&���ȼ�p?=wg2=����ǝ������8��Ѽ�叼�G>=�o =��4=�:�<� �9�L�O�<�_`=C��<��<L�;#��;Ǚ�;5e�<��7=���<����2��bs�Lm�=�Z0�����H�ۼa��<޵ =Z�E�NV�^�ci\=r<�ZŻ&�m<æ{�մ�;�Y�����M=��_<��ü���СC=�c���<U'?=��ܼC��<� �wЙ<���<�$h=u��;���;(�O=۝$�P;W=���V��<6'�;��
=P(����F<o��<��r<9�/�ɼ{p=+�0��!K��~�m$�?��fB���/�K�<3���o����=�)=��0=X���Z��� ���- ��ٻ�=5M4=�&�<M�=uB�򆘼�0T=h`<ά�<��<e���
&�>��<�H�<�c�<9$S��<;m6û�B�@w��<�+�W�<�� =Fu�;7-�%=����6�<��i<`�[=���<�҃�1q=:
����n�=��;��;=�DT���<@�"=��?�x���/�So�:JԺ;������<#�f�/n[=�U���l���~���<�-9=�;=hڼ�ʜ�3삽uP�x��t��Eڛ<�`��!/����K����m:�=�?
=qz<]o0<�Ӽ�2�<��û3�3=e=|SX�۟4=.�1=��8�
>[�3�5=}/���܊�zD�<x�=A�C�+���|�1������*=��;Ƚ<hk<���<�5	=��z���<|LX���k�M\ڼ�Վ�⒉<����+���(a=��Ǽ���=!!�ƍ�&?|<�8�<��=��N<p��kA!<��k��rR��':O.=��U#-<��=|݆��=< #W�̶~=Ș껻�j=+�,=C��<��<;�z=����<A�<s�'=^eB=�Iy=N�(=��U���t�����Ja9O$���m�*N���:JH�<43=�Pr<�=qUc<��)=B�s=]ˆ���8�k9S=��<Ӹ��P=�����<�_�c>�<�*�<I��<ˀм�<�g� D=�
��H)=	�J;���<"�;���;���ku=�L�x߻�3]�P��TQG= A,<�=�=;��a�<n!=�BX=+=�=?s@=�&�>i�<��i=�R7��N�<�?��k<
Έ�u�:/��J>=�8�<���)Y)<�8�<���<$�l��r��#�<'<��^3��m�=p�k<#�=hFw=R��<9{1��,�ࡩ<9f �l���H-��ö���
�U����-=�0\=:s"=;�W�w�̻�j�<�ƫ�/�<X��;�jZ<�q?=L�a=�X*=)g���e�`c=���<��ּm��<��<��<�\��Sv�V��</y9�2�E=/�?��=�����뼠�J��m�<QJ��8�;.F=�
�~=9�1����zU=���<X�ռ�7���,*��X���F<\$�/�1��'m��3ػ*�);�C�<�7�<�f���b�=��<ۂ����_=�7�|��<bg0��N;��/��
.;{_�;�T�<�h����q��$�3�ǿƼ�T�<�g_=fY=F�=�H�d�ּ�-2�ة>=H�O�E=L��;$��J��<K��<��Z�H��<�3�<L=O*b�O��<1&��vڼT8��!����\;��#�C<ܼ�����d�Ϻ���;^�\=�Es��i�hA2�1y�/�?=��t��;��H�Ｏ�^;-H&<#��q�����a��j�<����E�ɵ��4y`=�+`�f.=�|<#��^��;��O����<H���7�d�8=1E|�l�u��Z=�\\���"<S��<SD�;�钺_�μM�.<"R=FL�k��^��<�����<j����k=gT�M�H=OAe<�����Ex��="�o��h�<�Qv���.=�H�N�_=�e�<��Q��k���J�/i|��/=IX��|<<M�Y<�������Ȇ<���>n=�T�G=���<���ۂ;����O�dc����D��?�<ʦ��lP=ǄU=ᕼ;^�)=Uv�3{<��.�1�����<Α<,(ݻ���ߡ<x�Ѽ�ւ�EPż=��:V���޼���;H��ބc;_{8;lY=�Hc<�N=��nJ�	��<�z�=�|�<f['<�1��tu�����]���;?�<)"���ȼlU�<,04=/\��_���C�`�?J3=4or;�;�n\����֡�<��@<_2������Q=	�:�G=D�A=u��<�>��&��<Z�M��$�MH�<���<���F����=_$Z�L�����<��=i�;_�*<Q��<-���Y=�%M��V;=��#���=��[�^�<H=܁;P��<�c��vZ�C�<���;���y9i0o=�p8�-d@=��;o�=b�&<ӎM��.�=��=��������:��+���!�[�<0)*�d�����<""ػT>`<I=��F=�5�;�F�<c���;��;���\�A=����I�m@�ʖ=1ۛ��(�7�;渀=���|D����<���<�c���p]�Ty~���o�G���߼UF������{=L�Y=�����Aܼ�G��,6�<�W�<>�-=�m<�	�<�){<���=�¼�������;�2:=�v=�� ��#=4:�Y���{�=��9�� �<�"=\�<�|�L=cP=�~4;m%�nl�pQ�=#�����=�b�<��=S ��b3w= Qn=k��<�r�A�N�2hc�(!���;?�u=�#�G��;T73��N=��G�SG<��t=s�<�	����$<Xa�,l����v�==���<�at�R�L��:�<y�����c+==�RZ<�ib<�˃�la=;]���$<*��9�r���f����<x$/�y:=���uM�Q�׻�M|����<� =�B=�@�<FhY=�XR=�n��� ;�qC�v�]𐼃9���݆<�Y�=�j=���Ju�8��O����:����<�I��[o�<��X�p�^=��<����<^J
��<=]\��O
=�Ϙ<�Ѽ�/����<��G=&>�ϥ9�b��T�����<,�d�L�<Sy�;���:��b�]C�<��Q���1�1/���?��Q)�p�M=�<��mMt�|�����<��<}�G=P���~�y����<Q�;ĝ_�Ӈ�<-�������Jp<���]�;��#��m*=h�@=Pg=�c�<Nj�{�<��N=��I��
[�8p���i�Yʼa��;�����Qݼ�-�L�=`������}~Ǽ��λ��u�w(E�����	����Ԁ�<�f�<�ͼ2�)=pJ�=�)P���p=��S��4��r^���EK�"��<N������3��=ڰ�8 �=AN2�O��M� =�(�� =1��<I�P=X���e,=���K��m�<�HU�R�<��=FV6�<�D�A�;�6�<e̊=��=%F6=N_�<B��+)|�g��;PUj���U�9�d�<�Jl���q��<sm��8��E6$���Ǽ��=��<�9�<c�Y=�M=q�&�[Hb=6��kp{=�６��<n�8DH�l��<	�=���y�R=f^�;�(�Oǝ<B�H;R��<�[0=�[�fϟ��ĭ<S	�<��)���<�p¼*W�.�Լ
k<�ƕ=wF3��22<�Z)�IR����O@��V�=��<��=v�<$�t��x<@=M�=��0=\�=
��=e��;��?�|P<���;8@��Ћ��	���<�1=�"h��i���V<���;-Td=?��8�7�Z�^=��<�!=e�h=��:�	�<C镻�
�lT���4_�\z���ʼS5=|�%��1���#����h�^����skͼP�2=X�.<�>r��83=�sj�45�<��~����<��V��˔<L�������5L�K�;m��<=��K�m<�ܒ����]�,w<ɟ�uW{<)��5u�C?9=`�0�"���*�V6K����<;wn=�gK� ���4����<M�}:wA��`�a��*O=��W���R�Po<L�<�~ ;�h�=;ʊ��]�<>�2�׃�=x�4�|��<�=��=���<ׅ~��Z<��<'AO�LHE=<�0�c���=��>=-}u��m`=�>�<gY��
���y�:�g;�QI��4�;��<��
=�9��?���:=�=��=�Lٻ5  �mf�;��<B>���ac�%��<�J���5�����S�_�����p�⼬�N�ˋ^<݈4�b���g����Ӽ?��<��O<��r�Ҽ��=�=Y�<zp�<��F��k=Ӥ�<�"�a���6 =3���6���<��V��4q<�|�<�]=�͗;�DQ���;T=���k����<q�̼��/�W�B���%�ӻy�==�d�<3V�<)���B�<���<��=�=�/��]7�<,=�Mϼ�=e��gO.=�^=��H;2�ļ�9�m�,�`����E�	=>���h<r��;���;��
���߹�����κ�Qo=�]=���q�X=1*6���"���[�*{{= �M<-�E<֧��y�f<��*<,�E�xW�<K�<����/�<(���W��8d��{<2@=�2<� B=���I=u+�[�<��#=�(μV�d=�53���=8�U=��=�b��p*��={<(e<�z;=�*{�5��~�����<��f;���ɹc;y����c�s���W=�
&=W �d��<WU[�{���\��Ӹ�ZY�W:��h�;��==��0=vr�=�TE��E<@�ټ���;�+O=�P1����<�@����"<�)4����_=����<7h�<j	���<�ƕ�4|M�7��;�J=f��x ����J���<�
�<��z<nH��?�@�L��<�?����M=�!@�N=�!9����<�R;Z��;�K=YY<�L���G��<��B�����U\_=���ՕM;"�<YD��{5*;d�=��j��ޣw<�(��&q�!��gÇ�%a̻�>%;Iߙ���o:�Y���3�|�$���м�ZZ=����R+<4���o�S=M߮<1�T;�s�<�V＆u�= ��dO2=nK=�KƼ`9<�=[�������3uI=. �<���,�!=:`�)*�<��O<��e3!�1 =�F�<2-C=zm�)��;��;7P
��<MF=np�<��f��c�i҂<�I<^�<�~��NU�<��=�]=�J�j�<G`�*1Q=�i<հW=�|����M:�K��Gk�z4��\{�����3����bB<��<��/�`�����A�8�����.���׼;�#=������;�G2��=��;���̲c��=�Z�_K=`>"=���<W;bkӼ��5�E��<RR=�~�<e@=� C���<�}z��=+���_=����9����=�9�o5��mCC�S�<��0=:�=��h=���<�������<��F�޼��Լ C=�UC���"=���wP�<#-=�}t;���؅D��H�</!+<sb�<�E_<p@/<�VL=���V%ļ���D�h��r=�>=E�^=-��灼�80��*B���N<�e��G��@�8m6=*�A���=��<��=��e��Ӽ�F�C�c�4�$=)�.;��=���<I�:=L"��S��^O=]7���}q���o�X�4=�K@=�[,<��|��C�;��q��l��YX=����sV���G���<��<�=�ڼ�	�*C{=[�=㎇�ն�< =�hL:�b�������1��\C�10�޶<�Ϩ<6I<���m:2���UI=m�?=��+�1=�V�<9�N��}�<�s=��=��x� ���{H�D�	�JI�<��@�,��a=��<FT=8e�;�lo��;!�U=Ć@�.�b�ڣo��B}���;°Z�{e1=,���UY��P�;$a�<�*2=K :�Q 7�K����Ƽ��M���#=\`�<SWa�Hok���>=�P{�~f�<��N�V��<��=�C�� ={W+<v;=:�E�R&�=Jf=t��jU'=���Rg;�[I=h��U�$�.�~�1=u�����<J\�<I$=��G<�᳼�$.����<��輫�1=�a<=�/V����\��P�Z�_�;����n=��}���k��uW<��5���������D�m�<ZV;o�Q=�<��k=�E��Ȃ���_�<�C=f*=��;�a";�';]�"=��ɼL��<NY��P=H��<a�/��A�<��4�H��j;ZFw���T=�C=^�;={N1��D�<D>G={WZ���[=ό�EM=Jq�O��cI]=�"f=���O��,��<�%�9��<Q��<�Q�<��H=H>�ѫ������v�<�H���t=M�K�|t��]�=�/=�N*=�p��1<�.�<�����dB���==-��;��=�kҼ��������/�&A<�7[����<"'�<^�=��<�@F�-�K��Ӡ����9��0�>���=��2��B߼����/K&��<��O��=���<��[;]�0�==M�E<�Z,��i���4=�Q�<���4�;�k��K&�<S\-�Ej��m�����n�<�s=�Y=��<�=bu�<Y�;��=��Y= �j��
9�Ʀ<C|)=��)=NvS�
�4=ۻi��̖<W�<��zfW;Dt!=�� ��j<�0<�/s�uWݼ��{= Kr����i�Լ��<�0|<��<}��-�*�� =u���/�<m�^�h+{<��=�03���'=3 �����?�8��<	�i���;ny<_&<�����3�A�����<�H=�根-;�<,�}�4(���C����~��S������&=ݦE<�{=���;������<b�=�@(�V�7��<����բ��OL= ']��J���k<�.���?*�;�]�ϘM�SCg�UǞ��޼��3�<��B=��<�\W��L��&s=J�<�`=��4=VW��6q<�����Ѽ��<H�ۼӣ<f2/=m�1��䟼�E=�P����=��=t٥��:�<���սH<�����w<}��<�K�<|�<�r���Ѽ[���c^��ԗ�<��<r�a=tom�U~�< �;D���&<9Y=����,�;bs�<Wk=�k0��;=z�1�
��<��<+�G�5��<��Լd�&<A.�<�Ģ<=��<-�E=��=�#����G����#ֽ��ZP�S߀<w�<��<��<6�����Y�Y���^=F�x�W�S���g;��?��4�T�<��<��;Q����V�Є�<�?�m,=�?��Eȼ�ļ<
<����|:�A	�"�n�ҷ<��;��c=5U���ܼ��K=~L<�/�;D�
=��q��I�����PSk<��&�m"8�E�=�R^�5$=!$�<��j=p�<�<v��ͥ���Y���/��K^=1�H=������;:�{���<��d;��,="ż��û�����G=~ؼ�M��$��1J�=���<���<�U����<=��4��υ<
Al=@ߡ��~<�F�L1�<_�L=�t5<VȻ�<T$�<��l<��Q�A�M=��2���<B�<�D<��,��+W<N�f<��;Ұ@��V�g����;��M��:��� =���~�<G ��ӿ,=��Y����<G��;��;���<�!=%�p�i�	�N�:�o<��<�v���Z�=tP�;�W< B=S�<8Ou<��<����ܠ<�~��=ʮ�6=B<�����H=��;9��<z�B����<7=|�.=h�<U
��9ĉ��ZX��WS��`S�»>=��W��<�e<�bP=U$�<Q�%=D����<c�������a�= ��8<��L=��l=�2�2���NY��=0i*��w`=h:�Ԍ����/=�����b?��g�<2��I;==�8c=�BY�-�/<�+���r!;"�>��F�'/������*�@���=Hg)<jW�<����9������p�<�k/�EV�<����Nf)���'=.FX=Ŷ(<�7��謺�S�j|=�,=χ@=mu.�
$6���+��F=߇a="��<����[�;��=�]<']����'=�
=�~=�C%=�u�����<�~켴�#=dd��]A=��<��<u�;9R=�l<=�H�<T�{�;Xd�<���<̖=�<�)=|[�<3�\=dLe���7=I<�ͺ3H[��}j;��~=xa�T7[��=��=�f�n�D=��<��0=�5���'�&J=�7�<n=�^0��&�<�^�<4z��������T=s#=g:<��b���<�M"=~�-=�Dd��{S��q= 7=!�1=�D?=�G���<P�=2�=q�;�-�b��<����e,,�I�+<���=M��<3����(�t��<��U���;���C=%ּ�=��<t<{4��<��Q<� ,<{pl=B�i�<3=:�a=�4*<��R=���<��8=�¼��;���<�V��4�<�$5����:��F��\]�mW�<-�G=�9%=�5��N�G=4)"=�u
;�(Q=k����%<�L��M�<��N�/c==�?=r��<v��+����Z%<�:��Ua�l��<�5�<%]�<���;oC=��μ`tv<Hb ��i=b��;�\9��H<�x����ӆ��!,<����C�=�M=A.ݼU�/=q����9��<�u�<~Z=���(=��;�4_<Mǫ<��2�sf��+������;��3����\<�����<�i3<�p�<9=�^�����:D��<�/=��>��]��=���4]�<d�P=ȳ������@@i�IԻ�t�Z�=Ԑݼ[7=F:ּ;�==Y�=	�м�4R=�#����P�Y^'=�%ټ��=��ż�L=\<v���;J9��ټ�,}��=ּ'���A�8]��{�9g^=z;'<߻ͼ��;h�	<��Y��$�<5�.�}��<G�=Ӯ��O Z���0<��<O���b��<�@"�P�켤�?<t����:�<e�=�U+�<�~<�(=��n��g��5�<����D���\e�i��<"�I��� ���>�	�<�t��o><��"=q[<l&��ض<��h�u=h<�P�gV�W =Y���U�O=�Vh=&v4;~�{<��)�P=ks���Y2=�+�<��;����fő�5{X�M�=���<kZ�<٨=l[��@ؼx�F=2SF���$]Q<$���8�<J׼0��Oݷ����\��<3d��=�H)=�� �u�+��5W=�Z�7�n�hw���0l<�8<�
�;� �<��6�J(��_����<�?��
-�՗�<�O�'��<�¼�?�<�5����XV:էG�)��:�7q��@�����<a�<���@»�����<u�g=��=O�<�Ǽ|�/��<��N9�f������=��=o�6��I��[��<�/�O/� *<��G�=���9x,� ~�<�%���;��K��3V<x(�<�YK��<�@���Ǽ@�4�e�!�Ć�:6VD�1C���W���� =��P<ĺw=��Z<ͽ=�=��H=B���g<=��9���<=<X���=X�<Z�=���ʨ=ʽ�T��<u�.=�U��5Y�<F�{��wh<&��<b�g����;�9.=-�=b`�<k;�<p�S�<�ʼNd���=O��|�<�==.����*����f�s���s�;A�>��8`��=zѥ����;e>>�S���~<Ы=���>��;�V={����������`���Wq7=��y����|c�<��%�̻C=끂��b������fB�g2f=��N<q�S�M�b�O�8�����:sh~���X�9a�O	ۼ�p�����;�P==�.=��^��>��\yo�g�<ry����<Ӱ=�V�m9=o��6TA=E�>=����&A=R�#�N$����c��M=(#�}�=C�X��.�J9�\�G=��!1=�p%<�M꼴!f�v���g��~d]<�*=��P<xT���oȼA�R=��ϻ�Sb��=�Ĝ�]�a����<��7��@�;�=n����T�0G�<�߹<�;zg���==�+�<�F1<z�<�n�;�UO=1� �-�L���Ѽ�HQ=�Sj��l�q����Y��o=���<?*=�R4<\eH;i�e;S�3<��W�$vʼ�߸��p�A��@S��U�<��o�ݼ8��0��=oR~9�����D�?� ���%=���<˗<�#, ���<7F`<r�x<�̊���e9J�8ż��/=��0��P=�� =����˻�^�7=��f=����;W%L���ͼ���^c@�;Z
=�a*<7=�=��`��X��>=��f=�n=^�A����;Ｓ|��ɼ�W=i>a;��/=ڏ	����=�=������{'�!5H��绷�ԼZ���"3'�O�Ȼ��V�;�#@�z�=I�;�S=�}�<���vUQ���;N��:�g�Vv=��<d��u�\��v�<��,=�X��C=՗���V�<���R��<e�!=�稽�e�<N�=�v�o(�cp�b=!#��V�*%漜�0�4��<T
8�PI=ҟ5=���<�=�`�;��Q=�|��д��6z<�
��r��v��ұ?�OO{<kOR<(=k�u��j���`%�٭�<73R<�u�mvd��t*��.,<��<���<o^<!�<��
=�=��,=ZF���t��w'�@�,��v�΢*�tL�<�*���i;��i��S��W=<��<rʇ��=�����=�4�<Bu=�f<�!���P=��=f�ռ�5���:� =]R2=�2M�WJT�QT�;,MO����']�(K=�F)��~	=�	����<r��-�~E�<R�̼����x�;�S��
�R$�/� �E=)�	����=B=�J�;lv�g�i=)�T�p^f�cn=γ<����4W=�t0=��$��<e������߻<?�=m�=k_8=��@<�=������L4=D��=����%O�.3�<_�ڝ;��׼͐˼1�Y=�kR=ge�fY<����ا�<�2b�W�@=���<Q�K�ͯ��9���-S�����t=0�<?���� =X�@���O��dd<���<_h�;�oz�J�=T���];��%=�洺 ��<����#;/�uJ<=J�.��]u=�bU�
j �@�<���<G� =8�=Tc ����<��
��#��t<��=OO*=�c<��]<,�C==[l=������C=QP=�r�^�C<2Q.=+�L��B�]��<�*g��f"��>=���પ��ຼ:f�<���F槼P'=��<��S=�)<J���4�<��<�!g��=[=����n<���<�M���޺-�̼Ѕ�<�=�r;O
��G�<�TX�Y$=�ݥ<Ic+=��=xP���rW<�e�<'�켊i�<L&��9�¼���B�*=��1�|�,=0��;l{<]��<&8�<@Sμ@�1��7j=��ɼ�G��J�<Am�̘=��=�Z=�PU�&I=��"@�kU'=w�;��<�t���:<��ټS�ټ����apb�u
�\��}E=���P�;7��QA���5=.>�<=��<��H=P8&��5��Js=�=��8�(���cr��?����<j��=gT�<V�����<���%*;�=9� <Wy<��.=�ms�yV=�¼�Tc�l��<��w�',���(�;X#���R�W̄���1=������Ogb�T�;�[��~4=ہn� �B��`{�	��<�e=�:�=��8=!��NWW='q=@�I�+�=��!=�|'�IK_=��S�J���1�O�k��u�<�V��
��y�:䅢��G%��y��uv<�ʐ�4ʱ�}�?=:��;PO�<Ӽ�[�<�_�;2W*=�6�� =����� =(H��2�o=��I���];~ib=]����f$%=A��(��@���p�<0�7��2��;�Y=w�3="��<;S�<  6;S�n=\Ǽ��<��;��J=�8��'L��{0='�;�b/=F�;/!�<��-=��D=j�6���?���伸��<a�F=��`�Uo����<n���߼H��<�\<#�+<}��<��9�^�<�Rؼw�5�r+�;����(��|�<z��;T~=�`׼�I=		�<�;-�Y�<���:EY�s���.���`�������d{=.�P;�� ��JS��_ �zZ�<Z;A� =��*�3�w�����D�������<'X��&���`��_��|1�:F���\<�Y��=�qlj;A�i<�<�FC�����=�x޼o$��U��C�<���l�<~:=��a��p��ak	��H=?Q�<-�=���9Լ�<BU����B��O=�y���t�<�=[ =�\�k}<��=ǧ�(�?�C!=Ą= ��<M�J��i0=F�7=X՚�<���9<8<=>Q/<��5=s�5=���<�ɀ=�f����<T�E��7=B��=��K���X=gK<[�;��<�[R=5㞼	*���߼��-�o�p��EԼ�y���S=�9�ѻm���ih"�LE��kb��oĨ;W���Q�rq�or��8$'�>ݼ=�n=L,�L8˻ɿ��}O��Q����BӼ^j-={�=�b!�<����l��f�����;���<
 �S�����B���<z��<I�<���<b��;�i
==���=eH<�vk=
 �Ծ<^O|<:�\���ߧ�w�"��E�y�G��vb=	�B��U9=_L=�Ǣ�ѤX=�2�������$=�h5=�QE=�ر<�����f���=#32=x�i���9�_���#=���G�=�5����<��L=_���"<=�ͼ<t	B=�6=-��<�<vJ*=��:�d�'�9ĉ�;��l=�d�9��;_`!;��_�;5H��ü��<�ꅺA{5=�4= )�8k�H�j�=]�<P����:�T,���+�E�gG=���<w\=�<�w
�Y���z=��)=�Q��`.�ϑܼ��<I�2�S�<q*ݼW������;;p��=t-P�ą�<��{=� �ʩP=Qg9=WO{�˭=�� �q7����<?U�<J-=���<��༼�<ذ~=�e0="�����Q)<�WX��I =�)h<^Y�:^k=�#�<	y��^?��m�;L4�;�+=��q<�;^�'���j�D�����a=��a<���<��%�v�+�����Q=m0|<xW��f�< �5=x50=G�<�#����U��T�<�E�;/,ҼW��έƼ�uƼo�4�zI�<��:��/�<x4�9x?:��̻\_�
P@=���<�8�<���;�Oh=Jַ���~�$��<*iL=���� �;`}=�î�4Y�<���<hY=��r.M�&�i�]����
N=�u��/%�}0�s�*������(�]�h=l�;=P�U;�?��6�x�<=������<�Y0=r�<��H=�c==�R;�J<�&=:�<�
K�W��V�x<?�w��l~��A=��E�2��<��1���<{D���I=����t=��ͼ��<9��Fޙ<o=D�H=tV����r<BX�K�*=���<q�\=ڏ^<w1��+;,���߼겗<��=���9y[=�!�٘9������B<�y��:(�u�\q.��OK���e�G�	=��I���.=Z�����<g氻)�==k4n��LH=��5�=WU��Q�A��;Ŋ����<�轼����9=�K	=���;}���:�'=��߼��
����7jS=������_=�u/;�f��]��<r�}��1��TV<�N=��=|�K=�Q�<�=e�N=�_$=緉�ޜ�;�7^=�=uz\�5�{�g&!�.L�<�f��."���ǻK�:{�<t�<n��<l�<<􎪺�׼Ŧ<=��9=�Us��$�<�=�
��E���h� �!�A=�� �<&�	=��=Y��+;L�O=��x��j;�ܼ�W#=�ђ<<݉���9<�.D�=��;Y��W�v�4�I��?=�-�����`�;?�=���<��d�#hT����<��/�y�*�.��JI������D��d��*�<ڂǼ���<�}O�ǔ:��N`=��:i�&;��=�
��̽E��`�<+7�;a�ռ_�="�����/=�-��h=��g���j�/=�m��}ļ����ȑE=�䥼�H������-�Ѽ��м9�4�LX��^�9�ἀg=r�9�n�u��<~3ڼp��<z<��мx��<k;=�N��v�<I�k���.��_]=�"����<Y5��hQ�9�AN=c��;`�"=ct�;��=Y�w���\=́<��޼<�z<�5�$=�&<@��W'=rm�<� ��@�G=�\=��;<>�6=CZ'<�����ͼ�9��Oؼ�r�
�eF�،Ƽ��m<4�����L��<�� ���<�i��k-���F�2g¼��=2�~<v�<=�=�<��
=t�= ��<��t���>=E ���K�/��5�<��{�P)��}����<��G<)�<�2=K^�<Tؼ5�S<������8��5��
����<Uv`��T#����;�g&����;�A~��8X=5K������M伡���=����F�<����.=���<\���&����<E�<��;�8=�Y=ߙM�[B=h�w��μt���oZ�D�!=*�ؼZ~�;�`H<=�:�@�<��<]���u�.<��=�ע;�{�)�<��<H��<S�!���ٓ=��R{0=��<�uy�����{�!�2=4g���<*/��PZ=�Jn����\��<�J=���<�CB<�7F=k�����<�=�u�h	=�����%=�w	=$)ܼ3g5��P˻�AP<��<���<��=?)�<���7':�HD]��� <"<R�:_6=)f;�.W=�:+��Ҋ�	8-=ډ%=�J�UJ=^�;����BQ=W��Dʼ�H=��:=�Ld�"��;C�R�-g���]�V�}�#	�<��<B2=��=�:<�HG='�����<�<�K�<f���R<W(�<�h4=��:��S���üj�;l���ӆ��T�<+��<"��<�=ҡ�,���>�3��v=8�.=�S'�>��LL���=�3<6����N�<5�b<ӥѼ���$�=e�=�?=��8=���<|���˼n�	=�;��L�<�=y�<@��<0�;^aJ�����(BE=sYx����������6�ph�<�%�D{k���<i��<O�'��=����<�Gn<���%���<���GJ��o�K =�GM<�Vr=`�9<*=�D��x�=0�H�s�<��<���:��1)<ɮ�;�DY<������,��=�Ϡ���;�z8�߈�<�i=#���)�=iX<@r� �=���l?d<��ڻWb
=��<�=�t�<�1c<����$�=E=:��M1=7'�T�/����;��g=�SY<����$��=�l+=�I�;���vﲼ�Y/<��<=-�&81� e���(ռz�V�BZ?<CE=!��i<Ds���<��P�l��%���,�.����R���V��ӏO���=kS�<����i=�<��ϼb;P�ԎY=���-���x<�����Q=��=Z3D=��B<]�;IW�<���<Ub�;YTZ=?�����<������:뗷��=� �<4-�<�I=�[�e�`<��{���?=�=�b�<R�i��T����<v&]�rJ�&���N=z; ���$�	?��ފ =iF�<��=��;��)<�[�)/�;n�3=l�����U����i>�{Ɣ;DC�:��y�݀T=��x<���<�	<�a�<2b��ߔ�o�<�^P�B�=��5�5-�s�P<�ޔ<s�=��<u��<�ۼ]�̺A?R���{=��<��=:�`=����0���P:=��;<��`�ǌɼ�㐼�fU:#�<{�=�d�:�9�����<�^k="�-<$=��;1Wa�z�<z	<���>��2���&=\�4�xм?�$�5���.z����=�r=��#�L<H!J<̓��S���9��&�<29*���3�����=茘<jU/=	bl�~e=�8=9[#=&��<��I�6&�0�Y��R��Q7=�?7��,Q��^ü�{y�=�!�/�D��Z�=��$��u��=���<|�ݼ�44=R�8=���ҳ�=:$��vk�)����'v=9͕�Y<Lɹ<e�>=7vh=�#�����q.������6$=�:�JKr:w�!<D'���b=}O=_nj�D��<oO=l[⼩��<�O;l�*=�,��zj��{B��z޻PB���<���m�<��<�����#���h�����q�<���;� �;O1ϼYO#=j�dA3�ӉO<��p=7��<�U<=qj;�0μ����� <M	G<��J�h�ڹc7��?;=
��< 8�<y� ;z�!=�Y�<�	=	+�Iy=�M�=�L�(B���#<�cg<����:��/�<��;�F(����jp���F�<������r|<`����;M�J=p=Ji%;��n�V�B=�f5=����Y�:�h��0�<�an��w=z^;��[�<.�+�W��;e/^=��ּ9�E=�l����M=Q�=e�<?L,��W��1ͼi'g�Yh4=���<�U+�`��c3�<��d����<F�<����%�<J<H��O�]@ܺ6��L��u��*�n�^�`��M��b"�[&_������=�߇<0�p����<H��<K����)f=�e?=��b��D˼���<OQ����o�}証����Pa=�A�:Ӧ���G_�h�(�9�/=�^��+�-�(��o�<@�
��u�D��<$���PE=`�=K��e����� (+��������<��<��8�0X �*���׼��S=��"=V��<b'<7=�+u�:�Oy<��D=Y� �={=��e��Q���ݞ���=5�A=?�6=j�j��?�����$��<��"��T�<�W=�LK���O��Ƽfb9���O�1��}�=�kl¼�/�<��h��==�2��"Ζ<�TF�&|�<�Z�H�����9��,=���L��;��+�
~V=��'�A���	K���7����� =�
�=EE.=K+�̢<���<�苽��<�)#�O���押_ɼ�z���-i=���<[z�����=H�=�h�r�4��zq��!\=��<=�ߊ�G*Z���;��<-�<a&=Nxj=N��:'
=�儼��q� E����g����B�;��~�W�&�}���6=��_=~T��`�{A�;��<�l��K���'�ʗ[�M@�~��m��<v�=�I꼄�X�z,�����<�l+=V�D=�;�=<�D<����{~N���<w9=�b��Ʃ�n1�<��<AQ�<��\��V�P<���5� =Ƣ;=�!�=�K}<C(=�[=<��I;R����<�"�+�����s�z=$�A�P-��U�2�4�9=F���}1!�m1�<)Q=&=Z;���H=aa�;]e�M�<IMp��%�;��� Il�k��<��<��<^N�uv0;&�߼Uc=w�6=f�Q�?�w������Y�_e�<��v=�Pl����<�.�i�=��8����8�!�<ht[��W��<��<#�ʼ�`<U� �$=�!����;��:=#�;�k�<d18=��	=�rd<��#;j��<Ň[;s�=l�<�E�<�a�t�R=Z��<��;=�ؼ"�Y�p=Q�μ7I<�B=A��<xH���d<8�=~�T=FO��W��Q=�?7�I^V=%'���I=�b%��'��"�<ݛ����f=;�#���;�@��$��<���<d-X�4N�;�A��-�<��<u'���/�i�<��W�u�j=��2�6��<7Uۼf��<O�=#�<`.�<g;d=[I�[\:=��<
d#=)�Ѽ�ϵ<o�,���;��d =ڷI�-=�$ȼ"��<3nZ=��/=X��Mo9=��=���<���<�jG<s��:�S='�>�azl=��^�t傽৙��S��4����=�J?.�%��0�<�&��Q>;�沼!c�9J>���]<�p�|�X�f�<�e7=��<gj��޺x�<�~"�� #���1<�MR�g_	��!�Z}���<���`6";qN�l�7�袾�0�T��c޼Iݣ<�[<����ĻlW=#�Q=�=�G�=��M=F�Ҽ�fC=X�E���c=Q,���y#�T�:��<��-���v���6�7�t�{?��������P3=���=g�!=5�U��)Q=�5���mּ�N=7H>��vw�S�<�<:3r=�ʍ���q<��+�]��5�9=1=t¤<PJ������C��f>����<�S	=��;;��k� o$�r���%��*�1Y�<U-q=Qn/��_5=	.j�o�<f�;|�H=��g=�&�<>E�<((=K���z��B�$��;V��<��cG3�HO=�����=\=Z+�Z�ռ�v%�L>=�[0�LZ=k�2=�".;���<�ļ��E�4-��B�Z�N���<~�F�U�=�+=�Nv��Y=Q	�<Ƕ�<�$=��׼A+%=H��/��x�]����Ҽ;���m��Rd=�O9�9��
�d<HLC=�v�!�<��=�p�(=�I��t�v=0%H�/ۼ���,�k={�P��[�����<��G�fb4=��5��;=�K��(P=f�A=��s�����v���߻�B=P\<�= 
���g=��g��,�=�(k��އ��l=�zX�"�~�UJ�<��ػ�!=8<
9���5<=,=T鹼'q�m�4�]�:�g�<F�=��r=�:@=؛�:XI�<V��'��]�<�I�(��d1���=瀑<�Ӈ<8xW�&W�;�\��f%=�T��{@���X=��|=�4!=��<r��=�Z�<����=�<���/��9IU<=0����<|[U�8^��jHY=�6=���<+�켳yX=1�H;��q��׼}|+�W�g�p����O6=q=C��0Ex�����ݪ=ǃ�=o��%�<;��f<Q��<V|=-�.��=��&=*�{��b_�"�n���<#�$=@����=�R��|c��-"=��=<��W=z�=u�@=�zn���n̯��S\��T�<J~�<�"s=��ɼ�e0<��*������O�y�~;�;8"��ظļ
���~����<�����/����<����P�<�:�<�a:��5=v��;bV&=X�V��I�{)V=��n=G:�a��<C��:�.�!�	=�[:���<݉A=�8�~ۺKdN=�b<�Jy�d�<�V�����-X���-��۴(=H��� �f�A�vO���>=��?��G1=��O��IM=%<&����q=� `=�|V=�D9=zP<r`1��Po<�A+�s��;Ef�<ȧ6�
�T����;8;)�i�����;��`�F��5���g=&���;���;FѼ����0`�n�=��<��<��;~���i<�Ї<�vм�[��4ZY=��$=u3��?�O�U+=�eg����T��<���<=��몼=�=h�<1�t�DQ"=�=���!�jݽ���N=��=C<^�9FN����<���<��Y�l�C�b;L����<�l�mb�<g���� �F�����=Y�<�7!�/�<���<I/ȼI�A=��4<�p�;�k�;��X=�#y��&
=fj=���4�=�j=L_�<X9=���;Q;�Y_���<mz<=��[�Gp�=!}I�Zr�<	�<�=�Tz��q�<j=��z���
=3�h�u=�D�
�Y���D=&�'d=�oe���2=��;<X7��
���U�o�Z����<֚B=�1�<�)=c�}vF�=|`�̀i=�O�kL)=bg=�8�"X��K�<�'=��g���A;�R`��~�<�=�;�ݼPm��&��kۮ<SI���U'�'ݗ<�V=a�<-�d=�e�<�n�<�y="=m�|��e,=��s�K"������â�<xby��{=�]=)n�yd=���uc���==R_%<^�������3>`�?�x�P�9�@ʯ;��<E��Z���=3S=3��FYk��"�����<�4�;��r=��]=q%<�P���PU<��/=��R�)P%<��ҼjE=�p+=�&������*=����A<ʦ)��#=�?y��q<��:W󜼒Gm��wN=��<�}{=~�~=S�=\�=�z�;ñ�G7�$E��Hf�".�9�<1Vr��N<rQ=q@u=��ʺ�f�<�	V=�*���q��E�</C�"�����<1��<_%L��	.� n�<ų:�����Dj��	=��<l�C=r/�:Q�X�:�"�;m;:�=#�]=%�ͼj`	��'��t)�qK!�ɿ<���<���{���~==�=Q��:e��<�+�M#=2�=�o(�Q<��=3�7�\����9?<�;�f�<��j�vK=$�&���F��%�zs���B=/r��H;D����<#a-=C���>�F!X��G�W���!�M=��U�M�<�=�A��쬼ڥZ=��y��C�����6�z�S<6J���D�$=?&��E�;	"��hF��`��eO��ڣ< �M�x�<*����5��<�2=�P¼I<�<	r�;teb;?˹��6}=Z�+������<�O�!��ձ<I�D=�a.�ڂ�;�i��k����;�Y=M�<9��)�p��s<�PG��6<���+��;)��<쬣���:��X���\���<ߏ�MH<�����a�&%W�
��<������=��=�Y=�w�ý)=��$=�?N�_j��u�T=����i�<�d����8] =n��<�q�r�7=|[<�$=�L�;�'=���<V=����_*�N��G�3�TR��
�<@=e��벉:_����'�<ߦM=�Ҩ<M�7�gJ=��S��\��м�
���>=��<�X��'=Ƕ;��[�r�H�m,<�*�<��$�N&ǼF9W���-�\�d<�6�p�1����~ݼeڔ:�6�<���~hf=��q=/2=���<�܌��}��}���=���d =������߼�`��v��� ;��d�8�l���JM廄^<C'=#�$<��<rs�([����<@��;�ü���<���<P�=�)M=[}X�����=;��!=�<�3޼��P����!�����>=c�f=m����(�䳃<�Qp������(�z�C=y4�N�/�p��<x(@�-A5=U!!=^8��,�;��<��=�Մ=�L��6��<FN;�!&�T <�T<l���._�k�<�U�������!���H�onk=�=EG@�k%�;,�7�ɫ�uuo�(ǀ=%c�:e<��	l\��c�<�]���[ <���<���<���;��<i�5�y�;<3�%�=)��<��$=��z<
`�H�<T		<Q�=Ȧ���ɭ�ʥ<��
<ݦ=�Ha=4ԏ=�N�YPi=j1�<&g=wn1=Xy'�¦�:��0=�O:ɼ�\;���<�0ܼ\�<z#<��$���y��Z~<��Ǽ��<�g��ޛG�'M��}��-="#�<1I�<��O��|�Ы��orQ�{�%�q�h=��r�������<)����A<=-Z�e|I��"^�(@���(���2��=���3x=;��'�}�<�-?=���$��b�<�f=�����N<l��,<ƻ"�i�����RC\<�O5��!��5�5����2�<�u�<�A'=�<�������D�m���;Y����X����1=�J7�E"=��j�C�b�.ę<���< ��;�K��Z�U�ar��?1�$ߐ<��9��<=������f��P���/��<Udj�)���T�</㙼^�B�gom���<&��n����;=R��D�l;�<��J=��Ƽt-%=��<oT=DB=���I=I]!��5�;��
��5y=wz5=m[�<m큼YN�;r�
=��<Q��<��i<f�>=+7\��ao=��,�e=\#�:���<:�J<^m
=�DӻK<b��E��
���8<���)ۻ�].=F'��qS=� 1=�_���_#=�o=8UǼ�<!��:�Ő=�B#�,����/=o��<�l�<�����s=4}���O=�fz��o��U5��}��b�<<L��=w2�*�@=2�O���!=g\�U=pC~<ʵ`=	�x���*:-	)���=�-��)��'�aP=������<��;�T^������m=kL���n;�ha=�.t;��3U==���N6d��Ҽ�cT<����]�;_�Q���;�n�y=
�ȼZ�<�==m���r�g8x�%<���<98m�$��9�<��2=F�=H���Y>3��VU�s�2�t��8=L������~�<E>[�w��<I8b��`���˼Q[���g<L�h=�ĺ���<;��%
���@���w=ݙ�P�(=]㩼?�<�u<R�Q���*�^<�a��I��Y�<.H'=� �Yf3���<3��<x�͓��h�<ϑ<��=��"�g-�;/-޻¢<=:ý<:T�<��:���^=��]<��]=8�P�O͑<5�=���=tx�PM�<���<^�/�B=G>��ތ���Z=�1����$�§*=�XG��j<��<��s��MT=�gJ=~{�9r����6����<�/ϼl�%=�=@�a�b�У�<���B����H�Ԗ=����]�ռ��ػ��s�0E�<��;3=Mo�0;[<��<_X= X5=W%��ut=�;�<>^,=x�,�~b=��>��":]��<�<�<�Y^=�Y��K���	<�Aļ�@<Q�B�9�=Ȱ�;��g97�=�=�~��I�üm�5=m .<FļPc<��=��I=Vfo=�j�=tZ ��%<&�E=S"ؼ�灼6^�<g�;��y<ԑK=�1<���3�<`�Ҽ�=��ü����@�39H��<2���6�<�/�<)l=^X��H���<k��<B,<�z�S�<௅=�Q=��=֦�X�o=��<r��;���<N�F=�/����뤂<���<q�#=��<�Xw<����T�/;���;�ݎ<[�Y=�3=
Q�~(=�D=_�A�9�d�$�����V�/d�;�,��T9���<#�=h��Ib�;��_�L,�E�\=P�����=�o�+�7<��<����#�,���a���
��I�<2��,cN=2q�:�A=׮�<E#=�����7��<R�t�V�=�/4=M�;l���sx㼯G���f=Z�ʼ��Լt(�7i<C�3<sIW��퉼�u����<x&ؼd��<�/Z�cS�<���<�eݻ��'=��_��:="K�9������ߺ�k���n���<���Լ���<):>�O-^�z�]=?��c౼@3�R#h��A6=WF>=�~���.�P�~��l<<ұd=E>������ͼW�!=�#T�fVd=��<V`��	��<�P�B���=�G2�>k��$��̹�4
=�j=M�1=���<���<2�\=ۇ
=��ջBP
��o��P��q��	�e=�g{=�ip=�j,=�#!�[E=���;]pB<1<C�Z��0��C=%��<��9��D��^��������X�8#�v�ϼmf=��k���U��<�;)��PS��A+�DV�<%�<��Gxs�|�	���K�����|$s�wi��d���^5=�"f��xG=��*���|}N��
=8"=����=��D=	=,�+��2;�����
��+�!=s�'�Ҁ<�\A��h!�^G=�:;&�\����O=�I��<��f�;�2=�>!=G=�^:���<���<I'�Bc=o���2=]�A:	ꪼ#� �9�6����<�I���%�o6/=ؑ����=<K�=G_"��U��K�S<�/=�tA=Rf�<>�n��<���;��k��<����1�T�Ȩ<�&,=Z�=�]���Y<
e�<�Z'=	@==�f��<@JS�������;J�ڷ��:=��6<r"�	!<������wQ=� O�Zk��v���>F;���<90���=C=N?�&V���嚼n`�J�'�^��X�W���d=���/���=�
=z!�<�nh=��u��U�<�<�����ӖZ=���w[=7@W�6/(=J�`=�m=FfE=J]=/t�������>=&.P=h�\=�P�����2<1�P=e �AET=m��<��]=1 ���Z�����<?;�j漓�b=�����f�a����=g�Q�T���"��<��
������z�J�ү���:�=CF�tE�<G�Y�Lty��Ү;�~˼��8�e�=x�,=�91�Vԩ<\�Ｑ�Q=��=He+=k��iD�ݦ�<�������:y�C=�`=�NA���w<=��I<�u���=�ټWH0�����Yr��=	=��<͹㼚��<_�=)X�<U|��ض�����;\�s�QA=o�޼�bi�hQ=�'�?ż�K=V��J���<�j�~=�������;i�; c��Ӑؼ'�;�A�<fN�=��&�<�Bx=���<�n#<Ǽ�+�����7Mp=��<²r=�P���.ʼ��e=d���E<R�=�'�{�<��=�f�<r��q^=��=�O?=@=*5�<@��< l=E�0����S���I�<))=ij�<,$�V�=A�5���S=������<���G�t=ED=�l�9��[?j�� <8�˼�yi�� �I��Z���o��b�P�*3�j���=��;���<�K==�oZ=�u#=q��<�Q��<e�	=��:&=�E����<o!=z�=�L̻�s�<'�̻�+�&X=�ҙ�Ki="�9<ԒR��T�����ص<'-&=6(���Fz���-��<����Q��;��;��μ��<�����+<�f�<�R�;�7h�
�ڼ�v��3��)L�&h!<D����T��ћ<���*8��<A���:��<c,�<��<b�=\	G���]����<)�/��U=�<�T��7�@�ڮ��El���Z;ُo��.���]=� ����7=�.��k�<�Gm;84"���=��:���<��`=Ʀ ��c=/�,��<��O��9B�@v{�Sa���(>=��m<P>�E嫼'd=��;�P߼>u�N�3=�d���d7�¨P��˘�kF=�6�0�ڼ�<T<�=����,�4����<���<-46�	Ja�h�;��d=��]iǼ:����;<�IM�w]R��u?���������;�f�<T$;vt=Q�i=�O���������p��,<�Dk=*Sg=v�;��p��K\;qG�<�T=*F"=.都�&9=�<T=7<��ӻ�'ɻe����}�<�������|4=�x��<B���H�<�A`���{<V�<�:>��%=<Nۼ���58m<�w,=��n<o4\<�!�=�
Ǽ�$<w2=�����\�;F��<�>!=�J�<�f=غd�d�;L��� =-g׼��B���-	=�3��ޘ	�H =��i��5��+=�!=I��<��=pO[�1�缧ة<��!���\�<:�<�w*=�������Y�7 w=p<<D�O=�{=*)$<X���E-�/;
=���<�T<��j�}�:ۗ.<�x;#A��[pQ=K��7@<�c1=� $��{Y=�?�<(�=<���<��1���=�m�K�]O<�_��y��<��N=�,*=��:=�2�r̻i�C�ˏ��mzy=�h:;<�S�E,ݼ��|<� �C�<]��<�I=$Q=�%�ßF=b.E=:�	�ヺ�}�;:�����I���<���Ce^=�������<N��<ǿ�<���<�$�<uoL�eeJ<-ĺ��|<�K8�Q2��/(��A�<�;���C=74<���<I�Ҽ�)�<��=j�μ%��<� ��"c�������X�@m.=�
=�$=1R	�3=�ǒ<j��yr=%YT=��k�����/<7�9���!<��:8�'=�˼hG��Ő�!b<c8N=�N��R=Y
�%eb��N�<��<�;E��*����D=�1U���4��\���a�<�}<�[=�Ap��e�-�`���J�[�c=� �k���{�����? =Hm��}	=m�<o���G�7�N��pc:�.I��fӼ?=�Z�Ű�<�`B�]�R�r�<�W/= �<�I�<���<ә]=g2<y�.=7k-=
=�l�<���;d��;S�j���S���R���|�6[:����>�����;NRH�٥����<�ZU��Q;F[�<ls���`;VI�	U�'rS�T?G<�-e��r=�=�L�;��#� ��<�V��M=t|	�7ռ���<	���<F�Z�M��=Վ*�׍�{1I���;<ɮ[���=�#=��+=�^���9�'��!a[��`=�$��k�:=&�p=O�� '�<��$=��<�򢼝7s=��D�*x�:N[3:��<a�=�!����==	h=�1k�{A+�SYӼ�ka=�C{�{�~�.Ƒ�1���=��<�TZ�L5E�օ��b`=�Jl=�='=*��%<����a"��B���O"=(�v�
�ݺl|N=%�μ�R/=�{�?
�;�=)=��<6�'=S����/=4Đ��==7^;)L�aU��R��=��?��L�������<�>:=rmZ=Я[���M���;\.��e
o<�=�{�}�p=�����<d�
���i=�F�>�m<쮽�ʑ�����<%���'>���9�)H�M��:����-{@<�`�<��=
�t��h�<}�<6�Z�6�#=����s=����¨0=�5�*������F�̛P=��9�7�=�ü��U=1k�6O��j�<*nn=\e���<�J����ؼ$��;����{�;o����;�<%����<�d�<D 
����<(�k�@���h�p�p �<ăJ=�<Q	�<6��<yr��&�c=V�u�.=����M���䜅<��B<	P=���dK�h�E�����L�q$X����A�D�9�V��6h;�R�<��=I�+=���<��<N����<=OQz��d=۫��'ۼ=)U=�2��u���T=Z�<=il=��Ӽ��⼉S =B�`=̣A=V�=�5�/T���e$�V�c�=��<YZ<{=O"�;�0��]R���<���0�?��<B�=�T�h��n�;��"��=f�Eҫ<��/ ��7�<�1��)�yp=w)|�(�����;�'�=_`ʼ:�����k�8�û��!��^�������*<�������7<����pƹ'��<��S=��F�aӜ<�=�U[��=9��N=,���(%��70���O��)=���<Іp�q�(���8�檰<��G��쀼J<�;��PF<ـ̼oO�<�E��0�=�Cc��;<�%=.0��d;jg�u��:�'�,�=>*��`���t�<P=j`��nl=��"��"���<��J=j�ռ&z��N� E&���4;gJ��$�=�_<�-�<W��<(�ּIn=�g�9�=e=�[=ᓃ;S�����뤇=U�]���T�}�=8"�6���ȼ��<8��Ot���?=�r=�=|���5������P�<�x`=�]�S�d=g=�L�<���t���|���K����;���<�|��OK=�g<���R�=�w�rC�b.A��)=�}\����<�2#�1�W�8Ƃ�г�mA=�F<�?=P�;�ܻ�O<}6d=��Ҽ��E���3=�͂=��X�8(]��z�=�-�,@�Ge��s+�,�(=�K��f��a�Ҽ*n=S>��@=��k�MG����U;�}<,"��Ν���ɼ�I�*6���:�o�C�*F�<�,��Ѽ�C=��<J��μL��<�<����`�Z7^=��
=ַ>=�~�<jE���j����+�����j=�������G"���=^�=u,Z=����l4��� q�,W�6V炼�L�<*[�<QPl�X[a:�
���c���K=��]<2g����<��=�� <.�<ɛ��r=���2�%�<N =��B��)�|G?�������-=�1�<����&�<1�R=��2��X=?����k�<�/׼��_;3�a=�5=�@)<�=�4=FS`�V�><�����=_p�<{"m<�}m;��W=��B<OS����<�
��:�u�<��`��h�;`m:�һ��=�=��D=��<Q�j=����kJ�(������ll9=c����Y:=�e=Oj<^����.�|E��b������<�[=��?��|)��]z�����j��[<�5&�����Z�<|I��T�=�����{��xTϻ��������%�;Q���a =��<�(�� �8l!=.��i⸼KB����<�.8=T�,���#<<b9�T��!>w�F�P=�3'����=;�J<�]e���<֥�!=BOe=C�;=z3;<��V���=���%=��7�"2h�Ye�<��=�K=L�j,�1�(��2u:51=��ż��<^~�<���� ���w=/�<"�={�D<l�����b:=v��<����]m<��B=Յ�<�{	:��=n�X�7ю�f�����|:����'=�8�<o�ѻ�Ax<Pۡ�/�9��@�<�(;+9=!�A�B=p?�G���d㍼�/�:y= �t����<'`j�-=/^=-�E��&^�C�=�ޅ�ܼ���;����Jx<;�����5=5=�o���ӻ��A�qLq<m0�<VC=���'���=��<�J=���<dR�;3(7���ּ�!_�6�c��rV���мue;�E�<������M���2=�:#<p���B=F�ز߼�=�5�="k �v`�<�j0�T[�<�C��E�<Q�~�(�~R8�m�<7l �D6*=���SR�=H��l���<�	=�j<7��<C�<s�?=��<+r�I�I�aN&=�i˼�}�	~�<�^=�ӥ�i�<T96�>9���=�R,�8��<��=�Z"=� +=���p=��t=��&<+�����2=�W��x��3�;�mb=�,
<�0+����;�����S �+b=���k8$�M�
=�v�;�k���m<[�4�1*=�Y��J��:򺃝Q=0�D=)�>��ʳ����:@Tf�>��1B���t9lb=+_�;�4,��
��)=�cS=����+=55;_n=��<��+=��;b;�<pD�<�X��9�z�[<��U=eM<J	ֻ�������=��-	!�cS���u+�=��j�+Z��2�<׳0=��R��x��ר<�2=�(N��t�?-<���<J$���
�l3�8��<��r=M���i�;,��%=�x�gx���s��^=C6��/�S=��^;Jy�<P�?����<���#P6<i�W�=�;�Y&;�7-=�2�xx4=&�<H��G��0=c�ռR=�Qѻ�%ټ��1�v0����w�ov(�����9��};W�S=����`!n�h�2�"�u=Q9]��mM<�~��忼�{�g�<7������,G=  (���G�&f@=�W=�84=]$��v�t;����D{���B�/Y��W�<��;Ds=�S=��<st�<�{7�KY߼>�<u�;���<�Ǫ<�5%<�^�;��+r=�)��J(=��<��'���1���	Nļ�B�<б=���>p&=������<���<�h=}c��! �=Y�������WW=㱼�u<�^�@=Eⲻ��u���d<�@=^�ȼ\=�&L:9\�����Z;�T�&/1���?a�n嶼�,q=����*{ʻ��<�72=�΃=�S�!�=z� ���3���Ȼ��;�(4<���\(=��7�V��l<d
��+J=&���.�5R<��i��<���:?=�h�<�m�<�*���M(=[�`�*�-=�q�+B���3�j�j��ݢ<{�b����<B��U�E��-e�b (<j��<���;l�ۼ�P/=T�ҺLj<��<��<?�c��U=+��<�K� <�-=M:o=,��b�O=�U�<a�=����m���/0=�^;�Z����<�Ҡ�w�p��0�0=z��� ��;��<&�?�e���P<��Y���;�#=�C�ue��v�;2{#�	
��E?��;}��j_=~��I']<<uN=��i�wj[=<"�� ��1K=�c�S���\N��4���+B��kѻ��<e�<w}:�m�<�r���<0;�˄=倓���=����q���<輛E=���<]���a���
��=}]�<�� =�k�<�d'�oQ��$ĕ��b=��D��9M=ܺO<�1�R7=�sǼ/g�ló����<���<�B<��#:��o�h�
��6�<�����<��h���<MYO<�T�"V8=�.�<c��;�L�/+���(�Q�l���<D`=yU�$B�}G��c�%<�&f<x�<�>=��z<���X�H��㕼xÎ<�|F���ۻ:<�<��=]D\�y.���ۼ"�5���G=F3o=ڽS;�Һ<�}�<�qa=Y���Ѽ4�G�#X���7��H���O(<��~=����<K��;��\=h�2==��:LQ=�O2��?=3''<�g���j��,��<��=�˼�2(=Z�8��,�<�iüxu2�#��<���;��#�&�<����蒼
/�<\��<+�4����7�I=�@����<�ڸ�IlV<��=��-���o��=��=�M⽼8bm=4k�;W?	�ʭ`<D��<��$=�Q�i��<�T�<�[�=�ļtH=/�<=$�#��=s�=�RJ�JLX<�X��!��G��'��բ;��=�/�/�J��MO�.�<�] ���~���8�R�Y*�&��DF�;n��D�;ǚӼ���͗��U.�����<h���6=t��;rD=R�\��*��Z���<���'�Q���<�蠼�Vy���\��8=��@<��R=���=��;�Uc��ۊ��T�;��.=Fw{�D�,����X3d=5��:<�`���T�=�$�; |K9�< P=�h=��<�������)C�<�K=���;�\=�a��\R<�_=��=�=&<unB���N�Y�;�5=|ż{�"�k <�Z�<��3<^$:����:x���P���Ѽ�|[=�5<h&ິ��y���Q��b�׼���;e�E��X�>����<8���T�H�.���#<cb=�/C�emD=��w�J4��%��;�h=:#�roJ��N=j�b=�#=�/,��=��:=�ݼ�W���=��3��tK=��e�5y�<����� =�=lYq=d���;4B�;�f�7�L=ׂ=���l���<b@G��V���%�ϯ�<8C�ڿ	=���;�y��K<��:��(�r�d�Rܼ�[��n�<=1�,=��<�g1=ibY==
=�G��X���9�A�����~�"�V���$<�\<s����� ���Ƽ\*R�z�$�3��<��=�=�yr=���<��?<3	����3=ŭ��$�����H=�6���,=��=-�4=Hk��nAͼ�X=��E= �7�qWD=`�� =�͂���W�	��<J�1=Y�{�i�=�}C�$=�z<�r2:���?�<�8�Jfg=�kv��뺼hk7���=A�����o=m�=�j ����<p0�Վb;CU=8��<��5���Z���.<,45�`�=��& 9,;|G����J��<�~_=,Q���hT<#Qj=������<QG<dߖ����
�-�mw�;�={�c�tm�L�!=�p=�WH�df�T�<a��,Ҫ��~F�kzW=��|=�!
=��]*3=Ԑ4=6��^b��Yk�<шٺ�x=��;<.�U=�V�<��$<�C�<���;W�;#,�O�=nr=$|?=���Vc�m�a�~�c`�:YA�-U�<��ɼj�����4=?S5�cǮ<��b=�?t=�<�'$==���
����:t[=U�9=���<�xs<�J�<�V�;�5�;�}<l�	<�CE��X�;,F���I��[�0=:����f=�c'=�$��q=J鈼����}���rt�:�C=�0�<��{��<�Ҍ<�g���J�.5����{�=�'�d�<��<sm^���\�Z�^<���<Ѯ��42<}Kt=��2<�#;�9�; OY=�/�;�K��:�=\oS=)Vϼ���<�qG��b'=)Y�;�#n=8�����Y<.�*��:#��a��aH�<�cV=r�<QU�;�^�
����<�o��=�7D=�JD��b��c�߿3�t&=��U=��뼄z<&+ռ=�'=�=C��?=)T=��=�3>=H�9�,�#<@I�<�¼ы.=S_=�g��E�w�r�p,�<0�1���==���B�=������ż�����[��;d��2��L���<�G��En�$=14�<,�=�y�T���s8��Y=��<�a�Ma;M�#=I6����`�!w���l4= 3��~�,0,��y�����<R�=��J=���<rV��� =�p{���(=�l	=�<��ȸ��ҼײƼ�=һ";��j"�����<B^0=�R�<Xz	��B8��e�<�8:�5[C<�����+!�<��=-�<�}�<�����0����r<�n�dE������?V��蟽�(*=�f�UX�=�)B�=�s��U����;�o =�@O��;W�=N�<UI����[�8=b�<�Y+$=tټ��E=j�<
�{;]�=������ռ��׼JSK=�R������F�<$�6�d���t	l;��K�J눽�t�<j1<=/��ѥ^=�E>�-�Z=���=�.�_�����I��Z^��̆�
�+=�j���0=�
�;�#�+t�W�~�f5�<���r��*뼔%R<(5¼h		��!��QN=ma=V��<�|����&=`=��@�#����`��Y= o�=jS�<�!f=v��5]{�� ��p�X=fd���
=��=ީ;r����Q��n����J/��+��
/=A=�F��P�;e�ͼ�,���<�Oػ,9�;�Lڼ�q�<�J=Db��.I�v�M=UJ������@�˦�;{Vv��ݕ<�<=�o+=��==L���@<�]<BB!��>���<Hˣ���=Q��<0���� ~=�G$���͹P��+�<ʹ�<h�=���<��ϼg�w<���V���`=��B�i4��7�Q<��8��0�Q=�Uм
��<UZ>�C=��m<�'<)�B=c74�����6�L��h�v<���b�[�*�R=�4<�*.=�y�j�Y=054<�%=k���ߧ�$ZB�g�"=���<��=�;�;��:=���j�;���]�< j� ��:�v;�=�R�4��}I=M'���v�<d�r�p��4�=r��l><�dk=�5!� �<�N�:���<~
=Z��<y=��O��'=�U�	���>��<��<eQX=��;$��<�;f=���;�'���i�
��<���<,r;;A��4!G�x�=�P�#���`A�<�0q=��=қJ����8�PƊ< ��DFE=p+�R0�6�ܼ9B���1=i��:�<�=��	=��-�5=�$=���<��L���<y=�;WD]=��V={;�^���T�<'0=-�(�&��<%�<>��<X����L	=g3�����?�<�v�:�dA�Ax�<���<����D�<�x7��t�|�<<|�=O}s=��ɼ��߼��<Ļ�<�_.=8���>ļ��;07�<�o��=�}9�,�]<�� �?Q�o��<�<:��(�Hio=�dm<Grh<%=�L��9��L
\�_������j`�^�<.fQ=M��<<��<���;y ,<,W���=z����$=�c(��Y\=W�<=1��<j^�<��<�Sp;R��]=U=��c=K|�;x=L�
���b���y<���rS0=U�7�%����<��<�,O�2�=U�Q=�����,=�%˼���<��4=�'ż�AC=�EF�<�ۼ�7Ǽw��9��Ƽ( =�@Y<��=Y�;��ź�?C=if3=��|=�+�T�=�/<�� =��O=m�<Ѯ�;~��y�<�Ǝ�l��,�:�S"�7��S�y:�pU<V�4�r	�:�b����<���JW���x<�v=����-�Cxf�0ǒ<�$��;f�=ۏ�<�t��
1��e$�(= 8,:�'M=�Z+��C=��8=��:��G=��T=��<�H���t���#�<�ϒ�nlA���|�3�Z�Wp<����݈=��4=���k��<v�=�Cc���3=��:=GK�=6VF=�GX<�|�\< @�j�ݼ$�:�R=�2U=����;��,=W
=�C�<���u��<1
��x
�<���;.4����<��\<��I='/�<�-4�1�<�R\���|�}Ż�^�m��� �ē9={ =����:���#�]xl<�P=�4�';bZm<e켄ȩ<���b�%�`=}��m�={��]���"=ӆ=�ڗ<�o=۟���V'=�U�=>���1���X=�?<Ri:�+8�UP����{q���<ۗѻ� M�$�a=�w������RS	�i+ļ�
�(�2�����+=� ��d�< �r������IY=M��t��<F�� ؅<9�@���=025�{7�<A~'=����fP�w�S=C�:��f=�+�7ǟ��O������=U=<��g=�=�t=�vѼ���<��u�)i�<��J��<,����CC<vs$�~���a8�=�<�$���`=���Vy<<J=J8O��������ݻ�0R=�Vv<B�<�?�ƫݼ�a������ʘ��k=��:���<
��<�^n=ob���z�Y�<<r�<W��<�:�<� �<F_'=+����S<VN:^�==	B
=I��<fꆻ�Q};�.;��@=��^��<O���o=8�,=MAA�I�x=RMּ'����S��L.=�����$����<��ϼ!y�:�n���<ͷ�=��=��"=[�<�,=w]<��[<g��=��Ӽֹj�R&|=�\;�,u<�D�< �T�Z	��%E=�*	=�O�#v�<z�;�B=r^
��ݬ<�ω<��2=:�<_=��)<���W.�;�D9��.w=�/<����2/=Q��;�
���<����2=��T<H�=�F���;L<�;��:��3�<��G;�	�:��m���<�=�<�6#�oK�;�S=``E=A��<�4�.�x�[O
��Q��ĕ�B�0=_>+��{=gbG=����?�N�<�U�-�6�|�r���ڻ/�#=ܒ:�[&h��,ǻ���6��;2���a=M�=��S<��;�^�����;���<k%�a9�W�<����O�����<
�<��=G�i� <)B������c#��,=C��:Qh�<b��/g[�k�-�<[=佛:u�4�
>ļ�^q=�|����(pF<�D��"$=�D�W0�8�7���Հ"=�!z��n��	����鼪�=���½�<� �= ��</�r�h��`~���c=z�A�ט���qڼ
��<�$=8��<G��<����9=C�C����<-�+�a�!=`��t'R����<"\O=�K=��<��뼕�:�q��O=��m����<|���c��;]8'���?�	�8���иm_��ڵ[=a�	=g�m� :<^k'���T=)����=��<�߁��4���	��� =Ee�<��Q��K<���3=��p�y2��a�7=l�)=�3�<sT�A���e���~=,������<=+;=��{�Z=)��<�ºF��:n �E*���M��X�<֔H��:5=c�`���<X�=!�M�1����3��{=�勼)A+��h=&���^���=�V=���#1=��=_�z;��+=	A=&�����l=) `<ڣ�<\�ƻ�;���i���;܁�<�)<�p#=c�*�oad���Q�K��<���=��
��8=���<�2
=݇�<�F;��Ӽ$w�;'�C��T�(�.;�11;��Z���L�<s��<4���ً���ǼE'�N�s��꼌6w<���<h
�<�9�<,�<\D�<�J�:�h�L�H�E|��1O]��	�f�v<�H}<�D�f�Ņw���<�ma<�p�>Ӽ��)�^�=p�F����;�F==]~Y=�D�=5�=�/л�RN��2�<�i!=�3 <�9�=�z<Q�<��@��ʴ<v���I�	;�Q��jS=��Z���n=.�ɼ������o���0=��]=؍�U.=N��:���;�)��(�<��Q�	ۻ��y< b9=&2��↻ 0{=�\Ѽ�VY=�}�<Z	k=9v<��<I���}$�<A��듻iW=c�
�>E�>�׼��żB�;	<��0=~۹�S��D�N�,�e;�4=�hT��	��nɻw�C��C�Ӣ��t�;4=���;��ѼD���7=K%�vF+�<	V<	��;!O=�5��*ü�p)��;�<��5=�����rX<����2?=-�=�i=�c�=l�S=ǩ��6��8=nE�;�"�T���p%1��Y\����<��b=��=���;r.�<�2�[��<�/��м�����c=m�;�*;h�	�+[K��d=��q�5�$:3�-=���;S0�x��<�
;�2=Ѽ���N=�[=�%���s�<���<�xo:�r��w��bsA��6�<�a�<,f=y*=(�~�C��<�;�	��QR�`m:�0$����;Z�0���};g���+]=��^<�N��%�
���P<?ٛ;e.!�9ۄ���<��0�q�1����=��e�>C����Ǽ���<N��R*=f@��*�.�j`)=ʟd���-����<+oY=4�f<��3=�yN��|�:F=b$<��<�Z=QXU<Fgռ�K@=�a��-]���఻~.�ݜ�4�=P�V=���<�M0=��D:�QT=��=�����[=�_=�����Х<Z��<ӵ���C=/l����E=tā���<狀<izt��:�<�7�=<<�=�gG=�����<�:����Yu<��V�,Q	�-]'�u��3�1=�0=�@M��t=�üM�<*�;R�:�-�K�0U�=��<��q��D+�	{,=�N=dLȼ�8=Lټ�r�e��;�e=P
5���=</B���\=�ę<�^ڼ䞏�9���\<�J=����<��R���`�X伯���9�<$��;��f���k=�$/�$v�<����;�=�&�
�V,=���
�<	i<�,|<L�<�F��=�B�<�	%� 5<���<rJ�;�����a�<B���v=d�#=�_�� ��tQ�V�"=�s�=�XK=]�T�<�c<T�m��<����M����YE=VQ��^==)S/���f<��=�-�=a �<8��<��⼧�l=�0���|��%=�<�;b�0=��ټ����=�о�TRU<�З���<���<ؿ	=�>ļ$�K�=7�<sSn=ZA{=����3�u�+�RE1��Ȱ���Y��;F.�Oļh�<�x��E�����G�\��>�����<�6=IW��%����<��M��S����<�|o=��J�ڢc��M�h�O=�ja==�t<q��C�<�\j�g���S����52��!;6/���o<��yR_=2�8=c�;�� =���[(=�a=��=�e�=)W�٨)�0y���ga��	�<�#����|s��I���;�-h=�T�<�b\;S�S;�P�&C=8(�҅-���2�x�O����<�UA��p=%:��G��nǼ興:w�i��s<�A=���;O�<��U���<��0=C�<i�J= *="� <�b�<:Ȇ=���[=��-����M��}K�5qO�꼥,Y��e�<,F�#�;�/%�-����`{�Ե�=�?�<hl=f,!;� I=��2��R��7����������Q=�z'=i/޼�[�<��T�D�W�n�;M���Z@ =����T}V<D�<l�|�MM(=�؞<1̃� #$<Ñ��'��e�+=�`<���¦�M���U= �<��#<�=�9M�G=-���p�%�`�z�':U=-����H=� Z���~=�o��p�k;��t}�3�<J�鼼"=��)�������\=���<3�Z<�o7;+��r���w2�mQ�<t����:�0�<j��-J=�����K�<�����E=�',���V=�	)<L�<�eL=%���줼��4������01���!���E�<�_=�:=?7</��!�����<� =��<���Bkp<��=d���Q��7g<~���`�ȼ�=�¼ʐ=�H���0��C=�?�<|�7�����/߼0��4��<�t��}<��<�U$<�/>=x�)�FO���6,;�{#7�[م=�Z��2��R�Z�a6=΋缐�����RA�Mm<�^��}�=�0=�ҩ��צ��>��o������=��O��0=��Ab�C��`��ɤ��.k���<��n=�WJ�B�=261=x����(ӹI�[���<Ζ%�:���"=�g�����q�x=�̻0��<f���ˎ=�b��d�]=��<S./��_X��t5=A7�;��C�*�o�W=-"���@A�Kz���˼��<��R��h;єj�U�����%=-=^�h����Z<�Y?<!S �7�H�ZS��6Q=q
ϼ��P�^=�H<�0]�`��~[==+���μ{_<��ּW�<���M���-��_e���C�}R���ߺ<e�-�}.+��)m=i���C�O&<{bS��W;��[�Uz:$=��6<O=d��f;g�=2d4=�5=��]={��;$	S=�a7���<ݲ7=��%��.@�`�Ҽ�[$�Ψ�Z;�<��;�w�GW<Q�漆^_=ȹ����K�A�|��桼��=-ӂ���H=1�F;�=�YV=N�>=�?���F=}�_=���<��<�孼� 4=�U��~m=*H�<G&=�E�<;�==A�� &��k�<���<�Pt=��<c�U���<?tz�����3�����`CO=T8<����� ��Mn��-)���h��4�I��;����Q"-=[)���T=o��}R@�k����:!�!���7<��T�P�0�=$��:!�<��=W4=�/=m3�<�qk�vE��<����<�a�ڧK�?�0�Ƚ�<X�<{���*=�M���@1=�8=�f:��ȏ��;�<��h���<oP�W��9J� ��(���\z=#%���<å`�w�����<~p=�H�s�!��u����_��b0��M�<���~V�<���<���<�J5��?<��<���
q=t�<o�I K���=ǘ=>�C�� <;x��?��=X���<8�/=>�0=I`=4u��Yʼ<��o<��ۼ���;��ݵL=�o�<����f=q�7���!<��:��썼��<�c�<
��<\�:
���4=�!�=��.���;�=�q�'}&��3��Cߺ].,=�{T��0
�J?�V�<$N<�
t��˖:H����D=d�-��#ἑPJ=H�5��__=��aiC;���<�zZ=��<4��0�4�Sl*�����J=u]�I�&=��<c+M�x�Լ�	��|�<��λ=t}\=`�m<����{@*��B:=e�<��t=�=�޼�����i%=y��v�[�l7��P�D<�=PV�<U�_�����@��;�n=^���Vj���ޣ�U��<dz��9�����<��=�@�=V�0=H4�f=׬�^�:X=��=k!�:G<�徼`¼�dK��E����G�E�����*=�96<������	��^U.�]�0=�<�#�P��$� ;�<WC�<ʧ@=�۬<��c�瑼mq<e0߼�A��4�S��
�/Q��r��<}��<�C,��@<�û�S���=���;
Y=�	{��<ڐ<a^�;ٻ��)H��<�:���<6���--ݼ�ർd�ؼ�:X��h�0@��<�a=�u=��=�A;�E��x�~��K�����@��:ګ���*\�腙��#=���<$BA��
� [X���;���=f�K�j�X�K}`� ����6=�L�<�X�Й�Q1a<-๐��<Lu�=AX3<Lz�<4ݦ�b�P=@K��뇐<Źc��A�k1(�:=��=��=\��"2=4�ļ^j����-�9;��������o���Ix������<�۷���<2�*=��k<A�A�ٖ3��G@={_�<t|;�.��<�ܼ�cʻYEt��	L=T�<�[�:�������<�K��KW+=��A���ؼ*�7=H�;��3�Q��X���ׯ9�%1N�� s=����Z�6л��'<C}5=xn�7�;�� =�[=hL9L�=�1�}���^=��U=��h<�'P�|=�@=DD��π�9��<p$j���Լ� ^��u�<:M<��=ʯq=?8���pv�{��$�5�WR=��<Ʒ�<�_� � �+��y��=��� � ��X=���n-=��8���A�(c<�fH��j�#. =d� �ޤ��d�"��1W<�<`wq;����	B�R�|����<yl	�� �<y7=���=�.�)No<��#=��̼��'���^=��|�q�.=�1(=��]=!Ex�e*�<>�=��湛�ں��=H�	���'d==�V��0��'ƈ<���^f���Y=�y�<1V�;.�=��(=�rc<C�=»��3�S��*|�/��4�!�V� ��B�<���϶+=��<q�l<qS�:A�"��=<��d=��<e�}=�=�<�"�<��?��}��@˼E[��v�J�NW��h�z��.-=��k���N=�(�:{���ٱ<� J=ø�<Y ��>��3;��e���q�M��;���<!�ۼ�΍<,o6�\��;kg�<u= p��%�P�Iy=�8@=��;����+�漣�<� ��%+=-U�<����z��|�e*=_m���&���Ǽ�3,�&�=�;�9�¼�c=�n<�0h����;=K~�7&<��E�Ï=L�7��	��6�����<�n�F ��ޓ<^q^����<P�
=�|<�!O�;�<���%C=�9�< "j���\���4����۰{��ly=��F�����<F��I�A=����~Ե�:�E�.:�� =J�a=�=�f=>��^������x��L=��O=L�0����;����e6:�i���f��<q��:��8�w���<i��
'���Aw���<̮�<?�W����<�7�����,���#= !D���+�ǩ1=]A=�d��%�F�*�_�:W=�D<�D�<cN�<EJ=m(��/Z�@�i���8=*Tc=�?(=�F�=S�~��<��6=�F<��M����^�9�$Iмv�;�o=3�9��Į��d>=��%���,<̶�<��<,�;��<KTD��[�<�"�O&�<P�̼G+��>I���#=Y];͂ռ��;�=���kN;=a�R�ܼ4S�:�ܻY�:6�<�<\�<�E�w�<�2xf�����h�<}z=��.<'��<��<`ռ���¼�}m�+�;Ғ̼ty9���>�1=I�@=4*�<�쾼��J��; =c{=�mP=���<�	D<mՇ��~ɼ
�=E<=�<>n�1t��C�<�ἳ�=c���L=�$���0����г5=�H{���O�W�N�i����T��I��~=�6�<�Wu=��\=0fY=7� �,:;�t'=�.��I�<�/v��F����J=<|� =��zÇ<CN8=N����%��S�D� ��=>�M�=	��<^�[����/�ܢ</�Q=s�<c�i=�<�C'�ȝ���Ϗ<��<�_��9<��=�
=�XP<�>��3m=OL�<��<1$ʼ�g�=2
���P�<u����Eob�_U�<�Ȕ���=Fv=�-�<(n2��;5=��"���Ƽ5�2��<�!v/=���������p=wo4��P�< 9�"0R=`��<<ɻ�Z>==V'�9%μ���2缧�+�,ǂ<��`=��=!F:��C����a!%���<���@>r<tR��H���;H*<ذN=U���j���BC��=C7D=,K꼴"�d?w=7�<f��<4u�;VdK< �q<���=��8=�V��jH���κ�+�<
��<�k+=�2��GJ;��<�W��P<�=��:0��v"3��3�<~�7=����C��8=���Sr�;?�0����<��[���<�u*<�F=	�=�7���j=X��dI�<��5<��<�[K�_�=���<#%=�mY�o/���2<��<E�6=��X������T�+��<b�<ټ�;z��=�ټ�&�<�����W(=�s�a���.s==̓.�Z�.��'�<v=��<޲I�<y�<c�9=��
��VҼ��t����<|�߼ia��`=�fv;i�N=�q$=c�1��H�B=�K�;��<Ώ�wlk=�����@=@	�aj=��b���"o�^�F��=�S=�ˏ�L+���5���<��<A26�h硼 5~����;�k?=&�<�9W���;<�<[�Q<��b��&��F�}���X���<�^�BY��s=�)�<(
Q�� ;�|2=���<��@=(�*�=�����(��&���J6�#��:��7��9d�$BS<�b&=���<��v<<�m���@��=�^=k�!;��ټ���:�m�`.3;�j=Q,<a�ļY9��-�K��̷;��!=�3˼g��<��Ӻ�	�P/��g9+�3<W
�$Db�Ñ=�^#���;=4g<"��;��5=��<� =&�E<$�L��<��5�(=��U=��Z=��k��P��:�<�K�c�=q��:?��;p]�-쪼�q����<�1�)�;��I��b�<n~�<�����M���u<���D��(d�<�$���׼��,���=L��D�D���=��V���I�o�g9h�<;��;ig�d�~=�p�<�L=Y'<�����;O���e�e<��T�z��;��3=�W.=�U�<98=#�ƼI��;
ټ���<�^%<��&<��n��<�ݼ�d����i=�'=Ǜ����h�R�ݫ<�h)<ݣ���P�;��=}O%�X�=�ӻ��x�.��� Ӽ��Լ�0=��s�B4=�g;<�y纍�X="/G������n�c�9��<�������<ܫ�9t�$=-TM=��3��<�<�O�
:����<JU%�L�;M�M�,�D=~3!<�ς=�ӌ�A�m=��<$����P-=��м�X�l�=@��<l@B<�7�
s���p�Xv=��^=���� �.�/��<`=�5�%�U�$-"��X�l�%=-�<&vp���Լq�u=%�
<�f>;y��(x�"_N;Q���Ӣ�;�l]:`J�=����0"<DbG�{A�<�@T<z�Z<��!;�=�<c
�&�#8��CՎ=SN[��1*��5�<��N;���<����,Z=�1�<��s�c!U="μ�߻�5�<M��;�f��p;C�ջKe�;��&=�q<�K�;�r�;	m;�=�-g�D$��3P���<v�8=���)=?�Q=��w�ϓ@=��V=��)�|+�;��)=�A<�V�<x�==�(��x��g]��W��:ܻ��<.�L���;��=��=�5��3J��:9=�9z���#c��Χ<�����==�;M=����0����<��=����s��<�qp�Qz�<��<�|(�U��<;4�<�4=��ɼ5�=�"�C2�<?_꼽H�<�P=KF����<���kG;=	�2=a�`<��=�T�<z6�fA�;tH}<�s@�>��-��l=zf�5%:=�?>=p�<Щ4�1<��r���鏕���)=�b2=<�ʻ(����K=���<�����ה���u�:��<��<2��e�=i�<��z�z�K=�<��H=e�+�����y;5�=q[�<�<<��z�=��"=�i=~�K=��=�0<����ss<�HY�|����vm���2�܅�G@<�	=��=�4˼ƐG=�b[=*E<����J���2�(+=�u�rr'���(�9<p�)<��ܻg$�鐑<9u=��3�\�=���;9r5=�? �)�<x��<=9�<^#��9O�6{պ`N�<4P�<m(;i#=��.<�,�;a<�up<Q��<� �%bN=+Lp=f1j<j	��eK<���<�=i���φ���1�A�����<��<�1�e\D�yռ���:|��}��uF�=���<f	��81�J��<�?[��)C<�S��'5=ƚD��y�<T���*�;x�q=������d="���Z�=[���Vټȳ�<<h<�3��R}�<�V:����n9=�b=��^<���< ��b=C#=��3=�<��D���7�D^`��Q#=d׆����<#6���A<�y�Oy�d\=�78�;�=&O�kU"��]t=h�"=��k���K=�=��	�ٶ=ޙ�|,`<�޼������|=�=<{������<��8���w�@�g����м����}�<�L<&�=�F��4<}�|=d�� �J����=_���+!0�����|�<�u<֏Ƽ˵=~xg=7a��y =��b<hE=t���u��-�V}üo�<͐R=��
=��v:@���&=m��Uߊ=8�*=px�8t�i=���[m�<1�͹��л�T�<���X��wּO�+��r==��q;�u3<�Qm���7��ZE���`�rXL=�n@=�bH=5�Ls�40=�����<ED�����6�<��= �E=3=�0�;�%E��="�=Si�:�!(=/���V���5����	��^=	=�9Y���!=Y����\�򼐻(q���$��d?��."��mL=�I=���4��:?=��;V����A=+��<�dм�`�����Q�O=0B<��=�X0��36=.d_=�U=�m_={0��w���	�W=&�'=����	��ڮ<;�<�"��s�<�ro;3�����=�WY=��f��J�ѣ�<~;�<���HF��lɍ��	1�m�ռ�'=C�:=�6^=�7��ZC<�*�j;��uȼ���<��M=ׂ{�ч;��h��<j=���<V�4��:)�f$=�o�<��=,�0=��J<�Ȃ��/�<dw����=�h�<B��<�N<�_�<3�>���<�wF<tT=#ql=���;��p�(��I��D�<���ы�e4����3�Ա���C��U=v�z��n��5�<�m"=��x<<����G�Y��8�C=�4�� z�<:m=\<� E����<cf>=���<Y�=��;��4��aE��w�懗�Elc�x�+��s)=O2=�)1��h�<��W���<�0=0p��
�D2�<ʰ����<�UZ��%�<��b�x|��[�;V�����'=L�]��xW;��]��ឺR夻��}��F_��Y=��A$���CE��V��Ë��,'=�Y��56=*�v�	=�����="A���=d�F�C^ <u"?=�^W���=w��B��-t=��"�����
��=0�z���;�ε<���<a;�;d�<Bܽ�&K�<H�C=��-<��������k���9�0�V=� ��v<�Y=��)=�q�<&��;��(;�N�=�j���<3ʌ�ԸF������=��=x)�<cAy=�I=�oE���#<=6���I+��=&�k=��=���;"�;�� ���W��g��^=5�T-=��;6��� λm���c��U=��<��6=̥�<�"����N���Z[�|$�<�:=��X5������4�I�*��G���-Z= ^���X�F�t��L�<��=�s=L���R��V=+@0<;�=,м������9����|=�M=��}=��:P8O���=V'��<�w?=dI<=��ɼ'~(=_��6�<�==�u���=��Y=��n����Ċ��[>�,\-=lT��ɶ3=/��;f����Pf=i�7�`�=����%�X�Y\=�V���y<��<��
=�*@��1����=�Z=��(=�L-<�-h��a����4=O�^�:���_ϼQH=�G=�e�e_`��eg��W�<y��;߷���ټ� �;�I�5<(�ڐ=S��!��<"ּvڼ�<�,�*g��02����1@�?���J���σ�(Eƻ�qڼm�;c������<o�]�Y<=���'�<V�i:f4���c���(=��ۼ�߳���J�ɦz��o<�B���$�:��<�(��Ks������]e�1��:$�G=����׼��m�2�1���=�3�;�F=��ܻ���;���<�
�<��j=�@м+'����<�a��$=j�G�ĞZ<�z�<��-=v�;�(~:������=�o�c�{=B�?�mBp=�cݻ`VO=��o=�=sL���0�<��c���(���*<��W��	�V�-=��=���;��x=U{�<�� <l���_����!<�8�<�-߼'�=i�)��,���@n<fA�6�"�b�=Q�y=�ͮ��	������\��|�;`�0=��7���'=B�R=<���=G=�=�<�������D�%=C���ڟ�d���I�q��;6�3�E�����U��K=0 ��zϙ< O=X�<����%=N#O=v����4��м�xѼ5v)� t�8t�<��ļ۝i=m4=��G��jq�q�R�<�=}:^=�����/=v:<�0=��Z=��y<��߼ƥD�rh�<3�f<�'��x�5#�:��4=iN<G=k�]�����s�5��1�+l�(L����q=(���:��AM<t V�=�-�nim=o��&��<>ռ�ļp��A�Hwؼ�G-���0=�.<=M��<�$��F�<��)=����y�=�3��]l���o=�i$���
=.��n�����<�9c���<W&)<e�N�g�=�=-�����:<p�<Ƙ�=w�;���/����<#�&�;��=�:����\=a���&=J^o=a��1#�tj9�2��"�T��6�(t�:�3���*=k̡<�)%=�H^= .}<{����]=� &���>�s�$�I<.G��SC�ˀ�<�0�<<�ܐs���;�U�:������9=�R��G���x�=��TA���)��u�<���<I!�<�Kl<�) =�%=De���w�<m؞��=���F:�s=�K@��m�;N��z�D�y�U�+w�$߻f���5=֦����6�W���I=��a=��r=��+=\|<U����w=~�=�; -=L<|r���¾�<&	5�:�,����;)�w<�lD����<6�8=�f_�Gx^<��<O��P��2�=�8=r��j������ҵ��z-4���=ߣ =럺<��Q=�S���!�K=��C�+c=�C<�=u���=�
r��:�z��<9Bi���=ő���9�p��Dsӻܟ ���V�zż�R�9z�A�:�xUr=h=��t༂�>=d=Kiۻ�'�<����y�������	��!H=y���X|ּka�;k/���]<��a<��^��h¼LY��؏<j�t��E=���<(e=�=���=
�7=�\0��~޼�~-=�����W<�m
=�N�;��R�p���/ݣ�܏=&A=L��:��>���/<�;���<F*E���+=Zz�U&���<�P<�O#��;X=���X�<���9��"=$ꟼ��7�vꓼ�<�-=��Ỿ�<Z�C=���<�F<En�e��<�<�#�<�+4���e�*�q=�q=�磻�{�:��=��Q�:8�̄T=��<r[3�
�C=��<~�;<�4�*�Ἰ�G�z��:�0<����F�="�<�HE=0+�63(�S����'=��)=��=Y.�<98V=�*���������;#]C=��;��<R�H<M�м6/H��ҼsA���I�<]*~=�ў��
�1�<��
��_3�ī|=�Z2=ӝ;����TeU�8
 �c�k��s<������;��!=�-�<�b��s#;hd��M�U$O=x���/�b=�n����\��=��<����	�.UO=��^=��<���������!�<r$�;�kh�Rܐ�޾<�< �L�� o<�92=��
�+�;���~8�����;*�
�(y3=����q=s�<�JI�f�]<�/|=�%�u�I���=�=<�CF�W��'Dj�{>u�x�<ü�8�}�=ڭ>� �o�Sj�<#6ż��H<0������<bߔ<$�<�3�����<��.=��:5�;lP�D�=Rt1=ȴ!=Hҟ��
m=�6<^KB=�*4�W�^9��Ƽ��_��e���L=�=���<U��36�kr8Z�D4����3�пb����<�.!�Ǎ��䑻���p.u�De= V�<���q_��dJ���#�px<5=�S�׉��{=��T5=ŉ���=��뼩:�=UB(�NL��eQ=��?�k�o����M�T����<�9�<D��<�I�<t�U�o"���=~�="2#� o�<��쥙<7�8��j�V}w;!��<6as��6@;�=�@<��z���{��̲;f�B<��;���S=������N�8Ǽ���-��<C��<�(
=�<=p:�?�6�\,~������H*�@�=F�X���Z=��Y��%#�z��:���<qhy=��\=2�*=�Mk=7��� �(�;�R��<1����n�;9M�	l&�
��<��=^cK�w�Լ����ÀּÛk;<G;��7O�J�𼍫�<�K=2�8��t=�l<��`���=tp�I�6�s��� =1=.�+=�=�>��"�8"A�s���^ɻ�'D��
���=XOG<2�=����Q=h�s�A7~;�p =��={o�<is�<b5.<K�9=�y3��c��+ih�X;�=�=ք�<��&�<\�<�}d;�kT=����9�;���AY<;b<�0j;��伤 ���=Kq�=���Sa'��F=ۧ�>�,=Z����༿�|��?'�<xw�~�*<S�-�K+��Hy</x��I�*<����/k� /I��Ѣ<*s�<<���܍�k�<=c��D�[7e=� =m,�����<"�;��R�W�K��S��^=_�мe�<���<�A輏4���R�;�<M�,��}��<" <=���i�K=!��X�T���0�F��\=x�7=��<6��<j��<M �<#��;`$&=8�I�m�������<���;֎<^��$c����;/���1�W=6W�<�O�Y��;A���G=7�=Ƣ�<�DT=�J�<8R�;�!;���<��\<��t���p=LU=z��<��;�������;��c<���<��\��?���/=ȗ�l]=ӟ;#)V��B��J�Q==�� ��ѻ��;�4=�0�<O�;7p�#v�<�{��PHO;�@;�J�A%Q=��<�,H��p��0Q%��'=]r�<��<�#!=%,��ۦ�1�H=�1�~�<�}D=�*=�3�]E0��ـ<;���cͼ^�=M,����E�d��=���=s1�?G�;H�a���鼱C���^N�< �=�!��2=���T�{���W<N�����t=��<e=Y�ߡ$=ji�=�q<Eh�<J��<]N=�'�<,�<��� ���{u�=��<�m[=��<j��@�<����W����^	��G=g�<�R�wv��,�r��oj<��:�H���=8k�;�*/�.2=�k<3��<b�M=(���bX�x, �-�T���i���<��<��m����1^�	 <Vn��z�d=K=��C=�R�d����꣼;�l<~*e�<�Y=T�ļ�/��/������ Z=(�P�!7[<;m�J f:B(�<3��<R��<��=V�9��;�<lj7��T��*�9�D��_!����8O����Zr�/,T���1�ڌ#=���<nU=��F����<!��<����7K=���`K;<����p�I=�#�;����&q�<Y�R��,�<�^�<r,ͼe���t�=S�t�:<�
�<8�<�μ��<4��<3�.��;<eL�<q<$=�����5���P��U�����=ɠ_�3����|�<�zǼ8�=ĚN�H��<)q<� "�t�<b��2�`<�=Sj�<a���Լ��=��W=ZE���:�<��<�����<��nG(<��S��^� l�<�t���~w=>r��-�O<ؔ���C�eq���X�!�8=r
=)T�;�!���E=�k6=�]=��W=T
K;��:>N[�,�*��漩 '<<����=���<�a��󲼗+=E`[��Vu�!H'=�w,��> �$*�=�`S����S�8=Zr:=L�=��<��^<۵���T���;�����MYV<O��<����&��;7�=Rg9�pQ=�=�A=�{=<�5<s�=�A���n��
�����0��r�<NО���<���Z�K��P伽�v�h>h�T �<�t-�g��;J�E=<�=���<�HI�R8E� �=�*h���=�j=E\��#�0=$E���/<�-W:u�z<��,<����۩f�g=�a<;��?=FMj;��</�2=��6�>ԯ<%�����<lY���|�]W=m5�W8���3=F���x�<*��<%����PU<^
��l$=�A/=�j�<���<��	J���ζ��;��м�t��DC=���<.�<�$���4���������}`��7<�����?=��
=#��<"�Y=�-�;v�\����<�屼jg<@L�4�B�ƝG�((��A<E�#���=1�л�͖<1�F=Nټh�/��m�<v'9��U��ف����=��"���Ǽ�ձ��d�<H��EI9<�;�;L=��[��������w7=B2&=��d�g�"=P&�<,\�;Zr��Տ!��l�P��:]��j�����<*�e��<i�m��*��]�<^�_;\�-:3$o��=]��<�+D�i*�<n��<Sq�C	=�W ��uz��w ��l�6!��6,<�~W���<�8�<UJ#�M݃�=Ʒ��ڔ�\�P�r����c�튆=4�6=�Ty����Vr�<�`��QP<G�</�I<I�#�}��v��q��(�!��t>��f8=�x=yP�0=e V<�X�:��;F�x�C�n�k��1,=�w�"=�����*G_�1�=4����S<m]5=�#�7;�}{�<�&Q9aL�;�L�<�Q�<]��ȴ-=�H]=#�ѻyx9�Ӽhh1�,==�
E���=h�P�h��Y�0��j���@R=��\���λ}�W=}Yl�Պ;�	�A=���ϿR�J�<�ނ=�e�N�2���<e0=�N�Yd���&<�g���S�T����<��@<���Ë�,!�`�=['����$��щ��9��<Z<M����T=E���b��Z�U�M��&���ü|�x=�t�B ���6�Z?Q�q =���l���f�*=X}��K�<S�<���<<��q}_=�$X�!V�<D1��vF��ew�G��<)Eq9��x=v�l<E�<L�X=,<��A��%=���L��;��=�5=ɿ�<]%Z�?[�3�=�>/��]=.4�
	����<�QV���Q�Z;� �/=�LQ;ߊ<��6���<�L�;��<~^�&q=��4=���<�<v�=w�<�(���T�B<=Yw�<��<��#=��<�3��W;H�Ƽ�5=z3�;���<��c=-2=�\�� �<�@:.�l��Q�<`3��;2=8C$;�	*=��<��=��<0�=4�n����:�n�:�<=<��@<P]&<���<y���D�7=HO����w=��<<4�Q=dV�}�"=&�żIvs�M�<��3=�w�<"�=���<C�<�9=�w�Q;U;Y/=z��
�黀ː=KS�<�(��;=1fc=�|�<�z��y� ��<�P�<�p�<�d�EN�<��7=Z����켈�8<�u�|	<�h\=5�F=R!��&�<u�<�!�<1G��{�<��̯����;a�B;t��<]	,��� =g�"=�5=��<f"�<��<O��;��g���<uVr;f<���<t=��=_���������� W=�|��A��;�����N=�mi��E��7�=x��<��=�*5���L<T��<o V=�_o=�ؼf�<>C!=��^<%Di���=�t='�;�Q�^oY<���<�N1��<aI�C���<
X</;Ａ"=�+=�M�<�%�V����?=�������<g�=��ͼ�=e�=Ν:�q�
�8=�<ᭇ�b=-;[�YƱ<B 1=7)<�=�G���	���*��`�-��e�p<��;�'��d�<�i=sS��v6&��w~=�h=$a�<�
Q��Xi����;Ɵd�j
=o`"�-:�<]a;�{�<��'<�(�<`켼���;aE$�=� �P=��ú}Z=m�="�����X���7�<���5�Ļ� 8=&�&=ˑ�h6;��:=�D=���;U�=�H=�ʼ׽+:�D��l=RG�;85�<�~:���ü\͂�C��V�<=)�]�vv)��6�u�c=w���K⼈i�:�rx<	��.�v�!�
��7M=j��<U����c�	(ٻ0�<h��<	��<�m@<h�#�0�H=2���'=T���:�c3�rHr=Ӝ�<M�<+=<S弈�.���<
�><pZ�3<Y=�*%�qQ��] �o�%�M�������=P�;��|=)·;@��<�E�����Z�<���<��h<���E6*=VE�:����o��>ۼ�A����c��%<\�<}7�<a@/��+�;ٞ;=|c��9��w�S=C=�i��幼ɅF����;�G�#�_;%u��Syy�"�[=�:�<h�����<�y���=ݼ?���LOL=��㼯��;������#�6�=H�)�ݡ����;�u�=��M<�FK<�[�<�nQ=PD�k�"=ê�<==W<ik5��<��^=)��<��<�e�<�h��!��;�1���B�O"<6vn���ۼ�6�<�n����T=�3��Y&����<L����׼�����0=}a�<���f�h��.7=��F�W�ż��=0X��� �=�+;u�N�C#=m�7=(�!=�2�<s<�@9�;�[=�V����=y��<j���:�m� �������F�z����-=>�<�I�;��û�G��jG�<��?=( v�|m�<'r�<X���'=c��<�e��2=Ȕ�<��}=��<�ex <){F����]�!�_:�B	�� M=�d<a�2���A��u�<lAC=��;�w=E?�84=8�<L�`�=tԼp��=�A�=~�\��#c����9 �`<�Ol;gp,��w�<oY'��ԗ��"�<z��=�L�Lp��������$=8�N����;�=�uT=�&���<{ؼ�F���<���;H�Z�!a<��t <,n�<��|]!�d񈽾�׼�f���c=]�<����iD�ּ�޾;��<��;+�`<u�Q��H=�,=4
��O��<�<"f�OM=Px���*Ӽ�~�<}5v��=jnK=]�<V�t9��%H�)Q�������7����ʼ�M	�yܼ`�Ժɗ�<{cB�]����%�b�5��e��_�����<��{���r9�!	=�_'=i?Q��=�;�/�?�7��r=����i�|�5��~��4�l=ON���x9���X,=5�=(iE���E���4���UZؼ�;�و=�[���@f=�O����/=���ļ��<Mmu�L���h ?=��<u�_�0�=,A�=����Qka��=S��=uVj=`�8<l=�	��+μ��V�w�J=^y�p	�<e�/���<p��
~=xY���B<ğ̼�nn�����<�'��>l:�NB�f=߻!�B:=]p=7�<�3!�n �<v$=�v������cu=�=�-=eB5<�#��^B=�j��)_������a9<��#=P/���-=����M=ؗҼ��B=�x$�'����<�̼4 �g��;�if=%C =��8<������u-��=�=6=���;v7�;dn���;�ޟg���N�#�R�Y\;���Z=�	/���<�f5<h�1��8�v�;���;-I�<�7A��<a`&��s%=�>]��we�~2{=���<c�nf�!�<"���#@��4��@<b�g�(=q=y~�������j=%v-=���<w�Y�\�G���i;��"=�G�n==DM��:��'+=�>=/�"��N<�(���p=�]�<��7�E�E�`3�����<%[K����<קb�Z�*�&sd�m
�<5��<�I<�	?=b�!�����3�%��J�X� F�T7�<d��!e<�&�<oӼ��C��CA<����B�&���<&x�:Ě޼g��?�U=a�=�w<��<��M=�0=�K==��=�O�aAA�IA=@�!�MB��1�[s=�a=��f= ��<؛c�^�n�w��<
�<=l�w=�K$<o#.������,<��<��z�+�q���
=ء)���`��j����t���
���S=�B4���=��=��;�*�<%^�� �<��H������2�A���LVg���=l�?��O=\�<A�'=��-��j�E����'μi z�,$:��h�<�V�<z�<���;�;�Ա�'������<fB<��7���=����q�;- <B����<��<v� �p;»��<������<��n=��=��Ǽ�"e�Ŝ<�]Ҽ�=C�G�K��{���b�F�_'�;v�<�x��̻���"�4k�<�,V=����7�F鋼D�o= y$�Lm=P�.����<�}W��E���o<-{z��)���bɺZ�j<��=��<�5�p?���<��;�&>�l�η*= �<��=��-<c��<Ld��rQ������.���J=����$L�Pb���<�gO:`�;ST2��]z���=�ļ���;fl���)3=+'��B)��ǂ;''Q����G��<ܒ�<����Ǽ*U�<�B#<a�='_�D|���=*�"=�4m9`jw��
�e=�<����u�>�/�,��<�e<�@X=�=0��������f��7���ZF=�W�;��<)��9=���$-��˾�A��<L#�<W�l�`�켫�B�	EA�]g�<�_?�ZË<Q�2�"�:���<��r��݄��m��I=7��<>m��0�-u�:
�{�����sB�<6P�7r�<=���<8��<nJm��������;���Ǝ���H��~=ۥ�V�=�>�3�W9�f=���=�������Y=���W����8�;%�Ͽ�WB;Ǡ<��@=���;+�;�I�����Ś7�?꼽t�<��<�+��L�ٱ�<[�C��ԝ;؀��-��$(>=;O*=��=H�='�]����<~�<�Z�<��<>�=�\�;��#��<J��;N/����@<<M���9\���G�ⷢ��	���<� �:��+���<�p|���5=+�=��k�l���&�<D3���d�0�;].���y<*�/6R���<ˆ[� D�<9ͺ:$'<)��<�fU�]˜9gO�=jm�<�B�<��Z=�O�<���v"+�a�����{�W������&0=R��<�jN�=L�b�<�/.�M5!�y��;�2w=a`��o�l=���񎤼�j��	q��Re=���;��V;li=�gF���<�M>�hn=�*<������Ū��,<�d=L�J��h-<[�����$�����@=����7=�����<��B=��=�}��/��L=�1=8������<m���h;N}�<���; \��c^�O�+==s��0��C�C��ļ��<5M��D]�;P� ��<��
=��x<yE2=7h%<�7=k^(=&uj=���< ��<L�`=�:}ᘺĠ\��~�<#�@�^G <c[J<.Y̼ ��;�5#��-�dpB��|�� ��(M����?�r���Y���Ƽ��%;�A���1<=��<�g�<�*�<H.=�8{�π�z=U=6%�<�\]<�,߷XN�;�d-=�ņ=� �"���p߼�0`;#_��o���l�䈶��)�<�En=>����S��De��_��������<�恽*;���V{�cN�Mx���%)��!<7t�;�!����G5��^�<ѐ$=�/���f=`LO��=��x^?;��U��=��}t�L1=��^����<-u<������+=�\c<�5#=͎��?�@����5����;u��<#�S<�R,���=����2|=N���]�������"ּ�j�<�2�ᔺ��T=ñ	�XX��R`2�!�u�]�=5�V=yk�� ڗ<I�v<�~�<���p��H��0� =��E�R��<K�޼�a=�;~:��r=�cT=\�P=}e������������~Y��B)�G?�;C���6?��>=��I=�&�<2Ӳ�Ӻo=qx�<�Y� ��=(�T=:��<�U���U/����S���ۼ�a@���8<�3�< p�=i翼f��m%�.�<��{<eM&=���RG=��=�я���!��i�<΂�����<4��;?靻���R1�)G���<?�� ���FӼ�9=W�I��˼�0<��4<��< ��;���"`�f�,���,�r"a=� ���<��B����6Z�<b�&�PrE��/�=�`�����<���8�N=ZG/=�]<Ssڼ�a=��I=X��<�i=�W[=�S>=��~�۠����;��=��3=�˼a�<0����d`:�$=����@��o�=I��L66���<x�V<U�T�V0�<ݓ���h=:m�:ji��jV= �y�<�v=���b=)�=�ʼZI�<�c!���;9����=��=Ȏ�=#��:V�ǻ����\V<��3��L��3�y��M�rw�<�+R��1=z䠼�h���z=+� ��%=}���p$�]�Q<M�:�=��Ҽ�9A=#l��}�*����<�;��$=���S<X	9�P�.���K���i5C=�����+=8��<�IT��1C������<Ɛi�sk�;��.=�,�0�<�C.�Mu�<�-�N��<$n���b�<��f=I5;j'�<�N�<�hA�yM`�w����<N�l=��Ǹ��1=�Lk��YW�q�n=He�<�:�<ɍw<P�e=�����s==)-<�f��R'�ф{��@���P�����0`,�JY»�d�<�OB��U7=��!�-�==!�D=����%=W�
=�v=֑�2��<%Ss��~��E=�S"=���<�8�s���3�<#�)������u���ʻA�ػ+�;=p�w<؀0=I�E�q;�;���=��;�E��gP��^=[�1�6�.�#����=�ʉ:x�"�薥�=9�%�	<��ú�R=����,= �=&�Y;�*E=:-=��3��5�������{�8M�=Vd=��L���ú<샽���<�ȥ��a�<F�=�<�9�R;8|[��Yռѱ2��)�]PD<s�R�}��:�O��Hb<$�9���!<[^=U�=@�ݼ��V��!<���<gy��M�N�C���;�X!��ۻp��9�<��j�V�=�M=~C!=B����<��=���6,�LX%=
[��Bj��X<�=
=e����ݼ��<~�b���t=�+v�cS<�`�<����J`���<���DbQ���t�Q�O= v�S_=�:<<5=��ֻ�r=�K���1���<j?=^R�=�7�6M=_���3�=vBB��/�����<W�f=r��<8�������D�:�uA=k <�W����="y=�S;�K��<���<<)�;�,ܼ�ym���U=(�>���a=���<3w�<�Z=+ ڼ��<=�L=R�=�^_;�k�=xR�����&��;�v;&p�B��<��<�:R=&��=;U�<v�<IƗ<q׫����Y�/=u�%���92��\T=��<��'���4=f�y��h.=���;�p�=��L=W[<�Y�<�U��D�</�S��s=����T��.�<x�m�e���6�=�����=�&~m=��5=х<x%=�1�<�]J='�?���@��H��]�<��>�mú=@�=�B��xn=�%�;o9w�R=�p��Q<��J�r��<W�1<�uP�B�P�������;���<]Zx�C�H��z���<�o뼏+����b��9�b=�A�<@�=*�;=2y��D`�<A�<��R=���e�L�<�*,���h�����<)��d�u�|[�;�S�<��$=��<Ɲ����<:A ;���;^��<����8<�ü���<���:���<@�r�Pa:����r\�_-p=�욼/���<ݳf�z�=\��<�e��UE<v�=U9�<���<���ex0=J�Y��P'��X���<Nރ���;�@�ٻ܍�mX��#=���2=���N�8�SL�ˇ��e(�=���ҷ�~�B=�v�<d�:=��=4%0��o����㼶3��P��� =qz�g!g=F.�<{q�:֗q���2���w<|ڼ�%�<��;��=�g<���<�)�b�.=ӡ;��ק;a��llz=��h<![�<x�<�$=�^�k��<����A�<|�=K�a������E��t��<�L=0�S��(ἡ�V=204�%�A�\�<�f�<,MY=��Po=�#��pS='�x=6v�<�T<�D=��!<��W=c���,�ϼ��R��X�=Obټf�6=���<c��<���<��;{�B���1=T�=��<;�=�Q$=�=�(c���X़�8��4=TD�<�I\=&P=]�=(�=Y��;u1���+(��3
��zA;��i����ߑ<�:w=�g<��L���$<m:=z�7=�M���F���7<Dh�"���=����ů=��-��麹v�B=rvQ��\ �����e`X=b��;�T��͵"<B�,=�e����M=�%<�;�V�=4W&��FW<��i�$�=�E=��V�*eK=U�S��6���U(�j��=%��y	�;#�J�^�0��Xg=?=���<s�B��1�<W�<G?=����'<s�<����<"��8����e�?�Y<��`=��<��D���=g�g=����-���*�挼A]��(�*;�� <
R =��<��'=����i~��ɳ�g6=d���N=,�O��ҡ<*����q3=� K=^�5��5�P��<7�,�z�s�?H8��o��౼�1;|}輋�>�s�@�v�b=_f=_�"=��h=�X���<��u=�ч=}����<q�輸�<TڼD�c�?!ѼY��<Ⱥ��Q�:�ff9=�0�h�	�=��1�s���=f�.=�˯<�޷��g��D=��1=Z~޻�\�<�1⼺_.�Y:�X�̔��G�!�¼@�z=�N�:Bn��3缪.=�c3<����	=н<b[,=[G3�?��<p��:�8=��;|��<Tf9A�y�G�<�롼�8��D=�q�h�u��\^<��
7�r�
)��/l�<賄�Ks���!=E�E=��W��6��vA=-m~<0�)�Q���<Q��5~;����<�@���ݼ� =�I��!>�<�'�<3=1<��B<"��<�[���`=xûGW=RU�<^.7��+w��B�����?�S�]�����Y<WV��f�� ��;J�K���Y�'μL=3=� n�:2�<�<$���T#�cБ<�I���<�L�4��l�9=�=�;t��<��2=Y`M=	A===��d���h;�Z�<�CE=��J=Z�弭����Zżw��<�Y�xWr=M���=��.M=�Ǽ�Z2���ż��<(�=�6G<�'U=��=��A=0�s���;V�(���	���<x� <Yq�? ~<!�����L�o�*7����e�̨U���<�8=ji/<2a^=�?
=�=�A�3�<:R�<?"�<��W�u����%,=���=g񼴥K=3����-��N=$�\��W����E<!�����<1_�=��<��=��;�(���=�X�;o����$��<���<�ż����^&��S�<=o�<����<&��:��<�%#�����,=�����"=
���D�����<¡c=��<�"�:��AE��wz�<Q�;O�ۼ�H�<�=��<w�������5�X�X1H�t��Gb༩Q
�����T;(������<�m��*����5ּ�Ŏ��*�<�V;=���v�Z<I�6�>s)<���?�<�C�;�ط�a]9�=�=�S��e8m=�,&�U����<� !;(M�9;�"ͼGZ=4�˻Z�`��	=�(8�;� =0b4�dk��6��<h�Ѽ� =(�=����Z }�R�����*<�N.�>Y�B�<�@	=vd��p9�n� =U�(=�於�A<��z<�Aݼ3��<2��;RO�;�����v=������T�XJ�l���yr=t#�;�_�/�� ���Z���/<�<=a�E�(��<P�#=��żiN�Lq��IV�#R���X=uf=�M����<9ز<�X�<��=�r�<�D���6K�ޚ�;�H&�E�"�U�<�Fռ�b�=w-����l�=��;<~O2=��
��M�����꼻��<������<
��:�
O�^�;=m�{=thz���<�l�;ZV�;	-=�'<䜶<w���jW���X����<��1Z�<�:=�O��]�<p�7<�C�<Zm��!�<m����T���r=,�ٻ>�5=��=�~Q�]�S<-��<_�=����j����j�g�'=�������B�q.=�{B�}�Q=a�q}����2W���	<�$=8�<���;?�a=�lA��+�����μ��o�e<�q�<������<�e,�t�弽������<�  =!3<�]�<@���c�=�[�;�o�"j=��^Se=�>��=����)g���J<�����!h��)��wN��Sb�<�B�<���;�%�<+:=�u==��3���J��8=TD:<gu�X����|���4=b9=��l<���<ߓ�;0�n�Fw����F�9)�<��=b����7�<dD9�͖�;�(���<= ��Tb��mr=&j�;Nي�]�b�2(*��'�<���<�%W=C�R;w���,м#="��<��u��1��p)<J;��ͻ���;��D�T�M�#Ż<A�<H쀼��N��S�;Y,=�h>=�u�<O�.���<��;=�3�;�GL<ߪ4;3tj<aK���=f8=�Lg���=�ȳ������6м�I=1��<�;�BD��ea��\M=qm=���J<nH<�w�<Y�n=�	��v��
;��<>4���鼉A&=v����/=xʬ���,�a��<�G�f�]<�M�<��j:f}ܼjS=��`;��w���D���0<v�<�W=�/e��*��.伐�?=�fi��	M=Ntt�E���7ȼNf�<yx��#�N=8=�G̼,��x�=�F�]����z�����w�G�J�=�7����ٻ�i;Y����Ѽ��;*�	=���膼�����@=�a�<�8I:� �����B�s����;�T���#=��'�A�XǼ͗=�u3<K��_m6=�U�<�.�<�g?���:��=a�u=~^'��jS=J
�<�U�q}8�k�H�.����u��׭�J)9��vW��ȼbKc��U=����O~<��ؼ���<8z�<�
��G�·|���<����[��<%@Z<��9=�Tl���=�GS�I�=zn�<P��y�<��n=�j��]{�zwX���B�+<����<��;=�!=�L��vm="!�ޑ\��%�<�0�_=�YY��B{=��@��vd=�J�����<��\��mһ�<��6�yç;"GV;<Ѫ��;�c*��,�W�<=A����'�<
y}8�*���<R�=$s�*S�;�
�C1@=W�_=��J=b����[T<1UN=�?1=iG��&�<�Zl<�S!<�.���5�Κ@�Z�M=T��<�m.<�]�<�o	=��8�6/�V�<j�<2ǭ<Gց�k>�<tHa;[6c�!�@��[���<U�ڼP�-=��%=�(ٻ`�<1I��"^������8=�d���;U\��B ��&=�9+�!:���B���I����;��x=�N�<�f�<�uG=�����y�v�G=T�,��4�< �»�#�<ܸ���"=���$�P��A<=��=/�;<9��<���;��;�X:��D=���<���<]q=�!=ĵ:�~�Ҙ��3����:&P�<}�<��v����:��<j�`�6�R�l�YW=�,<_}`���Z�0>�:���3ʼ�*�oE���滜�����=<8f���+=3mQ��
��g�3x��3�9=+=S]j<��������+(�c�	<�{;�=\�t��C��[/��>={q8� �����="E���5_��Q��d~;��i='Mw�[h,=��>=�5 ="����P=>�,����q���d7=�`��[��X�E� Y�;��=P:e=~��v�Լ����x�;�5	=QQr<[�����һ��ϼ��<��K�'(�<��<p"=�Ls�9=��I��M4�hG���)=�Ї�cT����X_^<�М<��8=l�=a��o�,$ ��^?=� �;�e���B���;u"�;�&��G��6e�9��O�w:=���<J;�?�[=�+=@�=� ��"���U�0j��m�6���󻀒����n�v<f��<����7�<R	��i	�;��7=�Vż��F��)K=�,S=:y�=��<=�.C-=���<�M�!�c=�E;��&=�[; �;��'=��
���=�*=���t���YB=�0=`L�;�`y��O��'<p�����;q/��{uP�Vһ���<=�.=��<�u�<�A��<����aW=��$��>ݼ��=�T=ˡ-���<�5���E;�S�L	0=^@=.���.*��A<�d��0e�;��򺈱9=����1P=�h��1�~:)%:=�fK<���!�=_=a\���մ; x\��G�<�=7�!��<�E��Tg=~e9�V��)�Î�Q;��<C^X�c3J�J׺<c���.3���V�9?ļ][1�*=�������87�9}:��$K���ؼ�H�<:T��$I;`���f=�*5=K�&�ٚ޻�_�<a�M=����d܅<o��<��m��':=�g0��f���d=zI��ܼ\4����lp�Pa�<��=�⼇�O��:=��S=����K�������;��<\����=t��<�G�<�J?���λ:�<�}Ƽ;ǘ<)u�=y�/<`"�g3y<T��<�`=F�ӗL�cl=�@b<U��<�`=L�<���;�dI�����m<Ns��d���D�6=��<t=cQ=5�^��N��s����<��e�uF@=�H
�#�a���=�R��|i��g�<��� P���M;ʶ�;r���犑�7�S�\�t�4��3�<��H<��P��Ś.=��	�:�+�oB����@l,��F����u��!�<w��<�>ټ�D~�qL�<bp<��Ѽ�o�<`�<HY�E�޼r�H=:=`�=Q���2#7<w��=`7w=���<��U��ꈼ��K�I8���#=�C�=$-o��]�<tB0�ʹw�6Y�<��T=:y=���<Fm�=�X=�]��t=�,�����h]=��"<]��6"��"=�F:=�S!�@�=��9	�|=�s�<��\9Ɖs=��Ի<⣼�Z=�P.=�:K�<P<���>�tG�<�f%=B-���U<�58��)=4�C��*��a(,��o=��7;�n;��u=�|(<���<-`'�O�(=(��σ��W�����A��	�<4"��i<7 i;�1��'�f<�6�<��f������<m2���Jc<�CK=W�<�2��!;�j�R= �ɼf�[���4�e��,p&=S?�<(���ph���V;��l�N�[=������T:h�<�0/=�S=�`q<��<��=�%�7�y~�;��R=_�\���<� -�hB=T/4�E�K����<J�;-{���=����#��<fe	=�Oq���?=���l�*����~��<�#��3��:<�����<3U<n/-�\�����:��x7=�`��dCc�FPg��8&=�s���a���<��;8���\<�Ҽ��	<'��ϸQ=��b;|X6�k$=�?���[�m��X=O�����X�X[8=��:�7u�<�����Y	=r�O�<$j�&<[l=���<���<�;*,���/���y��N���[=c��<N�u��\*=Z�=[�+<��޻!��<K[�{��ym=�ż:Ɍ<Y�<U�{��MV<�=���������1=�9=Hu�#׼��~=���<���<L=U������&O��J�<%���vD=��<a��<�o��س�V] ;7�_=Γ���<�"��R�1���=�����<��6=��>=
E�)⻾��LV =
���sF�#��<OѼGb=��,�L=�[<�=g�,<��r=���D�v<��8=GL���
=���9|�<u��<!/!���<(�Z=�=S�1�Z�o=;7���_�&�}�=�&��$��1=�b+=]�$��x|=�8;�@/��n]�=~x�κE=d�6�|�Y�2�����G<�)=|>�����e�Z�הS�`�q;ej�<�+�\�Ǽ�5��a��8P��G'��=��Z=6�:<r�X�_��;.OS�(�'�S'-�`�<��;I��<��<J��H{�<(��<��?���7=Z뻺:�;y[<M�=�
ἣ�����<�O7<$��=�='=�Ւ=~�_�ҥ8�HO�<(�=�]�;����@�;�e�Ad�����<���d���FO=$Y=��=*ހ��VN<�N"<\�=��V�ks��V#�:/�;�|�<n�<�H)<*�%�ة%=.�1�]����<󗃼�Q�����<�:O��R��K�<C�=��<�3=2��r��:�=Ò~=f�5�%����y=�n��:�����6l�<���<f��;�u���J�</)�=�<#eļ{��<����U�;,j<h��ڙ�<�Iм�#=�<�X��I�<7e$�G2<j�>=M{��i��<�=A1���"�+=��N��cV�ޖA��l��x<�$��T=J�<����:�Ӽ��=V)���e��=�=�i%=P@ļa�:SU�<f�b���O��?3<��=5&=.c��`��a�h�5��<t$ݻ[�a=Ӳ;<猁�G���9��;*ne;ǟ�6�":[�=9��G�?��rż�n<��^*)���?<a�<<��<�ӟ�*	=�0!��i��WK���=��U��~��)������;�ha=%��<��|=�V<�"���AY=;�/=��<s�0��'��Z���;�E	�� �}T=щ�����<Fx�;�K�<���;��<h�<�Y=��I�Mx���&=O�<�����=%%=����+G��n��2�<M�T����<i�?����<y�V�Cq�=�3��!=X�o;54�Pлp6B=e-=�F��"�����<5�9�!F=��7=O�=���+���p�T������J�d#��׼ '�9��W��E�窘�o��<S����~;k�=Y�	=�v�<s�L<�
c<��6<�;��==�\5�`���aǼ�[6��#�=���4�U�<�����`�Z�=������]=xL뼢^,���׼3�]=�̼��z�;M�K<Oa��i����\���(=�M��ZZS=Y�w=3�ͼ�d]�?�P<wØ<*B:9�=j@�oC �9�<;�9��q<S	+��k̼�ټ�;A��7F<��6=7,-��BG���/��t�E�o=�W���ۻ.��<����5�A���=��C�ʴ�;/�=K�=��<����)� =�2W=U^����(�M�r={ �;�%=��'�wO;�[��=~��<��ͼv��<O	=$[�<�/\�@�?��|=;�<�}�<j�:��λbȉ��*�<��+=*op�.`�b{�<���q�<�P�Y��<2��<�c����c<�4=H��<�;�w=
-�<R����U�j(5��E8=�l�<��,:v�<�+E���-�s��<�k���;���;�VT��4�= 珼�Z=oP=�ba��
=�	��i/�2F=� ;ހ���1������}^"�֑ƻ-)=�L=�=�FH=�)�� O<�p~=ķ�����W?<f6�<6�N��=��=�\m���Z=;)��F�[=ɼh=U�<H����O�;��=��.<��̼��E<�y�<��Y=�P�<�6�<�@�=;=�Cv�!\;2?��_�<X��:.���p=��b<�2�<4��<�ɜ�i�<���;����e�@�^А<V�}�J����$=�	';q����:�@�����y��o=d�<���<)������*��:�Pg��_�<P�S<��=�uM= 
M<�������
�ټ2ή�`qǼ8���K��<�!=�-=�zT��R<�"Gм*h���������� ��_��q�d�P����CC��m%;�|j��T��O�<��c=��<��H�c�<�	������V=b��;r:���H�_n�<��!�h�f=yj����<,/��1��D��]=�3!��8)=��A=Q���=��<����6���[H�<�w�<�k�<-�8=.=��=����z�3�t8=�����m�<�8=��^=�q�R3�C갹�y2="��m����2ֻ_��"q�� ����-�Ϙ�<%�=��s<��ٻ��Z�ŒR=<�<��*����!<�WD�P=�Z;f�U=}�-=�2���ؼB�<ͿO=�~9�,�<��f=4J<��z����<h���T6�<_o <��}:3YQ���<l�<au.=��/��Q=B�8=��;8�;�\*<��X<��1=T�/=��g=z/[�0�=ElP=ճ����-�'�;����=h�My�:�"+=�>�=-H<�!��"��ݱ��U��3���伌R�<M�#=�t��z25=D{��/�==���<#>�<M�=�@Q=n�a=* V�8H?<� =&Y�<p�=Sc]�t�<o������i�����9=# 3=yE��D�EG�x�
�ل����?=")<jT���Tܨ�D�8<��;|:�,����;
G=�Ĭ�f�0=?=�m7���D���H�jrS����+�$<�QO��YO�ƼE������<�ӵ<	嗼�Pe=�G�����<H%&=fC=�yY=��ʻ��̻��T���ȼ=F���o�Xk�<��мrgɼZ�~=<	,���5���W�%d�.p�<���:�<3��<����z=�."�mr/��7����'��=�J��N�_�m�\�,C��<�<*�=�=��
�j�W=8�����<$�ǻ_k =IG�vǥ:�{L�`ּ��W=<Q�V�ؼ�n=H��<�T,<t�Z�=X4|��@ݼ��<�(�<NF==�K=�%<�;=��<:O��oS=������t17����<al�<��5=�=���⟼{q�<q�@��<���mA=���<�����7=�p�w��;�!e�x��ȚS=[J�w��,(���o;��ă�@�|<b9�m��;p��	�<L�F=v�\=�H~�fż� �:�}ͼҚ���d+=�ۍ<�;a�@Oٻʬ�k�P=O��v9��ټ������u;J]�_��ɀ��t���K	<sWм{=�J�P=��=��=� Z<�C��5V@�[9="��<��)=�[V=���[�O������U=��w=-{	=sΕ���q;v��<ڇ6���^=�l��o�l�.��<�4=�=�;�|���+%��c�P���;@u�o��F������<�B�k�<0�N��2=ۑ�<g{a����{ǂ<��<�a�~��<<�<7�;�?���=�E�;��C�[��<����dD=�<�+F�������<hc��kL=� O=�E|���<���<��<<�����;�v%�����I�<j�V���b=V�7=��̼��/=������;� �Ojj��A��N#/=��<UN==��<Wp�<��:��˺+��A���m���xJ�����!�Ѽ I=�	;��!=0
 �]K�<�0(��="=���;��u��2�<U��<I��<-"����;Q-0��}m���N��+t�-n�;)C�<@�'�V�]=h�"=��X��;�T�<�Y4=sZ����<�.�����B�<�Dռ�$ּ�$����}���jA�i7�<�=��k�'*D=�i�<��V=I�a=��� �2��ż�$�����H�=��b�T��<���+-{��Ã��C%=0QT��FѼ�fq<�׻<�%ͼ�D�����G=�<�%6��V��@ݼ�6�9%v;���=Y�:<��]�ogl<��M��N=N6{�i�0�Օ=��0<�f=�����)��fX<��0=|�@�8�Y=t_��T��/N=~T5�C̼nW�<��ռ������#��z�<Q�N<|�G=�m����Q=H��"ׅ�X�Q=z�;�ą�>"@��]=E�;sZ:Β-�cs��(�����풱<�kR<�#=fG`=<�:�G���-���p������,һ��==� ����;��@=�TǺ#Mc=�Bw:݄=�G]�[HҼڍF=�4��%�;���<���#�8=)$�<s�G=�r,������<��9���мQ|P��O�W�-=����NX����<�)<�HU�I<C��<X��4i<f��G'=��<�1ͻ��<}���+$=3�k����;�1=5��<�*=ЗԼS��<��e<\�^=8($�<��4�#=R	��d/�;�%<;�=l����U�U�:=�bc<g����m�=5C�n�G���W<%�;�s=<OG�uJ%={Q=�jH�(;���<���;¾=n��<wk���W����<�<�!"��I�� ~B=2A=�`�<�0=',7���<�o	��9�OFg��7m��S<�) =%��"��I:=$Ow=�f�:"O���:<v]�2�=�ǚ�W����\�������!��n��<wWF���!�� ��w7��.��#R=�p=�<;4=��<�HI=�p=O/�k��\��<�p�<x!�>t��uU=�s=N=�;%e0�+b=�L�;�1�<0����c=�64<p�<��N:&H��oX�2�M����"w���������JA���8��<s�
��>l���i=�:Y=v_%=��8���&<��:�DG��Q��/9
�t1/<o�D;=�<�������H<<7'L�T��<&�_= �Ȼ���qr��9g��8(=�d����2�8=�=��/=��<�st��
����Z=��Z���e�hlL=dqa�)�%��#����_�2=<ud��$;���@�NШ<�p�<eA6=�YԼ��<��=�L/�,B��~^���j���<ʕ�=H�<D�<C� <, f=q�����p=Ԗ��I<a�{�=Q-�<�T=�B
=���|���<O_��qu��4"�;������<���<�ă<�7#=���U%==%^�v)�;Gy��}P�<J��<���;��\�~<g(=��<�擼��A<g<==�����%��d�=Hl����<�����<ƺ+���� ����ȼ� �W}K���3=���<���<S@"�B��<˫�}�q���(=��ky"��w=3(�<F�=��ȼ�Bu����3�j<zQ뼋^��!~<�M�9�Z��8hI����<0b<����2�!�b7=��7�2�ͼĝ;3c�=ss:�
�J����W������<	��G�`��^ =��S<��=ɞ׼#�s<�.�:��<���b7�;eƻ�u<�һ<�D��[�<iX��ü7.=��N=� ���$�Υ8���"=@}�<ْ�<>�I�F����v=�1 =�^U=�t
<܃L���=M,;.����<�jC��@�>��<~
=��<v��<&��H�;�V^=�A���+=2��aO���O��C?�쟜<`�<u-'��<�Ɨ<���� �<�Ǽ�Ђ�[$�<}�t<�!b�b�2���zᏼz��$=�;�X�G�#�Q�*�������!�0�ۼ*�ݼ�u���<-�Y=a#�x_=���<��`<d�5:��.�=���c�;Mѻƌ=6����=��v�==��N��1=C8=$H
�l"�<�]d�(d���<�wH��Ѽ�%�=���<8�<Z怼��P=umb=u��q\�V4=�j���_=i�?;�'�{�G�hճ;ѣ��������`<����9�l]Ỉ;���<�G<=o�?<u�;� �����B�x<c/��;
=b$� ��<�,;;H�<��ԼD��[�?=u��<�.)���e<�v�;�~o�I���y:��r2=�'=TV�<#W�jNa=��w���E=c9�<嬪<��<=ƀ߼�7=<�/<{#i���=[Ձ����X&S��g= C�<˙Ӽ�Ȅ7s4$�C�I=�э=��	=ʆ�;�=0=fT=�j�<N�+<���b�<��;Ey���������,�&�|�;�k=�{���]�<���?/=��=����̼�$���n:���'=��Q��u���LN�s�6�<g>��=*�;�<�<�=��Z�Q!|<w�̼S4=9���5;�*=�CJ=��<�.=��P=������>��=?�R=q���Z�7�VU<0BP��h@;����5Ol��|^�;sq=�����<\�H�b=A\���̼������<�� =�g/�Gfμ�b��hP����;.�b�b��<8_X���n<�����>=����@�Y<&(=���v��9�=�_w�7���JJ=kHY=x�7�Qc&�)t�<�Sȼ�^=���<�h�9��L<Rn<=�:_�ry���l#�����g��_ٳ<�zӼ%��P��<0�<R,A���8=����������0="o�;&�=��R�R�:<��<OɄ�Z�z<��;�p��n<�ټ��-=>�n=����=�%k���!=%���ʺ�<�%���%;��HT�<je�:zO��>_��O�<:��=������tZ3<�P=��x7=�C��ZC��<��̼��R���X�3�)'9=?�f�<�pj�Ck�����R�<��="����Y����;K�8=1����4��]=�B������wT��;b�D�=�ߓ�<Y�׼����?P=q��<��w��/<; ����A�V;;����n��y��<H)ݼ�XP�`==+S�=cs=���|:ں����[�<p�'=�U��m����%-|=tI=˼�D=�i|;�<��M����N�'�Eqq��RV��ŵ���E=pYԼ�Q =�ug=4���[=�RO�����P��/�F�b�	�ϼ�Z�0�=��<������>�E�_>�;�O}��j�<�ij�| A=�n��S=�w�<��=	�;^D���&=S��<&�
�1�Ӽ4넼" =�ZJ��F����=��;��6�� ߺ�����p��t�<[��<4?d��� ��:����<gQU=�S����Z�{�a�BY$�t����K���D��g;��(;�9�!�;v=�;��<J�s�JO�B��$啼]y��	�$q�w2�<H������<<7|=Ϗ= +=��=[�{�7�u2?�V8R���+��3k��Ѽ�*l��Xo;�m=�z��{)��()𼫗�<�Y�<�˻w�\<���<	��;���<o�=���;Kv =gf�buJ��a�t�F=������<󉻑;!����Y2��e3=��v=X�n=-��7��<V�< �� J?��g;/I��-=vIϻ�Y��M6�2�F<G�T=N'8=�];��.�1Љ�}�<�{��CL�h@ϼ<w{<В)��A�c���ubP;_��أ�[`��]<*'�<4��n�<
b^=��R=��B=_90<>߼��x<r��ד�:�-O���]�2��<d����<G /��)Ҽ�Z���(�������P���3_�<Įɼ������)��
n�����Z,��3��d��cl0=�k��ٝ<=��^�8�I=��<�^L=�S�<����s=��,=A�J�Dv=�,�=�[<��p�?�<���<���<�Jg���==�U=.�*��P�=2�M���W=	�o�)�i�
����=��q���<p�|<J�<��=�,"=��"��Q=��p,5�4l=��<�Q=��q�w�2�6�����=�[��<�,���(��C�<��=I"��E���D=:Z&����;T��:�4=���;�@��<�=\'��!a��Wq=,Ӽ}�=t.��F=<`=+�R�<��q���süXe��a���!ջ#�3<��=�KS=X�<��<��%<���:��O=�Um�S=S3���P�#{ʼ1�<�xb���;���c�W��]O=B�d='�	=��9<��=:���/HS<X�:-ͼ��6�^u�U "=��K����<✬�*f�*C=��x��ѓ�I����<����sor���U�#<�=^�@=!�)=8�E=��/<ӊ�<�'=�"�<t��9�l<�1�<V�M�-��r��3j�<��<7v��v�w_<���<�pD=�aJ�>>�x���?�<�û��P&x;�����ٷ�`-=�nü�8(�|��B��ɻi��=TmR������u;�3B����+����+��@�o=Ga9<�Y�<�=��Լ�1���a<cE��<F��{0���׺��8<���Xg�?<<�;��<�;�/�
==�<�|�<�O��/?��H��TA���z輄F0����;dT;���,�[=��
����=šM=�A!=�`�<�F�<ꗯ���9B׼BP�<K��<�%{:Ũh=�o��+m�B� ��!{= ���������:f;����S����j�����:����g�=:Q=�V
=�8�ZY<�G�=�Q<���<4(�;�[u�'�=�-=���<%�����<<��<bE��p�<�b�:ߩ���ݺ��=smI��*ռXT=C=Ҭ��|μ4n7�]����!��f=j�-=�)=f�<o.�����
=��G=���<]����g��R��"�<:���7�� ��<9=�žE=�;=��h=��B�N�I=���#�6=��c<����6��Ԡ�C�;@?=�H�d~%�X�<9�g<�Bż���:l�8=	�˼�Ir<��Y<�����@���?�!�x�=��<��3��~�<#<�?��_�:�=�{��oV��Y=LKQ=_$:%��<\s=�ZA�.IL���<�����<�=�4����<��*7=��Z;��<������m`��䫼o�)<�OZ���_;��<���<�uF��}���r<���9�=�c=��<�x ���7����s�w =-n:=��Ov�m����<�*<=C/ɼ<$�e�ռ)����	;�W <z�W<�eR��9�<|P�e�=Gh��u�;�>E���"��ֆ<��Ӽ���=�8"�<O����¼#�R�.Y+=��v�|���okL�Ѹ=zN��/溦��<�7���\��&�`�=�?u;�J����=��+�tXr=�Ʌ=3�==1�<]��;�*=@E&=~�1�L��;����j^H���"=����2#1=N=MlE�"x	=f��<�2�p'V=��d=l����W�X@�<�eg=�˼��)�<���<�<9��ڶ<�E��w7=]Ω�	xY=�=�"3<�ϧ<��/;�>��Bo��k6��Ȼ��(�ƃ�<B�=�(/��%!S<A���Dy��#�YWg=��<��S=���P?=�@=��<\3|<��<B��<*��;z�<��`��W�.E*��C$=P�=HF⻓`F���<�X=ߣ��<R,��Q{t:�u�,�I=��J=�Jq=q�t<ђ?=J�=i�k�T=�7p���<z��;�A�<J<�V=�kW�myW=�VM�rޓ<ȋ7=�$�:�J���B= s�=u[��Wy=:��#�W��tI���3=9�;^O=+��*��<��Z=�g�;���V1����<��s<eGL=;I(��Em��W�<;p/��(���6=�+=��T�;($={
1��F_���L=!���;=�褼��Լ��Z�+5���%�91=@lj��?�<�i���A�<�Fz�VM��M�<�-�?a^��?�;�ꪼ��=')��V%=d0�<��2=�},�0=�2�n&���=��g���Ku�ے#=�=	���E�<<�o�H[�<'�<լV=�-�?^��@\��Q�<��<�?�;#�(=kc���3=U=����l�����Ю&=�F=�|<�,��}b�89���|n<��Y<kY���&=?�����=��;�BI�;��i<�6����ӼvUպ�N>��'�<�$H=�'��*!=��M���H��8F=ז��_Ŕ����6[	=���G}:�Gڟ��f��wA�|{=b5/�l+�� �<��;:0=��<�
�<��=>A=��=����Za��tڼ�D�z`=�n8=9::�Y�<=�H=LU��K�!�L�D5~=��H�`D=�5[��u$r<m=?��<B&�<�p6=O��<�����'��<4f�<	�=�!�<`�$��#V=�1�ꢾ<��K�Q���4-���t�<�dT���_=�ȱ;��1=�`:��򱼌 �<�w�<��<=���c�A=�mC=3࿼qY}��檼�[��YN��T��%@=�TA��k��o),��@=k]G<�F�;$�Q<�="�^=�e����;��f��8=i�I�b��;��/���=��ѼD�|=m�1��� =f��;G�X=�6��c$<>�=f�Y=>�w<��*=��=�p<�Fq�~a�0� =6�<�Y�y]�Y�;/*=�o߼��+=�xb<����;w��)4ռ��<�
O=�n^��>���T�<�=�<<�-=�܀�׵����G�A���m=�49�����4���x=V<s=ЁZ=y�n+=��<��3U�<�`0�4�=L =a{�;�Cм��f�P�|��G=L�4=D�<�/��;��*��Ҁ|=����^���������<�P-=3���7��<���<��<�����#���`�b5���b;P��<�b=�����>����ޤU=!H�*��=�U<c��<Ę<^�s�P��<��t_�<�P=�=[<�IY=b�<�]=V�#�-[=�Q=".�<�5Ҽ���=��=�%@�**F��v� O=�+�b" =��_=��r�J��C~�)�:��V=�Mڼ�<#
ȼ���<��<�iQ��"#��?=ޙ�����=�U7�<�¼1hR�0���b-�b~�m��� ]�6A<N~=���;%��::s�<��=�H�9b/=���~t}�z���9�<��+;u�s=��=<Q\h=h�=h)�}�*=�+���09��!=I=�W��N]�<O&<�w����|���;�E ��%|<Y�\<P��n��<W�1�a/]��Z;(�=���=^u=I���⼨፻�Z�`��<Il~���M==1=�e�� ;N1����=��+���a<���<e���3�d�,�-<�v=��_����ռ|
*=���;�\a=k�<D�;
���o�X=�|=����U�<+�˼����=C�=�B=�&���;�VE=�6M=o\�d��<k��<�<��O���q��Q
�<H)7=V%���@=Bϻ��_�tA<S=�<G\@��d�;��ɼ�!`=�j��ռ}�����;���S��BY���O�"���߬]����:#po=����o;3:=c�D�?��r�1sI��W�2r<C�'=�Լ�(��!n<*�<)�t<�o�V$X���<]0�<����˲9=A�<A��/Z鼋MջL �<�NU���ٻ��	<j���q�<FO�W!A�1Z� %ּ	=�<��*=��=ll��/+<Wz=�b�\�':nj�<�KX=�Hw=��4�˘4��7�=s����Z����D=�^M=<!H�����=~Wd=�|����S2:�����'��l=4��<�ZB�Y=���F�<$�=�5��Y���7V=ޣ.�x�<4�\<��ܻ��=�5�<��d��x	� ��8��*敼���b�U=���;0ɭ<A��<K�3=����JW׻>r(�w =ġ#=��;{.��"�P��O�<��~=�0��	^=L`6�!�]��Pj�P�]�<d��^=H#<n�=h�����}%*���i<�q�;+�<��6=�t���v��ϫz=��8=(���R=2��=��<�r=���<�B������ ����n�=�k<�L=��<h�.�|L#���绽ك�Apc���;Ղ=5v=H@I=��/�P����:��s�@��"0	=[�3=a�v<�gͼz�
=C{�C���BH��k�j<��O����<EG8�iX�<�	"=GS�~�<��o=��O=�g'��H��y�c��G6��ck���8<��N;tn#�V��<5;-�n���A=+"�z\����<�<lNp��?<H�C��dS�^3��6B����Ŀ�u�;=����=�{W�f�H�>�k=
�X�!�ò������� ��4�������'�rf�\�h;�A�趢<K�ӻ�QB��O�9��<܅�;�`<��S<��ϼ���<j�0�:�-�<�7:=�F�<"t�<(?�<��%=_}Y=7�<�Uԗ�y��<NU�)�[����<:�~-��� <Ɩ��."H;�C =�g�<yM,<�`1� �;�t��;�@;z��_�<��<O1�:���<���������.F�S��if=G�='�
 =9�м�ȵ��ؼ"�= �<�4<=�#����=� {�q2'�,V=��]���{���J�,��;�N>=�~{=��"=�YD=��:�o���*<�%J�腫<�~�;3��<@��Et��N���<��><��k=R���6�X<�(=�R¼�}%�
]m=��R=M�ͼ�z�=_V0�/@�;mp�;����z�Ś[=��p��9s�ꐼicx�&_Z�6=n4��L=~�};�
=m4<i�Լ=s�i�X�a#~� M�;�0<h�~=s0м�0�>w�<�}�Z��=�9��X�<�6��oT�׼`=^9=�K���$<�!у����-�<���<�>�L�ۼ<	=
OH�K�B��|����
��u�����<�t�<&T���M�����Q��^$���l�_�7=�ȉ<��o��$='�(��#뼁g4���M��Kü�%�<ʡ=�o<�"�<W�@�:e{�=s��<"��<��;A�+�L���n)��+޼Ʃ�P�:����Ƈ��hR4=P���_=��U��v"�"~$=��Y<�м���<�~�<���K-�;к%<�,>=Dw��`�]<g�Ѽ�A6=�#м�L�<�	<�z]���9Jz��l=�VR=�i߼�7|��-�6�j=Vf�;�o���ټX�����{k��L@�<=6]�;6�
�I޻p
5=�Z�YqA�����W��6=�B$=��=�K0��r˺�$=ǧ!=�ݍ<�f��'j,�c=��"=���ZL
�o(j���߼)A���T�$S���j�ZL����2�Jfa=j�޼�J��{��_J.�齚���;L�<�� �m<WPz���<���k=��B��-��eYN<��6=Ă	=�S
=Ѐv=�Q=�y;��:w� ��
=���:PS;[�<���Q���M=ďj=�%= A;����]����o>
<��#���Y��5�<��j�
=�]=[Wd=�=B���,�2�f���<�̎������Aڼ誫��*��4m��ע|��=�q�����-3b=د�<�F�<z��:YT=x�@= �w�$�<� �a=�� Y<H�f���W�@7=�A2��4=���<{4�;���<}���mz=�҈=�v�PFS<����r�~<Jp�C:�<0�ѼVWW=s��%
=C���d���{=܏ռ�iw=���>=�D�`�C�Dm1����;T���k<�>_�q,B�]��<J_�x8X=��&=F=�"��s&�ܥ�����N3�A�G<�G*<7�¼Ԕ.��X�����:�wм�1��#��`��<g��<�F5<�C=�"<��9��A���N=."��`�<Ɍ-�dP=�����<�m��AO=}�	>�<�S3�<�1=ip=7�<��u<<(�<X@ݼ�ԼS+�3�.=f»k�>���u��eD�?�H<�8�P�����=�������)��S=�(��BC/<���p4|�����
�?� ��.I��#=���<���:��s��E����E=.�=��q��4�<��]���ۗl=�k$='�7�̻�A$=�;E=�J���<�.m=�^\=��=<�5�#��<@��<�b�<4B�;����^i<��<&9<�\=z?g=f�<p���A������J����<p�3��ӫ��aмv|=S��<��i��&�<0^{�p6J�H*<�Y�;o��o�!=�"���������;l �Im=���<� ����_=냉;����jn<��g=���<ݭ�<x�ߵ�<�+,<<�;d��;�c=��@=[��F|�<8�/�]fH�A�<��ﻟ��#�Ǽ���J>v���M�?=��5=2[�/��:n<�<�C����><:�R=xI<���<^��<��^=��a<ݷ��y=x�X�ڼ.+D<
�y�e�o���<�R����;�	��K�9;H<�?5���U�;VQ���['���{6�GT�B.=�`�:�1׹��=^>=�|7�����W&�]����=t+�<s�z���K=����r�=]%;(�P=/���uF
=�m=դM:�2Ѽ���<QwZ=�~�;��<�W ��8�<��7���e=o�Z��]`=e*м�X<O�+�������<Ҹ��#B��+�<���;���;D�N�4n��w�<u#"���)��)�<=�<��q�{��<'@=c�Q���R���&=��λ��|<����4ϼ �;��<�߱�S>���D=�N���;=I�<6.=CK@=�=mkm��Q��F���Gg�N<=POq=��;�=�ܼ�cW��S<@P=����(��Q�:��d�Ci=1+�}��9��%�@�>����;i�x=�P:�=�'���<b�^�<�:F��<%�d�_��T	=,=�k=�;�h�g�;�Cz<�@��U��<sz��0��	�$�%�!�i=k�7j��b^���L�<o�޼g=��_p����B�>�b=g�-�??)=�	=�o��/"�<�N�<��D<�{d=�7�<��>=�Ҽ��-����;2R=ƅ�<7b<�4�I�����O<TsP=l���)��<gu�wr=��ć=���x�=��޼z	�<�}|��
=Ֆ�<)�0=�� �L���+��<ġ��j��TV���E�4+S���c=�*{<�<G���8�Č"=B��<PH��@M�HV�e�J=��<�MR�fX�;�XB��G)���8��a�����f7<��A=�K�G�-=�E����M�oH2=H�<�8���={?�h����t����<�D=�x;�儹V�
=�+%=�a6=gQ=���;�w�}k���=⛑� �gh���h�A��<�"��f�<BU�U�	=���=]�;�n=`i|=i�<JP����<3q�}�ֻ�����X�a-I<J<�O�*=��==2U�<P<�8t�;�M=p���H����A=�#�w;=��,<��ا4=�{+=��=����C6y�����5�0��<��<��P��<�G<A�<r�A=�1b��©�7ׄ��I�qD���c3����c=-Y=�z�1=<T�� �<B�����&k<��Q�f�=ݘ)=!(�;C�<C�'=�s�[�I<��B=�e��{L�<�h=NY_�c���6&���U=#)U< �%<d������!=f�����Y=Fa/�,�|<+��2ǭ�5n��b	�<�"H=��<n�Ҽs��j�ڻ�m��%&=�v=��</�a�c[~:�p8��<f�}���;��h�-�<�x=��F�c��4�<� ޺���<f`=��=�d�<��'=@���$];)�;=DNC<�C<��L�/���2 [=|}�<�ta=/�;�=�;�<��l=9P=fV�o����˼İ:=�|=�a�;�J=�����z�+�i�_�{���4<<�;3��<��<�W=[Qϼ��g=�7����'�f;ռ�=J=�q=EY��H�z;�%�;Ց2=2U=m>	�_�M=�����pg=�X&�Q�L��|��F)<@"�n8��I���~����;6,Ǽ��
=+�^���L<��<�H=��I=�d+=�DҼ��C��J=�u�Jӧ:���;��;S����f$�Wp-��z�;U�=D9w�1lP=���<J7R=�c5����<�C8�^]�c�
��--�p-��C�k�7� =��U<��F����<Yh�<��<�OA=�U(�$�	=�o=�5��h��Z����e�P��8��AQ�
���kM�(-=��r=�)=��b=%��<�����P��3=�j���2=�/��iMe=7t�<:T�<�2=�R=�P�j@=�-=Jϼ���T=�$=�I�<�BN=��9feq=��%;)o�ᚌ:�y��v�������X�D>���9b鼖ۊ�Wz<����ء���8��h(��p�=M�Q=��=@'=*xR;��N<01R�#2�x��;Eg��� =�aY�+��1�|�+��bN<��<+�;>)"=E0����"d=&o;�p�<��!=v�ּ.�;��`=�7���1�<DƧ��i�g(���ɼ�1S��hb��K��e^=����Ac?=lba=Bfw<F��zw���-����\S��s2�<��<������u7�]�C=j�x���;��\Ѽ�<<_�%����<KRG<�D�e�t�B�p=�Z̼b���ˋg�����+?<�;��v�r���<X������*y���oʼ8�-=K���;�e=��F<��<�)�E���R��<��<&a��F7<�=ں�V�h	G���f��u�m��m���r�d{�<E�2=��<q�G;iM=������<9�<��D���1��<܈��� ��t=�R=�7�<�j�;�b7=+�E=�H=u�;=�C=<����� ����$�}��jr=�2r��=ܼ��;x4=��!|ͼ��a=�tp=��Y��W�<�<<��7=��9;�F��m�;ɉ#<����똻؄
�ͷ<	�=�_���U�4s��8�<݅�C�K=�B�<�Y�ΉO;{�w;�'I�1�Y<c/�<.b�<-�	�h��<%B=��N=�=JE������.� ��Z��$"C=�����;��D<��=���<�w�_��<
�F�3 ü�~<�X�<�2Q=J<�=�E=5�<�]<Y�f=�i��WT��8=�o=;lm<����;����<�$<WF6=�G=�0X��&=�ڮ�i�3���<���'=�Մ��8�<Y��U=��x;�^��s�Դ�<
�=������<2Ź���U=��,=ݏ���g=�b����s���|�Z=�����$=��<k�;���� �<T<�5��1d�����=��J�
T��h�y�0��b1��.+=l�4=h��<դi9�ol=�`P=��丅=�c�;> =���<�6����:�}<�������K�<�ˌ���
=�:��R�!���	=]�F��T��3�����<��n;�K�<��<�]="q���A<̰=`K�:�F�Tm=Y���;��=�����c����i�<e='+�S���6�<a���9�;�`-���t�'2F�#�<x�{=J�^����;=08=���:�A[���A=-�@����@n/=��?<$���v���~b�L%=�J�;��8<$����O�S�"=��@��A<�N��cһ�K���9=rګ<�~�<u��;��\=�h=�s���%��8_���C�f��~�<ހ	=d�5=:�.���F=!�#<2��<_�<��2�^�z�^�;=���<4�R=�S==��< K�.
��@=��n���t<��λ��{<������'=�x��j�ؼ{�����d�٧�<	�#=���qFP=˱\<*e���=���<Kz=�=���"�v^%=�Q��!ͼ��!���<�f<�� =^���L�<՛�=�K�<C֚���q��:�π�����v�;�ր�X$��5�<�48;`� <�~P=]�=l��9��'���ۨ:��<j��;U�{�{[��9:�J�<�gG=?�d��A,=�-�<�MӼ�k����(�qW)��S=��3��5�:#r.=��=��0=��ȼ��<����:wH0=��=03�<k�.=j�I<'6ܻ �=�ϒ:�{� �伷�U���B=
b�<祦8�	9��sӺ�;�=�E���3=s<9�"�
5�;x�;�g��]3���]=j������=�a�%�<a�8:�����F��n=��L����<3�=��h;�C;�	�:�<o�Ի��<��M����	=�]���=u�4=����M�<�"
=�]ļ+�[=�;ߜj=����7=�3�������:!�<D&����C��<��4��6��`_v��5<��p=`jݼ~	�X+�<��Q�Լi]{�T=.s.<�k��d�p<���6���,���G�۠�;�ʼ� �;"�ƼX��<�Mb�u�'��d��
��z�����3�v*-=��B��m<C��;��һKˈ<�ZZ���&=J2���q�v�z^���Sv����d-;&]=x,���e5��hn=��d���.9<e���X<�8�ə�;@'�=�+�<����'&�jռ� .=��\:wM<8¼as�<PI�΅���t����A���{�u�C�´�<��q�����c���=��<�p}��>�KZ��}zL����<�߹�Ѽ���{=��=�U �E�@<0�#��p<�a��߼<�P���R����=I�ļ�=~�&���?���=�}+=�����^=NG5���!=8$[=ZxK�B��v+Q=p�!=�nE���H= r=U+���<#\���>'���8�<�2=2$�=�M4�#X�<gQ�;�g=l|)=:d��=-�eQj=o4��9�<H��<Q��<ĖH��l:��_�W�F�3��h\=��=ғ+��'<��<`��=��7�z�=�-<��
=��V��� =t=	��<�<��v�h\<�����C�<BY=s�4�<�|�4&,�Lu�G⼙��<�Y�<{�W�c�=����j�<OIF��h���"=o�-<���(���X19=�@J=Q��i���gS9<���<��<�����KG�D�������ix������5=n��H�=򘖼#c�:�lH�Dj>�&��(_����cH{=�[<bp=_��]�=)�z�1�����=f�=�V1�O�=�G�N��['=�9A�%AU<����kü�4�������_�|�>�C���h�Թӌ4=ʵ"��~=��*=I�ƼV����)=jJD��+D�*�B��c
<�Cp�d�*=��J���<��=�u����<�>(�TK���ּ�'=q/�
݀<#(�e�Q�Ω��,<L�S�(d=�6
�41=范��9C=�=��\=㫔�.]��F+�����<0��txI�t�9�u��`�<�W��G�Ƽ�A<�+L �p�4��M�<z,�<�^;9	��p7c=V;���&=�� �����IN<�9��<�<���<��9�-��=Pu]<9�n=��D�f�;l���($=u{��
/�eB��D�:�v��%U�<�P�<���<M�@����gTj���Ǽ��l=�����m$=T������<���+�ļ}
.�x+B=���-u<e~N<�M�<#!)���*=Q k=Ә�<�=_��t�Ҽ���������%=���94<=mZ=��d�5�;����@��p3��$�;��a=�E����=�x<�$���o�<�v
<�bL�}.&��U=��X<_Z_<�a3�$
=|�>=�[W=\�;=k�=�����<$QZ=1���ͼ_��:�o�싽��M;bo=���w]��
�_=�k�:�f8�g��W�f�ܿR=���5��p�~D���p��K}3�\�<��k��6�;$���=J;/fH=��=}®<��<-��C��z�=����k��<��y�Na�<hF��� =��0��'p<Opu<l[v�^�="Zm�&弌n1�*����:@�Y�����@=�H=�͒��JU=M�^<�TԼL<y��;�!�<��<���r+[�Ts��|�7=��་�d=ȿ<3J=���:�?�<r���x�<��R�
���{�;��='=:�=ak,����<�1��hh�j6�<��?<_�'���=ا��{��:u�Ǽ��q=俠��F�ؚ#�f��;�G�<;c�V�:=3��:�k^=�*�CH	=�W/���<�����d��D�<k.D=I8��p�=p�ɼ���<(���-<'5=*o���GZ�C��|�_=�����X;=}�<C;=�1��3��m��!���O����D����<��ּt���Ǉ<��D=�(,=]�G=C�;�=mS<�3�K�j���R=�y=�>�;ѹK<�1=A�����G`{<
�#=�3�<8�2=�B=�ā=��4=4v?<v�G=׽ļ#�;=*J�D�;=c}�<�M�;:(#�]S��Z$˼����d(=М�<D�d���<�*1�Th�<�V<瓗��4C=�a
��GK;c���fl�<��T��x"�V� =��{=��<c���E�=�_*�n��<	%��U=�<�,xD�1�ټR#q=��u=/,=��=�8��su�^d=�:i<��;zt��lk=��:��r"��Z?<�����")��_��T��wB=�4����o�����;�yK=��J��[�Xɼ�|����<�v(=�y���O���T��?�;�B޼6��<"��<_�e��� ��V� ���ڂ�/��p��la�<�s�3�=\���8W>�D	��=�Iv���a�6QD�n�/<&a�<�ZF�q4l<�
���A<��H��Ř<�z<2ȼ��<��,=���;�=M@�����,\=�4<��K�����o&���
�v{�r! ��H5�����0�r�Ǥ�� �;86=	�=��=���i���-��O'����%�w�:�|0�5?%= �Ǽƛ�<�`�;e|���V�<�{ü�W=mt�;��:齼ǖV=&��;� G=�v�˻t��3�����<埽;�b =�nL=���+�����'�����;a�K���\=�=�탻��r�$<y�[=Ha=Uy�<t�/:fJڻ:5'=���r��%e<I��<<����ἶN���=�B=5@�<�f�;� =��i=�F=0Th�{9=G�+=���K�<-�y�nR<�;|�<\�Ӽ�=Ѹμxӻ-B/�����2�e�K=4"<�P�<)���<�X�9��;�����X=ڽ=��<���<Y?<mc<���<�l��`�y<b=;%e��<�K�<��x�9A�= =fL���S
=T�; �!����E��<(�V=��J�kF�<G<7`3�R������+2=@$�<�j�<��<^v���M_�-S@�I�	=ˢ��eY=��N��'<8�K���	=9�ֺ�r�=�3B���3=��!�(GM=�����<�e2=��0�e�˼el��Cc=CG=�Vm=�������=u@,<A�����\��Z����<�f^=R��z^���(V�Qi�s'�<� �<g��<��C�"Z��|m��ʖ�����9��:�#�1�G=�=1��=��Y�:���<~G:�4X���ػ&=3{�:i=d<�����`�C�3=�Z��g�o��4T����k����<���#�<��Ț<��V<؟��2�j8�pw�<WK�:�p�<Q�μ��$�R�\��E�;5�%���5��0��u�F=X׼2� ���u�|�L�ϺN�������.��{d=[�%=��=��̗n<}�a<}/{=W�<�[=T(�<�} =:7==ڀ0=���aK��I��T�<��;Fd���X���N=�{��[ � �5��������8��:=����+��C۫<i�"=O����������L�1=�@{=�X~;':y���<ܥ1��nY<����d��4��<G�1���;�� �uL=n=N��</�<��Ǽv�0=��'�?��뫼�3��3;=�1E=�wn<�/��"�:�lѼPS<��Ｌ�I���今�J=�W=�(�g~������d���<)(��Ƽ�Լ�6�;��<y�X=H61<S��2�8�d�\=�vy=[*T������8`<��ջͯ.�İ�:�E�=��i����;\��<�<w\�����<�;;<�Q=�M%=�����?߻�Bͼ��a�j�Ż3��;�ZL<�U=�k�S�{Ñ;q<���ڼJLG<_��<J��:�l:ɵ�<dN�<�K�W;���f<���;p�R<� :p�I�(�g=�S=\aA<�F$���;�vy=��������J=i ޼K�A�i�Լ�.���7<
�&<u�<]D=���<�}Z<����E=b?�!�=5b�<N�ü���9d<�<���_1�<�*���!=/P��}�;�v��ͦ/����"Q�3�e=��a�[j�:��l�A�R�<Vz8=�O{�ye�<���9 �>N+=�9�<N�*=-�*=��o���:��V=�a�<�<�=��yA�<� �<�Z6=À��,<)��<,`��$��<���t�;�ǃ=+U�;��뼚��p&�<ȴ�;BY6���l��+,����;�V�;n!�3o2=*?���Z��w;(Jb;%��<Ro=���;�e�j̺��+=��=���<1S=bȱ<M����/k��QL=���<�|���Hc���:����<	3Ҽ\.��F��<���<B
�<�5=(��;W��;V��K`d=��%=-1�<��f�{�<�j=����Q��5&�<��c��G�;�j���=z5����;�p/0=�*��Լ].A�I�Q���h<[C��n��������T6��:�< D��KN=��=��<7H<��D����Q�5=��]=O�I�2 k=����������<���I�˻ي�<*�;�?�<0��L��Tc=.
H��3�#Ӽ���<אZ=]n><3����6�<cD#�Ec�{dP<~�<���:���;+m��+=���:��3v��@&��@J<��<���<�K=|�<�<�&=��K�L���<g�i��r���
�<UL�A��^J=)��<oEV=X��� =)��<5�5=����K��C%��!�ڟ��RF���=�VG��V=�?�凅�.�N���4=���<L��<��u<e�a���T��k�D�w��`�� ��ׂ��l_����<�Y3�KC=.K�y<�K����W�&l�<	AS='"˹RR=�-�
�N<ɺ�U�G��%���$0�<�.�:��¼��?��Ū<ɼ&���݇�<�9G=x�K�j༓�ݼ!�d;�C��B���VP<�N��<���-�<��1�0��q9��Ul��*�M=ȟ6�H�L�J�;������\�8d���=��>1����<`�@���<C��<��ӄ��4l������7�f*J��78=L3d=�8=.�=S�H��<�S0��ĕ=�C*<>�#�P,�:�P(������<��p�Z{&<��=�Ҽ@#<��w���<!)��ز�V B;7�K��f=Ғ�<Ɠ=�ɼ�'�w�W=�/"�|M%�Z��<;�̼�9�l1#=t?=| 9=�T�u1Ի+μ�y���xs�18�EK���=�W��/�=���<gG=������żNB��l���RE�U�<�~<��=b�*��^�<
"��@,E�o������8�b;���<�L=��%=mBǼT���v!>=�}=ؕ�s>Ǽ�xڼ�'�<,���}=u��98�<���<6=�`=�} =N����+E�,@=፞<�OP=:��<ȓ�1�0�!�����-~<7�<߽=��2=@AP=caҼL�#=&dA<)�(=������:�|�f�ٻ�����tҼ,�\��h=����=�L�N��ж�o4�=�F{�����h`=�f;g���g
=�y=�d��˚^����#=rz?�β�<�E��W=�����;Zh��߰��s�<h�=�cV�<
a�<a�b=yb���=l��<#�<�M��<=��<�G?������z!=q$��W�=�򡻇b�=��<�}9T//��L�3�<�Ic���<-�)�O-D��C�<�c�<�G<7:��K�"���'�;41;r�+���k�-܎��a�f�<���<B�O=���<D��<�o�<�}�\o =��W=J�={��:�c='��o�=�[Z:;&T���}�u<�KY��m �6��<x*�	���jO=�(p=ǽJ�=f�4>=9x<tnO=|p�<�8���h�b�.�tf�;Z�j=���U�+=��Z=�0��]䁻=�;���%S�<��]�١�<�Z;F<�:��k�8#�v�F<mBK�W��<p�u���p��l�;��Z;�"��7�<'@�<nq<P��xau����:k�;:�E���:��4=Kx�iG=����ϩ<�os��5=�F���l=��=�4�<o��<3w=ݓ�<�l0<w�ƻ*�{��q=`�Z=j]����_���*�$AX<Ya�<����7(�͕���<�8l�CL�Xˮ��0Ӽ��=��:=��b�ߘu=�k}= 1����<��8�y���)=Vw�;���<��%<��=m�c<�<���<��m����8@Dr��@���¼���,�=N�<�M"=Fa� D@=��7=4L���="m2�
�i�"�==g���"�<��=�+һD_<=�I5�f-=2Ҽ��=ZR7����0ּ�_:����<�4=��<�=�o������Y�k��<f�5��6\�h��8��=2C���P]��U�� =�������"?=�Yy��}!<~M���f=��T��d����c=* �<��3E:�9z���6;�_�kT=��<��<󂪼�=S=��V��;=EBT='�)�a�C�Y���CVV<{��<�I1�E���?�~=�pC=��:=��-��7J;�����=-�N=����:"v��\�����VK�#�.<�O�<{�#����=�?�<=/孼�7#�<z��;I���B��u =��:�T��� �N�?=b�R<���<T4=�ڻ�z@�|�=�:��<�÷���=m%	�j�!�Y�����?����������<�L	�e�<U��<�j<��R=��<=�� =��1��	[="��tn=�M����W<�k��.|=��w=�7���^;���<4E�<9�=�����'�=Jg"={��;�+!=8>��v	=�o��ƙ<}*c;}��<֠�<_����=ǈx<=�<B*�š�=sD��=�ͻP�b��<-N&<rk��M�n�	=�;���<�~��-0�%@p;ӛ�<��3�����3l��=n5���<����"uy:k������-߼�Iż��s=2{,�C=-��6���C=;�V<��~��!�(���׼�k�;�^=��v�������;���<�6м7��X#=�V׼9��pu�O�<�<_=$���d�󭢼KEo=�M���=�Z��s=�/	��tb=��f���=���<k��\��Fe�+;�7&ػYF��k�'���];�W�ȫf=:
=�J=�M�� �<?��)�=&]=�;�)];x��[�==�_����<[���&=`N;*��ϖ���(�U�Y��eU���мo��<�W=��.<^v0�e�<UX=U۟����8R��Y9;�#��0_K�521�U* =p?=cT�Ϻ,=����r�=��8=�ư<Wb�<0��<��G�)�I�/<�@=����% ��6����<JY�<D�L=d�̻@�z�M�����t=�;<�o =IT�� ��<��Y��2�;NT�W�o=�jv��`A=���<R�8�,� <����=�;=?l��y=�S=��0��#T=*�;D�=����g&�	���3�ը;�a�2=Ƿ=OB�<t=Vĉ<��N=.2U=��=��)=:�k=��=�C�w�\<<=\�;�`>��W�;�� �}��y�2<G_��6� �'l�<ߏ:��e��f;�c��r$=�06=�a=B���jU�)UU�����s�1�E<���=X,=yC��OB�������_�<"ĺ;�,�݌�<;N���Mm�����'�K��n���ц%�n�'����M=N]��7�N=�q.���(�M��;�c=��;O�$=r
�;����1<||R=��<ݙ-�u,�i��<�����λT�`���Q�<L�Eߌ�d�f��L�<bh�/�i=�N=~�M`=��z���G�<E�b�3�b�(=�7Q�XЧ<Cai;@�m���U;R}r���d�i���$Em<&l<k(�<�#��D�e�$j��E<
�";$
=}n��x�=�!v��'��<ާ�<��G=��8#��R�۲+��D =��)<�@>��W�<��'=�=�<�i=�=]C��:����<E�_<�}��N�;�U�<C�[�1�=h�R<�Q�S)�<�N���ߚ=T"<'�˼��켰=\=p4=o�7;'���J�<A���X=��/�a]�=�t�0�]�J_w<��'�*7�<�p�q!��鍽V�6�&a��%=�;�/h"=�$N=�R[�fy�;��8=X�:J�=� ���8Q=l2L=�	;=�3E���<P�9̪X��<c�&><��<��_=��I�J+=���9��I=B�<4�Y�B�<=�S���!=���<Ph6��W�RtD=�G/=����Od��i?��-U<�j��i���m�<��
����<�9��zg=lxX�ƅ���< d_=�^�=��<����M=c��<+*��Z&��%��==�RK���
�؂=�&=���<?k�<N�N=�"�Wb�<��ͻmǼfn�<���<�j�<�E�<�p&��?	=V�7��2�Cu<�Gi�?�<Q��;�p<��$=#AR��M�<R�=�r.=�H��\f=$��A�<��w�ם��ʤ8�N�f-=-;�� ����e���h���*�;�������ը�zb���$�@�b��=�nt�z�R��{�������깼��
;��»F8�6�ʼ��<�xH��=c�,=RW$=��ƼwmR��U�	��<���]V<#DY<@=�KZ<�/&=��I�;�d=�ᵼ�����/.=Ǽ��R�Ѧ1=3x�L7�;��=��<��=��{O=`==����	�<�̂<��Y=�9��q_X<�ɽ<r��;E��<��<��h=�"�<N���L�,��L>=�N"��}��q/���.O�T����su=��߼��E=��A=�\�<icR<���B����<u.ʹ�oR=��;���;�EB<6{�I�<k�&��#<f��<�u�<r75�>�f���Q=l�1���	��Ɓ��
�vx��8=���qR�ۏ���Ŧ�z�2=�#��x�8=j�X����\.�<;��:w����Ғ�<�W��9���<aN!���=uw=T�������&�=��$���Q=�=�U=~3j<���(��<;qrp=a��?�; ��<��|�g=�&b=H��@�߾=ʳB=uz6=�H=ӭ*=����<R�;yq4<J���Z�O;�*<4�[������G��&�<y�&�b�*��u��iػO8g��p^��1�!�b��?�;3 e��k.�|�o�>��<W�<��5=�@߼t�j�d�<�T�<�`�����<jֶ�k�뼋�#��P�<�����*xɼ	}�?5<���E��(��<t�E�����%Z�Y�<�F=Q$���
<�3J=	J=���<�� ����P�^`�ũ�<��Q=�\<&�;<W���[)T=bxO=�� �����¤�]=���qh=Y�G=�=��Ӹk=$��<	�<��h=�
�e�9�ѨR���?��e$<m3����5p�:Kg��&��9�;��v=*೼��=�m��<ջ-����*��*�(=�>K���2[=�V��M=�7�<�G�"v�<�d�	O�!5M�wy�=��<Y=Q��O;`�=��O��6��Eӹ�Z��JX=��<�e���y�<�E���H�<?=�Oż��;=��;<H���(Q=X�<P�o=����W�<�q�mr���8��R�ǻaf=�g+=}�A=��Ǽ�(<�@6@=���<-�]�ʕ�eJM��^<�Ou<�����I�z=���śۼ;�����\=��X�g��� �"�	�}.<j�����B=pJ/=:T<5� =yGL=��׼�E=_���Y=�I=�Y��1=1� =o�X��B<�ü��=��=e�)=B�B=S�<ch���R=��<\e���_�;���<
�-��k�c	I=�Z1=.ļ0�i���<��ż�=O�H�_�h���U;�Ά=�Ɔ�}
�<DRJ�92��ig�=6*H���q;B��<��A=�F=�0Q����<�b���=;%��`ķ���G=u/6=�P<C�<�%	��D��=�e=SK�����FK������˅=qm�<�)���.=|a�:�<^Ag��zD�0@^���=@Ѱ<ℜ<Z�g<�놻lp��O�=��1=񀺉�+�� =%\E=Q b=�Ƽ\n
�L�d�Y�ӽ;�$Z�J�c=�h��J�Bn�<H�F��:5�1��;�<���<
�ys�<%߷�$�<��,��<�x�V�e�L�S=(�(��V<��\=fG<F�O<6�<����	�|yk��]�<!�
��ۼ�� ��En=�2#�U��WFԻao�<�C�<�5�����5;���|<��D�	�<���<dqy=7	��G< g�<����_ɻ)z<�t�<��C==h�d\�<���=_��Kt#��+�<X�<��)�#����р=�U�;zS��f<���i�;B��<�-q=��<	+��A\<4P=S�*=YA7=�NZ��3]=�i^=QqQ��t���;=���vJ=�6=1`�<�uƼb>�<��==�V�<����`�	�ͳ�;�k=	��<K�=�ᱼz�<̪"�<|h��aӻi�<M�d�̙�����a�"=2h�)i#�t p�q�<�γ� �(��v�;/n��� =��h=2(H:(/��`%�<`����;m荼�a��eU=Yϼ�Pм�x�<<*�"���`���<���<��7���"=u��0ļSf\�<���O�<3��<�	=��Z=��;3#
=,d=O��<�
~�⢯��L=�Q:����#��<h�@=?M:�U�<��i�f �<uF=�៹c��*@=�QQ=!�<�м������8�F��;4�!�l=�g��2=�4��+8=�D����Z<�-	���O=�����w�:`��<�C���yk<5��<r�+��׻�O=�(B� ��<[�t<3������`��(U<��
����<h����3��8`���WC�R	<@2̼�r漢�켤p�� 0��U���ɽü*q;�� `��h���T��<�_�<Y�_���=�f�� �$;�~*�x�d�R�B<�s!��������ͼ��<�/<%��4/ =:w��P��<ih��SN:�,���<���g<=)hڼ;�S��sV�$�������%@<�p^��_�<��{<cR=n��<�d=�ȯ<�G�;���_=J�<1�<=� �<�J�<4�<!����=Ż�T�H�����܊�<[
=+Vl�}�`<���<�$4�����*Ij���<�Yj�O����	��tA=#�H;Y���Q�;:���L�1=7 �<�����x��:���$�T�4c�<"�<�~(���	=i�L�4	�)�I�r�ƻ �<��=�;p�Q��<��0��ur�����킦<��g�HJ�t�"� $�<w�:���
=F�ܼI����F�0�<F�ϼi��.�μ"��%�Y�6�g����-��<��G��f:=Y:���!��=��=��=4�l�=Ao=����﫺:�W���0�\�9�*a<W��<�e :�����ƼS�ü�2><�:M=�8�f;y�k��=���<��<���=�T<��༈�R�K�@=�=�߼l���+-=g�<�y\=��D=2��<�k�<�a���V��ټ<�W<G4�x�7������<�/�<9cf��輗v=�wd=;).�Qv�,?�x�<��<"��t༎�`<��=�Vl����<�*=��I=�R�*<��o���:=�_=Ss=z�k��=�	=3-|=���a��;�����D=09��	;;��3;J�D0�</�H=��}=���z�8�,
�<ӯY=�J���X=�o=��M��K�,�R<�KC��M=�:~<�W�<�v�<��=�-\=<�(�7Y�'[W=��"=�D��ϑż荦��,���)����v;��q���l��M��<<8��2o=yE=VG�:�@a=��S=������<߯?��!=�d�<��<���G�4=�2�;V�k���<��R� =�dY���<x��<MR�<�y=�$�<�1<8(u��:=��B='�ӻ��C<�ۄ�G��t�����;�L�<ʦ*=f.��N=a�a=Ю����@=�e"���.;g�I;�f:�W�]��<ŹP=���<�V!��1/=#u�<��P;=/����q<T�q<��C�Ez�A\5<V�}�0t=�g�Ė�,���K=�s����#=z����u=]= @(��=�5��'����:oM�:��<~'�\'T<�r6<"
(��C<�{ػ׷��o�|�i=���%��Y�=3z ��=�7<0:B=q��<�!�;O�Ӽ[rݻ��w�L��;[�%� D�=&QV=����'=k�^=��]��60����\���`��<�6�QdE��&p=��)�#~�U
�<�t�<<�껕����O���9=˾�<����,=��@�R�T='�;���V=��<<��/���<�����J=4ڵ���<y*�V�)=��-=Xik<]>���3=2�<�X";��<��e�SI�<V�����;	#=&�;5v= |d�/ּ��;�M�<��&=kat<�h�������3��s(=(���L=���c,�M��<�u�;�4�<��C��4����<�Wl<s�;�����:7<=�����<�S��	p=��6��9=����<�pg�Sk=�U�h=R�4��(!�oQ<e�,�����yB=آ�����mC=Ͼ���;i�]��߼O~7<r=��:�_����Q��'�<�P=.�<+�f��X�<�Ͱ��PR=3��<��)�7=����Ut}���3=��F�e/��ѓ<��<�J��Ƹ���=0+�wy=&<\=n(9�J'�\�Q��u��aw��sG�sf<�[098�<���>�L��Z��Q�e0= �<f��<	�<*;[���<<dn�e�E����:�=��#;3N�<��$��A�;߷;�N�|k���5V<xN=�; �/�<O�<�NC=�
=m�C=�Z���op������o�e�H���ټ(@l=�B)<RJ�3P��>|�;3<A����;7H\�8�b�����u'����X����<=<�HL=fe��Lb=���<[,d<U=V��Uü| H=y�<�^l<4�<�=;�+=v�A=SŽ;�sA= �� }�:��;��$�5퇼�/�<N��)5��s!�<LN���,<�=O�]N4�����tS����</����F��N���O$=�_���Լּ#=|o4�:�J<��i=�7U��-��6*=�O��"=�����=�.���ټ�`=��4=E:��v �i2ȼ�����y}=g��<�Fk�<u�{w�WX��׏4��:� =߼�U��!_O��6=���;Ѱ�ԧ<�Z.=�=b�?=Z�,=*���߰�<h��<�Rw�e2�<ۘڻ����ż?um<�B<��O���d�I��<6#`��c��*=m�b���W�D���n]p��xʼǍ=�7��R��<�
=?y5�s#�u+=��<�\�:hy<v=�b��~&�n����4���*�5<��S=c�=dsu=u�=.��<��A=��<���OV��+"��=�<hV��y�YHn����C<^=�=�$���tE= �&=<��<20=�O3=ꘂ=�X=��r=���z~=��=-}3=	S1=x��NH���6�<�:�q�k;�v{����;�k��FG<1V=S�l=2-����<�鄼ƪ������м�dc�G<Y=4V���R�R�S<�2��z<��j|�<�R9�(CK9�����d4;#oۼ�L�DB=���M����j7=���<5����p�m�?�Ox���Gv��O=�*m=l�����@�A4=Fx�4�=�o;�S	=N;ڼOt�<�$b�w�b����=�!f��0=�!<�pּ�i=�=G�V< ^a=z��<7�=t�;��H%���U=X���x����\��Vq=�~Իqy�<�l	=b�*��d-=/�=��<�&���<��;��P��fD<�#=TNѻ�|�VK�x=�T���;$֡��`L�6�t=0�<�=	<�����ǜ��-��I���i";�0=]��;E��K��8�,�9e�=��=Lf~�z1�<���<PX�;�y����<2m&=�k~;Vҭ;��2������%��ܑ�<%�K���X=U5���z/���⼽,����ɻ�<�];%��=��<�x��d'=�X�� b&�z���%�����l5�0�A=� �q�=e%=���Y�ڼ.�=�˂�P~B<WK:�0=�ں;pR�<��R=�>g;�UM<9B:=;�.���=~�;�p�<���<C3�B�A<S���B�<2:��	\�R2����!Pe�M�ۼ�c=W��5�4�N=�;ӼLU=�=���<��<V5�����sh;���P�g��j�Z�{�=�)�<�#=�FR<��L=���<Q���''���a=��<뭵�X��<��;� ��}�n=��@=�篼RB)���ἴ��<]rb�H�=�|=��e=//g��R�;3`U=ݴ=�N~=`=Qun�!<��08=��)<������缄�D��{'; `=W�Ӽ��&<��j<�U���|���	=J=�*=��P=�Ｆ|���D��k9<�Mм9�����=;|�L<��)<Gm<(ݒ<u�<:���<�Tż������,�j�]=,�Y��ʼ������1=�=�c�! o�	D=B��<�V��y"��F�<��<A�f�e1����#=�F=��D�z3�<���XYf� �s���<���<�o�<�+_=�n���>����f�5�G�3�\A��M);��W��x{��G�c?�J�9�ۧ<M��O:�ՠ4=�3���`=�J�W!<��<=]�!���V= ⺼���;D��<��<�%=Z��HKE=�ކ��x��F|ż�@=b�H�6�[�k}��f6I�A�/<��<˵\����tM¼�_�=���GT�����ח<�8��9�<g�<��<��J:I<�^�if�<� ����-=��O��m}'=Y�<x1��n����d<(����� ��?�<9=�8�<��ʺ���<T~ü�7b=�/���4c��b�<���<X�<>�8��5*=�U<n�=�&����&]����<�/4�_���?�ן�;/[=���8üz�ڼSW�g,�m�$;f��+-G�S)��A`D�=/�=������=4���+M]��^C��i8��#d<T�3=��<5��
!2=wE�=&�a�.Mv��뢼��=V�˼�B�k_j=Tx;t|����n��<��:P"=#H�"	=Ckg=��<�>s�=s��A=]X������=�9Q��`�=��-��Q�<�Y8=�U���3����������<<H�;>��ʟj=��<�S�:m�A��]�d@ :C��<�<�Mֻ���YR'�5�*=9��<��<�ҼǱ��u݇<?��:=��<�y��6v=��$<���ɷ8�(�Z����?�#;�i�x����=�.��xh��=D+�Ύ�������;=;3=�-=��,�?��<�&�I�<������<���<�д<��k<����f�<N�<�t9��⁽'#`��Y¼Te.=h�ѻ�`�+@�<!��,�����@=�ʱ;2N�Z�<�)=�l=4�2�+Vü#�a���N<�7�'`=N�,<*�<��=N�.=u)=2�Z=����]�=WJ<��м�=�35,�P���.�O=��<BvS�����O=�dn�<k=�a<;Ն%��q�<�]r=+����S���< ��<&��(�=�� k=�$��z;�믅<���<�F����m8��d<Kç�����,��]=�D<�00��<ӻ�<)=��=���e=S��Dw?=��<�@��"=��8<9n$��cռ���<-[�E�/�5�	���<����,�G���&��<��=�ZJ����=z������b=��~=p^��"+�y�<���6����"���<I='����=���<������X=}���޼�xμ$��Z�J��y�9�h�2L<nZ=��=�~Q<#����1=�CD�Z8(��� =>���$?�IjR=Y����0�;]/�}7躣*�`�������4�mc=��#=w5�;�*��׻Hs\=�wy�q�̼��M�5��@�G=�������<��F��&u=��G#��
ͼf������;��;&�����D+<r:<r;A��=/hI���<�S=-PG���<�U�<F?�E�μ���9�o�=�=�����黼� ��m����<�d�<� x�A�=��H=�RF�u�s:C� ���Լ���<�a5��1�<�	����/��d�;)���R�=�V4��=�sA���6�����`�<=�d;ei��|⼽#���)|���<R�R�9J��<���ļ�����j=~����D=���7�e;o�q=���<�Gk�;�<���<�=<E1�<A_w��tl�Y�9�4=�ڎ<s�*�h�ٻY�ӻo]=�8��Ĉ=S�:���<m~�����<CE��[=���M=(��<C|� Z<�Ǝ<=���n';��=.��<T� ��)��\�=��3��<.��N�j91���7���F9ا=�?�Ј	=�ѻ���~<��ɼ��M=���<�����P=��7�<�^7�oXL=3�0=�:}=�T���`=��0��f*=Pb�<��5�_a���a�T+߼8|��z��^$Ǽ�+ =�����ɼ�E��%L=�hż#K.�{o���i<�W�i���<"���o伪�<�0���e=m�K=��:J#��4�K��O�<B/k���$�
�jb<^P�<pFY=����k�u�V��f\=z����nd�S=�@=��ͼ�,
=<?G�P�m=�U�<���t=�}l�;��K)=~�<m?m��ƅ<^wA<��>�r��;2��=
�!�6�w��ԭ�\=�� =3м����:�&��]7�)�.=�%��xe�Yr�<���<��߼y2�<Bm��N�,.,=���A�(�d)�<�*=p.2��R�ț����<i�&��#��=6=b��&=f��HE,=��W=�q�<�p]8���;��=��˼�B�au=\�D=�p��!=ǥ#��Cl=ٌ<��+�<}��;Iq�<֬=`�5�A�(=���<h�M��V =��-=$o��
YL�wz����\<7#]=Z��;�u.=��=�aQ=�ig�<aS�C��<�3�:s?�<$�!=��r��|�<�c�<�n;2�J���=��&���m=?L���3����;�^��T���"���T�s����J=�ӼË�:��< �;a� �sÝ��幼 \ӻ ��#z-=�.#�/�`=�6%<�% <��M=�ѻ���=��L���#���
�-{O��
k��V�<]���H
�󴆻dw�=y���8;�k4=5N3<�/�U�6;})��o,<�F=��[=ѻ$���b�&}E���1=l�,�����Ǖ����J�����^P=\ $�_�<���,����ܺ\m=&J4�P5$��Zx���R��y�<L=�t~=�����>F�ت༤=Ҍ-=���<]��<�Qi��<��:=w[<�=��_�0=Ӊ��FU<�3�m�S��剽�d��o=�`@���<Y3�=G7�!�<�帼8H����~=���"Ӑ�K�~=����0�<p]�<����=�;����=�)�< �G�H������=JX@���ϻ+�=�I0=�:I=HZ�<(rg��w����=�v_���9@K�<LDf=a�d<����<C=-�c=��/<�w�A�y��GX=�m�<R�`�OJ���<�$:^�{<�u=���<,lc�R���g�<�_�=�=�|���$;-bc��d-���:7����<5=ϓ<!�:x#��{=�}�<���##2����< &6;a� ��<�84;a==��v;*�@=��M=�J
�+d�<���O�=w/=>8W=�)�<�/;<^V`��H`�i�ؼ�f=��N��v��m=-'=\�<�X_=>�C= ������=4�<=���<O�
�[�;=.��⫼}b=	������!��;ף�<�mR�]:9=�"��|vW=���,����<���D}�<��p:�ń�k@��,$=?^�����K=�1�w���=�ޡ:<������X�=}G9=�tf���Ѽ�~:��D�izl;���<(�x<N��<H�<�F�_�P<����P��=��/=�?�7*d=�P���^=E=�:?��<��<3ı����;G�Z<��;�<n��M�<�'<��-���>= ^���,=м=�a<�]��;ȼeV��ȔԺy�<b�4<Z���s	=�yQ=n�<{<[%�E�)=DA=A(���ǂ��[3���=a�==?9��μ�拼��'=%�;�[w��I�6����D=H,5=Sh�<'Ѽb �ˌ=�?5=���;Av���&-���=@'�<�L�<p\�<:^�<�q�j=ǹ����<?%=]N
=�1��:E=�#=�������<���=/�
<�#H<��<��P=&�Z�̦��M��G5�
�񼾿�9=����,;��<<_�0=�k==6��Kg���ＬD��-<�%��o_=�	Q=o)�<��<��"=�Ż<�X=�I=j�=-�<te@�N��<���:��<ҲE=��= %
�k �{�A��tU=X5�<�[�<Hu=7�a���?=Hi��Aw=}|8=6�����&=����d��wڶ���,=����K�<�$Y=C�¼^�=^���"ֱ;#���J���W����/os�����XJ�:ܗ=u�<����D��,��qg�<ۏ�W#I�c�"=TM<�}�����<��;/��<%n<���;w���I�<��\=��=7n�;-м��u�,x���m/=����B��Bm�l��<5��;5=����<�:�<����#�3`�~�+��<@O0=�� =�;���<�� ={�=ye�;�х�}�h��pa�%�&�Dߔ<�$
�zž���;��$�An=DB=8�<<=}��<Q�P=j�!<�E=�k#<y�8='}�<G̨<w�@�������<��<�[+����;5���D�<�}�;��=���!<7�`�'c�<H��S|��X0��叽�Ӽ�o�}dؼ؃�<���;|z�a�켔�a=h�����9!���C���(=8��<Y_[<O=��^:3�P�p4���']<J�"=Τ�;�g�=
�<�9`=�E=@E�=:�F=�}b�z-=����~û5�9�`'�7h��J�;�L����_�(#5<.������<�<��D<.�<�	h<s��<E�<��Ⱥ\����~���G��s����<h�U<j�u=;�=���<� ��j��8=�b�s����=�82��C=��=�@^�>��_FI=���<<dX=�i�/��<�S׼���X`^�e~`�4�����y����<�#<9l��Y�n=��3�5w=)?�=�4�>>=�5��s�!�Ӻ�'7��j�HS�<�,�d|Z�J��<]���)t��:�У2=og�<>b;�?��T�,<�G��&� ��������I=T19=q����#�:7/=GDͻ��3���H;|<[=ж8=k��<B���J�;���`��<$Չ=��1���=�#K<�j���}�<}L=�,=`��;��t=.�C<p ��}��Aт�c�;�2�I	��:����*=�Xv<�qf=�Ș��x:�x����G�]���]L�<N1&��;��s�B�@<��(=]n<;:J<-f+�[�;eE�}� =�ª;�L����Am��x�=?���6�V<~0'��+�<&�b��g=vk����%�c�<q'9=�8��bļU�c=�D����<E�绻��<]�c<��X<$Q�ə�!�,;~ w<��y��U	����<��=�#%���,�p�<7Zj;�)=��=�X��vIm=2��q�M�\�Z=�8�<O_��V�<m���/9=��:����=UJk=H�;��w=�k�Sm��T���A/��}�<����TAN�&���E���?���<�c�<�%�<*��*�=p�c�c-)��<¿��L�;Ok$��H@<�^��ب��+=�2<�F�<ᚏ<���<��=/C���=���<O�<�H�<1h�;z��;ͽ�~-�;�0t��M5=�f@��}�_��<M	=q�j�7x�;~�O��*Ӭ;��-��+ݼ��%=��U<��6<�N����8� �=�l�;C2ʼ�����1��%+; +,�/��<+�'=&a/<��2<�b�:3�O=!��J�Z=��,<P�)=�=q<�< *�<�"��L�=�z=�"8�+N����b�;��E��>h<ڜ�W�='�H<���<�:���(��Y{�|=|%+<���<�>s�XU0��9�/�4��7<<�����<���k��<�<N
���c��M=!=2��.x��d�ܼ�s��k�;$�;`�<��0DA���<�Js�yb:�10�k�=�H
�	T"�7�!�
4���;�I�?-=pf;n��CZ��h�<>�%�e0�<�U ��ݼG��<#Xa�%.�<cŖ�
A�g;~ܼ�!�<��=���Уټ�u�D?-<M�5�>�(�h��~1=s�==x����<�<^ ��fA�I�H=^y�:
/�;@��<�%<��;=Ḱ��-Y��Ĝ<��a�m��:�:<��H�'l]=�5�<4=�o�x����Eڼ���%μ C;���=Y�:<�{=��<vz<�h����=L����W��jq�3麾�<��祼WA?�h�9=P6=�w���6����Xt<���Hz?�io;�=��<]�(��i@=T߾�U��ĸ�.��=/�'=Ϡh<g������<�w;H��<��<od=m����Bκhnܼ^%�<��Ҽ#�<v��	�w<�nJ���g���;��4o=�S<|�<�#����Q5�ɕ@;�GH<��W�w�μ�A�<�d<�j5<��<rFW���{�{T ����;�+=<�g=�&>�w2@��c�<\-=�'�<1��%�s��<��'��>V��R���s=�6<mQ��P����<�W�<�n	�q��)�V=V񰼕A���1��
���{�kP^���<�\�<į��j��9=�%=K�V<�z=<N�9���m<�kK���T����<�:-�!#=uB<��Z #�F�w������<��rK��ڡ�j6ļ�!K<0�7��ȷ�p-8��g2���=dOO<͵���I��ȡ:fRu���6���3=#��yi¼�z����)�0=UY��1�= 9�;c�Q���"=\�B���j���1�C+�<� =��m=�¥���R<��<��E�<���<�!���wn�!�=g�;�N7=T_d�J�1=<~s;n��׃<1{7<�Z�<ں��g��<�1=�X��Ƽ�,1<H�==�|M��g���#;=��=+.=�̇=[�"<"�}<�؊���<S���b=��<-#=����(^����<>{@=5�s�ןk��}��{<�g��:�ɮ���=c��`��F�-�JO��<�ik�<rG�;�A�<~2t�������к$�ո�
�X�#~�=���<zb��<�]B=�@���򴼥��<� =��;��5=���<'vK<~=���V֪���;v
s�A��6s=f9��N"=�&�.��<ů���z�܎"=��)�[�s}E=��-=��<P�:��=4%�FM��������;��ܼQ���#�<�!="X=�ɹ̛M=N7�<=~U���ؼU6��
�9�4;==�����N
<�`�;l.�3�%<�-B=��"=}��4�f���l=���1 =���<���#�=�<=�T�<�-����#��ǐ<�P��w���żZn0=Y5+���<ֵ��;=�3ϼm��<X�=�ռy�=:�����&=8�ǻ�hR�G�μS���\�~=A5�=x��;q��R3<r��b=��ϼ��2�Ob:<���i=����<���<5�<��i;�}�<'B��<�z��<��W=�J�7G<��h:l51���6= _.=�!=���=��;�/=��n<�EP�����k7��w��=�|�<~B�<$=8=�hƼ�,޼��H=F�мMP�];/�,�;�=�;ͩ���녻bl��q>�<��F�E��<�#l�h���ʜ=e
����;'�Ǽ�ʼ>�������j�X=�޼�N=
�<��P=�V�<"���&?<��A==�C�f!G=-:=C�=g���g�<Q]=S@	<~;1�#t��!�,=P�a�˘e=c�7�`K�;�-��\R= o�<w?z=�01<�LM=���ZA�ߢ��"=�B�;bA�=�� �8A<�<�-����<�Vd=&��;%�<�y�<φϻ�C(��=��&�ڜ������M��<& �����"�#=ut�<1^J=���K4�<���<<��<D����i=��g��D�<�|k���=�Wb=θ�;�F=##8=��R=��.�-���`8/��k�<�+_<#��<AO�<}��7�L���B�Y3Z=Z�<�2Q=8z�h�7=�_��5=~�<�F�=f���j'y��#�������V<`�<���q��<!�d=5�伉�V����f���E=WƼ��<�v=;M�2�;�B����<�奼V�X��1M�G誼I�h��l'<�	�<��=!�����+=ʥ�<��[<���<S7������[]��
��v�=��^=8�<R�=
 �<�F1�u��<ClN=�'�����tCs<�_<Io(��f=�xE�'���=~��<>޼�_<�Ɏ���9���<��<�O���<�-��k%����<��/=8'x����;���>�^=�?Լ�˼������ʼ�J��ϼ�K�<W�j���7=�/�<�dA�o�I='�=����#���к+��$���	�g�S=7�*�����G"=�P<�;�<���늼�6�a;1�=��X�wnA=70<ܸ0<!^��%�>�e�;�O�(�)�;��n�R=.Dt=���ipU=���d�<BS%��+,=<�=��7=�A=mH�.5<�䤼��+�m�r��{���<��<�/���1��\"<VO�<�
����<�@;%��;�R��f��6 =1��<�U�E�<�d���l��	�=ћC���/�0�q=����UF=?�J=�լ��� ���༵�#;�9F=	卼����k��?�/;���.�W.��ͧJ�9����K�?=�3����<ڻ�I|&���M�;��z= �D���p<��;<�O�<H"\<<���~��Eռ#�;�'`�	�{��v2<1��<Ǆ�;���t�h9�Q�Ō��_�j	ͼ����<*K�<������QU��؜?�k�;7�';���<ix=�\G=&R=x_;R=U�t<���<4d׼S�»��J=��z:���<S�����m<��l=BY��emM<�=܍�;�-=��U=��q=�gY�Et���<�I=��J=�<6�g+���'<j6޼�4#;O!�았��fD=�
=?�X��|�<Zm<FrŻ�h��w=�Y�;�
��JP=^�'����<��
�ɢ�<?!������=��,�e�7=M�����(]r�>�S�_�»۞>=��^=AM=X,+�qm����0=��-<�]=���etE;*N�=Z"�<S�w�izm�sd��b� � _b��/�H^+=���<���<d��:p ^=46�(�=��d=w��\�<����L<�ɺ�Cٺ61&<aI;=U�[=8A=[?J�ۿ"=��ǿ�<�����{�<�<~�Ƽ��9=DJt��G=�^�<�e����<\�żh\��b����օ<ǣ��L�Z=$�+�) ��@J+=�|i<ݣ5��y=R�O��b�<��	=.�
��<q1��?�<�뤼p=��(���F�b���k�h=1h�;À!��rK�aq}���<����0�[�<�y�<���
�� h�<7�"�j�|<�sL;W{6=)��3X�<��M=J=��^��Q���	;�A�<�H=�K<��=��ļ�5:=�\=�p��Jf��$���!`�GeT�o=拁���(����Y�b=w_ �5��<d�.����=�t=�1=�n�<��=��0��<@�e��r=h�˻rw�<MX�=O;L<�ma��_�j]�=��=/!���d <�^�<�3��ǆ�c=[�����;1ȼ"��<�|k�B!:=����\��v/�0Z=
,�<����&=��;��Z�}0 �p��*-�<��鼔�?=��<�>��0_=�M*���B=eӼo�
���:�u�I���o�ѻ=?���n�K�`G=��`=��<$d�<+�.=4L@�׉j;��k=�zI=��=�>���d(�̟�U�1��ٴ�u�<��_<�M�W �<�I�<R�u�4��#���$�	�˼�R�����oT�$,8<��==��*��F=M��:��=�=��=�˴<E]=f�M��Ek=B9�;r���=k�b��)&=�=���=��3��;��<��Z�gNV�1���%|<�4o<��N���=�a��<���<�I��.�m<=�nD=�'`=���	8<��o�=�=.��0M�9��<$��;��N=�o�=ZQ=`�=�Eȼ8;=�g�0��<�pR=�C=��<
��,R<7��=@�)=-F�<�\Y=c6.=`�;��.���O�]hټ�Yu�f/�<�84=!t��T��n�=���<��E:WE�vN�{Ζ�uz=�_���|<ݶ��I���_=F�����j=�3<<�v_�/=��[=�_�<�x���{:-�Ѽ��l�fD)=�=�C={�t<�ļ�__=KT	8w�f�6�*�j��XR��7	=^Vr���;+��u'�<É�	O�����~=!�g=ҙF��^N�K��:��=�C%<h5[=,ؼur��
<�_��G�<+�7�)��`H�<M/�;�̵<[��;�'"��;=֑缼}T=ܳ��5��j<�`u;����	���! ���N=�V9=��t=K�<�)�<1H(<��=����:����z�i���r<i�M:�a�;�L�<P�<�� � p��.d=7�#�4��q��<y)0=?� <I��#|�E�X=��;�h=�<<5Q&�h�<����� ��;���g��u=����-�:ee���H�IQx�>H�<Ĕ'�(��<^3=�H<�i�EO��:<f5��ٷ<�<��?q�<��<N9�=�=��y;�G<�f=<���<��="{��4�^�h� o]�['�;��<����tI��X��BZ =���<������=$N_�ؐ�z��?�i<U?=�L'��6��r"<8�E��I=)��;��M=|�s<��f�(p��(�� �(@�r����X��/=\�ͼ��=��]��}]�B��=�F=��=I�<eɼ>{K��Dt��}�<q��]e=y�T�I{�E-=	i�<T5��u(=sꇹ/�;u�)��[g=F�E�cռ���<�����N�nz�<7<��m�#��Io�sk��'=��Ѷm���(��Hn�.�K=;�~<��l�Ґ?�ⷌ�3_��
�R��<�=y��`�{=Ĩ�;�� =K I��SK=��E=�F_<��d=���5 T�l��P*�<����I=��9<y�=J=	g�����<{���5�M<�B=��<�0��p�:@�;�5;=3Q��b ��s�;Z�R)���e�9$<�v=�ܼ
]*=�ق�v.��b;������;�d��l�S�+:C=�� ��w�Rㅼ���e�'��!��!rd=,!����>��}��]	=lp�<1'��J�+�J<����7<��c=t�����g86=� �j���O:�����<»f=�,��;�<=c�=a[�^�7�곥<+���=Yb���H�<�{=��A;��F��#��='�̍\�si=i�X=��{;�n�e�=<qW�<";v��c;�Qh��;���<�t;<v�=�/��#��qVN�͐^=�vq=�=1	�<��=;=Xμk�#� 3J�)
;��,���=H����d�O��<��+�0G���Or=.J'��v=y�:;SI��4�<�����,<��<6_:��"�<@��<*���k�=�<��;�<LV��z�.=��
=��s<�&5=���<�ک<*��q����!�<�����<#1;cH=��'��	��b-��J�=��$���N���U=
���j<��4;�"���4/�g�5=�æ��Y�=�(��)<F��<��w=s�[=�K<u�k=���<i�#���o��=��p=8'=T�y;��<�t����һ���<v=-=��>�>ʼ� <!�<�<���<�$���:Q�=f==�낻��<��D<�4=Oʂ�� ��N�<2�`�A�4�Pc=Gf����	;�F<�8ٻ Gؼk�<Q�C==��;��<=�pk���,�b��;tr�<������=˲�C>��;3<�����</+�����<rL��7�7��
�<
��s�Ƃ�<���0 =�U(��$<%�-�٢�<S1z=��X=���.�<)��� �<$_g=bQ1��J�������̼��=-��=���t=a�}=z�<ͼ�x�1�:v�VmL���(=�Y/���L<�=���<zY$�����;1=���X�ܼ4�:�&f�<���cҼES���b�<���� =�Z <m$���s=�yV�3̻Ko�<5�;��<���Z����缂�P�S��;=;�<.M�<�1=���3�����O��^D=Kva=!f���=w@�<�	2=�.`<��<<����T=��6�}d�<�S���*�;j�7�����n� ���f�L�̼Yj.:��y=�+I=��<�E���Ђ<��;�I�<SM�y:[�<��4��Y�z�=�V=���v���#R�}�=�)Ҽ�
��h=}0D��<<���;!(=ya����L�Rxu��!<��:.ݽ��>�<���<Y�<H�1�<��<)[�<L/���k=�^~��n�����;M���:�+B==�=�D-=��T���˼_p��O�%�{<�٩�x�=B�ϖC��@����ܻMA����4��;�=��=��;�o1=�Bn=eW���ټ��ļX�	��jUg����<����<:i=4��;������8��b���ͼ��0=���7;���g<N
=G���H�,*q�WѼ2pt�ڤX�jZh=3�<Nü�45=�}K=�>�<K�<��+#=�$=�=F���7�P<(�<���<ϯ<��(�����}��<�~�w{;�bT=�=7��<QE�;)��<�+0=31'���=�X���s��	i<<�H���V<ֶ[=�ܬ�j�_�W	d��O=AE��u��! =�����f@<�Y�ڋ=ɾ=a�{�}B=��J�����5N=%,&�ul��Q^�9�N�����.��<G�&=G�<��<I���S+=��<=�B:�w���-=;���=�i=Gf@=��c���<�_<=Pۋ=^�=U�<�1;�<���<�$g;�2%;LݺL�6�@�D<BC�����<��Ἱ߼��C����<�y�B��5a�p����;s(�<AȖ=��4=�D�<���:A=��^�<�Q=�_�O���h=��I��d�;��<�����:,�-=y�w=�0=��7=)��4�I=��!=��y<�8o:���s��������":=3=�-����<����0�n6�<׳�<� J;�k���<3�"�`b4������<�}U��I�T�z��.ռ�I=M����-�<Ѽ�<��弤�N=P�'�ߞ%=Zd6���o=��=P
�;��;�Ľ�R�%<X�7�N���żē���<O�X��=��=-�����@3�g@��j#<o�]�V27=�7�� �9"�7�6˲��z����b=��O��y�~��@99��<Hx<�?��7��׀
=�����Y=���<pb�8�<� �pJ���#b�`;�^��<O�9��<n������<���h��;d���Gz9|��Tn=aW9��}�9�,8w<��=���<�<N�L<�-�B�Y��V����/E*�4n�z-=^6�<�u��ӎ�Y��<p�Š9�FД����<�-�W H�]�w����<��<k��{;=)�,�U���9=a��;'i�Q�B����+'=Wsn�C��Z�+��A!��`<䗂�C�Q��ނa=:�^=�Z%��eD�l�2=k�n�����=k����ؼ��'=AZ<=�L�� !=�f����=��?�*=;����8v=�J��`��<(CZ�S�
C��<uG=�y�<�O%�����Ҽm��;!�;Հ'�
fh���U=�=E���<���;!
=���<�{��iP5=�ꊽ�\U���8�<�e<Ep�H�Q;� =Т�<ws
�-�;�Qp���r=��	=j`�<n��<��<�_�2�(Մ�5�?�¼:��Iv<,�=��<�VQ�T��|�f��A�<���"���e�<��M<��R�o�_=i�B�B��<f>="_
��,j��3=�n=nV�<ԉ+=�m.=,�����Z��EL��N�=�,��B�<Ь���./=��;�zg�^�,=h���~�(�(�0��Ǆ��}��-4=���<�=��U=t�<
E�<�e=��)�E�7������t�:/ם�<�=<��W<KB	=C+��-"�*s<�$�bb�<�;�<ha��-%�q�H<�P=y�<j�H;�2���I�GC[=!Cd= �<R80�/ 4=�$<= ༼�0=
��;�u<
͗��]=+�����1�\=�H��;=<�L<Ϙ:�q�Pp=�yi�;�A*���.��E=P<��<���<���^�f=�=b��<!.<��<��=4G==�/==�w�i��!<M�/�
ɲ�Ps�<�#=./�/\�<À�
�<�㼴�P=��<!SM<Ah�Sർ���G$�;��������s�0���	=�&�5}�<��<@�3��g=`=.�9=�3��VڼNtR�>�$<����Fm=�Ȼ�=�
�R7=���(@��qO���]��׊f��B�<���<���<ăI���@�K�p��� ��:�^?G=��/=f��<�$N���G=�s(�u�M� G=~T=J�"=bC�����c�=��[�r*��A^;�����=��;�f�'=�a=X�<X�	=O��H>��;L������k=:
<�b��/�=�HV�)7���<}�M=on��ƭ�<	����<;�
�[Ө<aFY��=�2=�@D<�[ڼ��Ӽ�$�<��]�v^=H� =��<�8=�)=�Ȩ<�L+==.��
N%=g#=G�^=��#��E:ZWY=��}�mȮ��oP=P3=���<�z=��\=\/_;i�)=��V� 	=k��<�˃���<���<���<:��T=��?�d��<C7üe�]�B��<�g�<�n������l�D=Jx�<r�=pO�<T�%�Hrx��``��N2�&��<��.��	t���<��;P�v=��d��D:=�2=T.;c�%�th-<ؒz�b�һ� Ǽ�b!=	LN�6�����*<�r�<�-��{�m=�t7=�K�A� =�d���q<��:�==4�<У�;C�<ȽD�4�
<>�=�v㻭UܼEr�;����H�<�p�<?SG���;��7=�2�ȳ�;����F���#�9�����ڧ;��*���=�0��;K<�O6=A�d<x�=��I9w.�;U�v<���<��;m����%�<����G��E�\�'0ܻ}T�YOF=��o=��]9qCC=<����'X��0���O=ݢ��o��:��q�����*��U�,�L�<`�W:ӝ<"І<vȾ;,[A=}�B�M<��Ic����M� 1��/>=;a"=��9�)jV=�i�=g���z�<��6=HT�<p5��/h=���<��=��q=����U�#�7k2�u�<]�C=P|6<ؕQ;/�#���7=<�]�)|y=vN�<�.ƼǴ�Z��c=����2;
�<�d=jO=8�G=3��<�f񼫅Q=�?�M�(<�J^<��<0���(�q=��;`���>P���:;�9=���<�R$=3��<�I,�E�%�F,�A+���P������<{=���<Z�<N��I��<(��<���\<�떼Y�B�xE����L5����<$1��T��Mw�<���<�L�)k�<b�<�Z��,ü��r�Q#\�:\���5r=N�#= m����%����IrR��Q.��>=��:?��9�3";)[4= ��I�<�Y���)U<�@κ%H0�Ue�c=��<�5�<8�5;��A���.��@��<gF"=�����O�<��=��B=�,�<�>!=>G<��+��1a�I�9����t/��xj�^G<�jW<�H�-�|; �����8�A���ϟ�<�+=�:����/��Y9��jcS���;(Yϼ�8p� �a�p�Z<��K�)��<�q�>�;��=FK.=X�I�m<Rt�w�K� �=�߃�Ԇ�0jQ=}ud=���X�����<[�;�l=w�< ߻⣼�\r�!�=��,=���<���<�旼:�?� �1=���<���,�< �<��:�M�<�'�<��3=,Q�8� ����;�H�<�h��S>=�Q,���f=�5�#�8�����X;[>��@��w�;���=c�c=�uL<1�<�̙<��Ӽ���<�b滐�=D�9�D�<���D*;�1O;�������+�?=4@=n��9P5��Ci=	��Z�ڼv�v��5�бQ�+�ּ�PU=���<>��<�W�8t����3=_�5�D�+�H�R=�\=ʲA=�w(=x7߻�K�;:q=w�B=ĳU=���<}Q¼��4��s�<f�<'��=<��<>���ͣB�[�J�rHA��Y=M3ȼ�f��;�3���<15;k��<}��j�}<�����Do���<F�a��E=��#<��6���ϼ�sY�D�;#���3g=BC=�� ���{�M&$�nX|����%~�N�?��MO=�0=��f=�Cm�9y=͢�<0oV=�:�<�jD=��<<�J]������?=��= ������v-<��<fK��n-=���;�L=��5�/�=0e,�'�%=�<k�X<��^=�a�<F�m���O<���<�����<>��<�Ժšo�V-���6=��q=�6��Na�<9���[S�**r=n��45�G�K���%<�d��o���^�[�K=�yq��)7; �q<5<�<٩$��T=��<��ȼE�i�-�<U�<n`���j�6���ƽW=�%=��y���|���ɼ�[q�R��NY)=�jV�Ď,�i-�RU#����kZ������ۼt�;<��W<Ŷ<Ak�#=U2<�/M��5���<�1�<%x}=�E;;����B�]�8=��<u|��}jC�����@��Y�:�m�<c==&M��\�s=�:M��<� ���M���2.;�6=�\ �ݯ3�i�R�����.�=��ռ��0=��0=� <�������&��:�-=9�i=�c�'���@��<���F&/��2�=?E�<�#���=�A=#:�VB�5+H=˓6��Ȏ���;��(=Ӏ9=�B:��L�B= ;�׻����<���I!�O�=y��;{5�<���s0�;�Vq�}���X�N<�^����]�ǼB*ͼr�[=�J�=�!�6��=|���2�K�
���	A<��&<����A>r<��<M�����㼢eJ�� �<�|���d����;�MT�_X<�H��c8��`G=ԡ=��f�2��<W���R�;�yQ*�w��<�Z�<��`�	xc��g�ز4=5��<� ؼ�����p�;�#���qt=	�<�t�f�2<(��β<F�-���X<��E=V���.ڼ�B��I	�� ؼ��<7�<5�>�/)<��SJ(=��̏�;�?��=�W
=�qX�7�s�i¼�E::�=w�F9Y��B��j<I0�<̲���և;�i�;��A��ii�g��<j���k2=ۂ��� =�o���)6��&b<��ɼ�6+���u=��K����M�Q=��мX�T=Fm��ʏ����<y����W=�Q�:s�$�=��2�F=�4��"=�=J�)=��C�(/r��V�<��^<`�m=!i�<"��<���<+&����;�W<鱙���-=��U�0gq;#
�(}�<��,=��G=A<�<��6����<����LJ=?:��T+;38=P�f=���<�CӼΛe=�=Z���a�)&=DT`=(H=�r;�����<���p��<���nԼ_�2����	�Z�<=��?=��<��u=.u]=w���K�_�i=%q9=]�<17<Ϙ���t���<�D�<�E3���Ǽ�����\=�+X��
�<�#M��r�< ��<�[=�!�6t_=F�I<1��<�Y@��2j�9n<���:�-�!=ѐS<�4v��[S=���;�?��#6='��<�sh��º���v=�U��0I<m<�<�oؼ/�ͼ��/=C��h=Q�=��;,��� ���>���<���s㭼�х<f��;R	;o�6�c�J�6m=���}�<�"=8�/�u-9=��a�Փ�;NE��ռ�[��C+�|�a<���<`�I9�<��[=��˼c��碼hW��-����;i��:I_d����I U<��=;�=���"�ؔE=��k<�4;��<� �,L�<<��"�_8�<�����]<�d��( �1��<A�ü��S����=��@=�!���r��ť<,�B�&=��&��}i<��T���~��T���T:����Jv�<GX9����<�;E��ż�7Ⱥ��neD=GQ�;D�ܺ�z���%=೻+ݠ�C�=��A�:�U�� @�P"���C��+k=�<Ä˼�
=�r;��e��Q�i�=\��j�8��yj<M��ft��
ҼP`U�>z�9�W�����!<S1=�;k='��"Tڼ��=SV�<�������J=�m�<v�����8�����]xX=���<�
<� =�[żn�=��<S���Ö���pt=^��ߒ��ݭ���q<��P� -=R5=�Zf�4�x=	n:�T��Ks<���<���<T��<7ao�x9��+U��d<�)�%���D|6���%�[W�!m�/T�<�z�I�>�\<ߙ��䘛<�rN���V��a��Oc=hP=A.��=�B[=���U�K<�O��t#�;�I�<	
I;���<,=��c������=�5��9ü��b��=�7��Fo=\����%��m{�k"w< ��<��X��+4�>���ĻU`7:8�=I����<����'`�<�a.���$��=l� <G���~�;D<�Χ�<Q�d�[%V��E���BX���_8zn�<Oi���j�<G�^��N�;�H=ז�n8L9��8<X�*=g+N��?�<G����<I6*��Ӛ<�F ���g�uA0=f��D��:�#���<JxT�$�&���Լ~��s6Q<�?���Tq�8Hz�ټ��=��,��˼�r�<�d(�8nD=�����=��o=���]ܼ�\+�3R�;�N��p>=�H��
I�eO=�k&<��ļ�q=�=�r�<C��=���:��<�
��1=� $=F��}��ǧ㼿B�<��=���Ũɼ�K��=�-X:p��1y?=֑8=/?���v<�
=w]=y�g<��A<�����;��>=2(}�A^ƼT�L��"�<A8r=���੡��[?=́�_���[��p><�&���%�)S��a���5=��=i�9=����+��1�9�$=0�P=�@K��l�<Hp��+�_�=5�R�{1����2I��Vq���:~=�[�n�(��=��<_ռ}�?=�+<;[ƞ�B�W=*m3=��=0Z=i"ܼ?d�;�=K6��	G����J�Zm3=�GA�&78��hH�΄B���x��
��~��"�\�d��X��[����3�/�[=�{ ���0=V+=<Y��<!�q=�F�
۰����<��y=��<��~�;�a=�nm�餝�S�<�c�; -<��T�6tJ����<֐���D<��a�#�.=������R=A��<��}L�<I�=�\=/��i�<��h=�>m<�D.;HX=��=��@=X1e=�t��KPf�"�<lU�'�\�Nh<�����᪙;oO�<���=H�����R�Y���,S<$6:���O=���<��Ҽ�����]��#��&G=�\!=���<Q��<���<��o=��T�v,2=��S=f|���<�@�����]�<����L=����TȪ;���<(@i��ن=��;��<dT-��'%����<.3���R;�P���b=2�������#=��;/�s=o<�Ɵ�<X��?�(<�i�����>�^�k��S�:�;�;�Y㼈��;���b��<��q�>T!=�%�m�D��s�-���怆=�Du=c�=z�2<��<� =�\5����<Ӄ<�*K�B�L<!$�]�='�P<��l��^�O�U=�-P<ki?<��f��Z��[�Z�#�=�3�VJռ�{
<�ɩ<ۄ�.�E���v<�Y�<,[��A=a�\�Dؿ���=W�6��=/=��g=�K=)��<d�w<�̖;%�ۺc�1�6�<�k�wZ<O0�lP�V�z��Q�.��<t ]=S��=PB�1~Z�b�F=�R��*<�:}���<č���M�y~�o|4��żۿ=�@M��R=�J����w���8=V�L=q����P=��;Tk�W)�<pJZ=������<v����7��-K��T7��<=4��<Z�T<�1�;��<Bf;69=<#�༤����0�D��;��\<��<W�'=/!@�N����A=�/�ջk౻yv�<*>4=yH	=�$Ӽ�b̻��-=_�G=����f+�n;���&���F��yм�1������O< �\��%�����><<P�=��%�g4 ����<H<=�p�<��n<Q��<���<��U<q�D�#mq��N�P'+=���y<��L��9� ��<d�}�C�4<V�!|O��yc=�n=r�+=<$�������=�HS�m�<[=�T=�LW<#�%=��~=s�<�j^��k5��~��m�<J^㻰Q"=L�<�0��Z�1=Ê>=��=!�.�-.!��TӼc�9���%}�p�C=�X�����=���<9��<��-<G�1���=�ѡ;fG=�0=��I<J���o]l��4+�h:R<c�X�R���0�#=5��<& 4<��D=H�U��p"=�H���c�<�T\=�V�&��� 5=3�9��������O�^�X�0\:��l�<��T=+�K�9�=�M�
b�D��b�/�,g���$�::{;���<�����|<�(+����A�<f0�<��}�-=t�W=�<p�H;mGz�˼1=��<��NǻId-���ؼR#=!��<��u�CL��2�4��T��֮ʼ%yZ��8!=�w=`������xV�!]��1^��oa����͖�<ۜ+=��={�1�:�@�Iu+��\j���	<���P�����{X8�d���=��t=E��=n�꼁�J<q�i��g<-3�<-�=�"V�&:;,&�;��{)��0z);ȼ
� =���<>�K=��Nm�<ƿ	=��_�W.=�(�� d��*�<��4<f����
߼��k���g��<z=<Ñ���Ƽ[ �;J1�����o$ջ�Z+=�	�S�F�� ��'<A���җO=|�<��3���>��'=$�<ˏE=�(l�:r�)L=Պ�����\=^��<�H���!=c�2=e�(�2W�<E�ȼa��<��.=�#`=Y����w�<W<= ��7$�ͫ=c���Wh�('�<�k@�&�&=�"�wN���M=�=R�<pN�;v�'=��<���<����|x=XJ=]w���G'�'E~=JWV=%)��*=%�� E1;̓;B@��	;B�(��.]=[u���q4��
=�߄��Z<8?�/��<a��<&�U�P
1<�>�?��<@�;=W�<=d�G�Q�<���dI=��=ns=�I�E�#:|=h�a���;�k:=b�Z�\��l�=����d��<���X�p�<!	Ѽԙ�;, b��J�<���<K�=<5�E��`�:��R����=�-�=i���Q��<o�\=��w;�r+=rJb��s3=W�L=�\	�\y�<6tH=ķ
���c����0=�I���v�]�2=U�;��<f
=��<��A�H�h<�l8<r�!=���;�%*=�|ü�� =-_̸��0:ǟ5��p)=<<�F�<?_M��=;��</(G=Ƚ��j�D�V�"���ѻ��<*����Q=t��<�,!��"�uCZ�#:�Ң�;������C�<�
���g|=�?=J�]=!�C=���8�==��8��IM�X�.�����'�YO<���<��/��l�;|�&�tgm=G$�<�V=�B=���<���<2<�V=G(P��s<%ޭ<��$� �=��l;[�d<��<�o�I������9�U�M����׼V�<��=�Tg�B7,�	���T�<�LB=����O�C<����,s�<�`�W�<L���G�M<z�=g�-����;�@=�&=�?�<��#�h=�N5=S2=Q��<�]=:�<)A�;�=��;,�7=4��<����}"��t�<�B'=�M�1�7�G���@�<�Y4=!h�=^�=U���/�����������[�]��m=�lC���
= �#<t�Ǽ�0�kV����<���KG=eD�LN�yz�;]�z<�N�<n��<�e=�y�<�?ػ�{���t��l=�0<��I<�x<=k=�eN�P�ϼ��=��I=<pz=�v=��b��	=(����	�<i9,�xR��,�&=��׼ǍH����===򳪼ǤH��.<����=��&;�&�=���<���<`�;;<<���sƻ�d��S?M=p�;Zt���-=�����<)����5@���p= ;�b��<�$J��l7�~���_��S<=��C�1�����|[d��63�Z�ûU��D�=�H޹�'+�*4<����-�)�1�A=�������/=+��<��T=ͧ�����oR�<_3�;S��<�;K:6��;��H�Mμ��ػP��=�6= L��O�:�!�;��<�P���?=+�k�q-����<r�=�?o="=����D$=oy:П,<���<�V���a=��¼b�{=��=֞ۼ�+>=�D����<��!�g-�<��<�d��'t+=6Gռ~��	��������[J�<C�*�;�M��d�����>�<q�����^=9��<�4�+]�4<2����;P��9ˮ<A�z�}�&��KJ��^f=�7F�j6���l��]	 =�9�<$V)��C=�v&=t�ȼ,�(�y ,=�b1=� ��<-��<Pѻ�|g�$-U= ˚�P�F�w�='�=�̖��eB=L�=��K;��/=卼����w�0=s��<Y>�=�B�u=��=%h=wg�;#*������!0=K;�XZ<��E�L�+�ɣ�3��<P|=�a=���)&ԼD��J�[<6�<{#]��S�G��<�3ȼ��6<D/�:mD4=V�����<f�=���<�ic�ȸ���-���<Z��=�a�<w�=�!5�#++�Ww漵Ƽ3;�-U߼����7�����9!=(��1��-�<�J�����O�;��Ѿ��1m=�G�<�Kq9(��G�%=z=�i�O� =�m�<Q@n=� =τV��>��x�)����<���;�J=��M;���P�<�y�;J���.�<= ;wX�<I8�<��;CZT=�}�Ὶ�x,�<�8=�ҥ�!Wx��^z=��= p�:Q�������A=J`��xx<���N�s����<�&�;��z<.�uy�<��Լk	��R]�7�ȼ�ؼ�W=>�J��t����5=�e^=�vQ�j��0m��,Z̼
#���O���d�*��:4�6=j�=�E}�~��8��B�c?=6�q���5��i0����< �:��[=�������=D=A=�F@���0�hN��8 ��5�<'��;��	��TT�ϟ-=ާ��K�<�;�ɸ=̗p;�^�<�Ĺ<�a�<�NN�g�<6�<�]2=�E|�7�<=�]=0j<��D=�/U��
��zq:<�vȼlb%=���=.�A�<�Q�c�:fH:��D=�#p=K��}b�<�����(;e7{=�~ܻ�eb<'�L��ŀ=�*B=�2��i<�����<=�<�	�<8�<	b!�r �ջ-=�Cr=,���@.���ݼ��Y=u�=��6/��2=�=�jz���)�x,�bl�� �]�j��<�H4��rf�@���r<�9���<�3m����<[�B�i�9��m&=ޟ=��:��<�������߼5;�A���4���<���:��<=&�}=P�<pjh=�j��=��N<3μ0�T=�����ü�p��(d=�;�̋��_<2[o=��=��=�/����<�J�<�qҼA�ϼ�m򼐠.=Q��8
Z=LG���(=z�/�r�o��=X��<��<U�l=/T�:}�*�#Yi�8eH:�T;��Q=���<|mɼ�@c=]�6=�����{=a�˼ c}<SI>�����s�<L���Ki=���	�p�ڻ�G���T;J�<�X�<�8A�-��K]�<�J=�:;F������<�<��]���=�>��H:=���<r���-�>=���;ZY�<�ڻ�q�<�'4�ͤr=n{�N������|�?=GY�<
�\�=aX����<U��;I�L�͹��B��oD=�
<q�<�"伉^�E@='��/���}�F�eo=˻P��=�X=���<�`���꯼����z=�G�<�F2�{h�l�s;���$��SlG���<��R;�W���ֹo1e=�ˊ��È��E�;��8��c���q�~�<�ԼbAy<��S=]V�+Y��:=d[W=
�C=4Ő��J8��9H�;[aA=�°�]�K=ʘ��Tg���T;a�S�̮;��<3B<�X�<_U=[����2�j�#=6я<ș޼�2 ������ռ\���G�<��;c�`�(�E������;5b=p��f)=󈠼�F<ԍ�<�xY<��I�0o�<� =�ZB<	Ia='�<����<wd'= x���xl=D�ۼ����_��<(.$=���;=W��)���宼��i�	L����;�b:=����+|<|�c�����H<>�C�)Pe��?=��b֩<Ifb�J��Y�����:�0$��Ԟ�U�	<��<$2�<󥯼=EB��2)���'=Qh=_��u�=9�X�~5[��㭼8��<P.x�E.�;&�I=�L9��V���3����%�b<Q=�gL��?����+�-�=����r^ ��j1��O��-��X-D=�y�y������25���m���9�F�=�;V��;�m�<�F ������
��F`<y��J�q�H������<>�B��<����)=ʥ�9"j�yؿ���@=z8O��PU=3g3��j���P=�C3=����Y�üH�<�s<�GY�۱-=�9�e=���<��|� �0� ~<|5�;��p�iE��eX=�����Ǽ�ᇼ�,�=Pٞ<��<?|�a8`��H<&�C=]Bi��;�<���f�m=H�*;��Y���W��w=����==uJ��U�����$=�u����G�� !<�À���=LW�2H=8b=��e�B@��v<\:ͼ_�ܼH�=���_=��z�7=`�@�_�L=aV�<6�ü�`!:�:=H�;��	��`=��<7U0=�Y�<�8 �YD�;�zм�A�<~�&���=���=�j���:t�<�T��@�<T�S<��;�j�t�n�=@�n�B�<E;�;_�=���I�}=l+�����V�F���`2K�VJF�}e�;v�p�>�m�;;�=���;��<њ}�1�<=�oļ�=��"�Z����;B =�u��X�}��t���ʼ��;�5=�H;'�7���E=1��Mἑ���)�<[&�;B�
=�?T=�4P�cR���Ƶ;Q����<ʁ�;%��;qD����<W[��< ^=]�&�O�ڼ�����~�����$$9��lͼ�)c�zG���񾼀Ri�@�=�.�<��ڻ��l=�@~���j��#�=���< V��v�
��J=�G<%�V=�#.�~��<ۤ�<5������=<,���+&=ы�<�=��b;�^�LGn�pN��\+�4`�E.V=�v�{�;BoǼC��U�F� 8�<�Hz��=D<0n�\;��S���X��:??M�N�q�,�O=�B=��6��s=�p=�G��CH���I�=�P=��S=�%� ˓�G?�=�w<
���6,=��4�m?��/� �]k+��{���+A�6h�ވ�b7=iYz=�)C=>��<�y���o�_.(��B=��n���Ƽ�!2�Ũ
��=��;7�<=���<��/<�_!��C���L,�G�,<z��=�wl<�Ҽ/���V=1�<���8�F =��輰�&��?��IJ��r⼽F=1��r����<�rV=DP��-���:�W����F;7x	=�,=y�(;i���:�<]��/-�
!�;!&=�L��=���< Ǫ���;FM�<I��<��x=��A�-М�6�	�b�7�&����=�&=>2r���<�9n=���' =F=�<��֡7�2j�&*D=%����<P�3</=h��<�k{��fw��=G=y�=�а;p�f<Z�{���N��Ϣ<whZ�Su-=V~�<B�7=1"��EE=�\D�%d�<Ȫ{�#Ep<B��qR]=ޢ�\R�@����=��E<oH����=�]�F�2<T��=��<W��B���IaS����<�w;�
���];/����<l�=4#x=ӽJ=����=�)!=}��m<�=����qKs=�M	=s؂=x����N�)�żS&=����=�"=�^;��ἧ��<Z�V��ϼI;I�i�M�E�μr�3�Q����D=e����&���=�%^=��+=��x���B�i�8�տ#=��=ف4������#伂R=�W�<vC�<�&r�`�E�-ab=6�B�A���q< 6`=�@6���!�t��i�#53���;1#=�ݜ�=��;��\=��=�qK=��=�-�i�0�j�<�u���K=v����R=\:/���;�#�a=Ν=��=�=X���2<�z�;����gZ�DU:W8���G��tH=��¼���>k$�A� <}+M�̾6=����HN��\X=�3�i�F�+ ���Y=�2
����<Ǘ�<J#=�ּT%Z�C������<K�<�/"�FB�@S)=�düVZ8<ԝ��r���}�W=ۧb=7HI���	�����҈�<ᒙ�U=k�&$Ż�a�i����<�)=ȍ}=·�<+T)=��<�}=i��<U�m�u��& ?�ki<N��<-�,��$���f=�p:=*m�;p,�{>�<,7���P�	ļ�
���n�<�ŕ�g�<kh�Ǩ	�y���\��uv=�A)<��1�\n�<g�<���<��<�uN�]0�<�<0KC=���]��<.w��G�8d�=��=Hi��,�<##���I��b)��t5���.��4Z<k�=�!���j<�h�����c�L=��-��~=�<��{���ʼ��L=)F%��)6���;�>�;. V�
�=��м�Y=�W�w�=mN�~ �<�~7=�\�<��n=Z��<���<���aL9��;�E=bA(=+쩻|����h������&�;޴�;A1��r�#<��n=`0r=��7�G�H�?�<R@<�lw=�i��_G��*�I<��<cx�k�=��=�����>=ӜA=�C.��^(���=�C=E�
=Vv����|��Z��5%'=��\���X<\�F�S�<b�5S=����� =w����Ƽ>L��L��C�;�(�	��<�y�<(̀=�顼�i%�Y�;��o=n!�;�<e���P��<����R�Fq=��	='`<�a�gqR;�4�<���0�"��G�<�]=�ۧ<��
=�颼з��͗<OJ�=H�A�\X���¼�ix�YH����N<WU�K�R������<P�n
e=��0<6:�<m �<�1ȼ'R�T8Ƽ����Ϳ<�&������޻�_���ü����}�<X�L=1n�;ؗ��u{F=�!�o)Լ��C����<1���I�9Z$=\�,{]�*�˼ʍN�5'������`�<-=��,������2�<i �<R���v�<������/���"���i�J�<J��<Mq�<�;�EǼs�*=a0�<l�=�3Z<!;��=$�N=�z��#H�7�=�B�	�@�J=-���>E�<	i=F� =�d;��aU�YڼP�S��?�I+o;�����9
xn=ϯK�/�w=�+D=��<Z�-���<=��a<�`��=Y����=
��7�<˩g=���<��撼�1�QP��܍���W�`���fM��
�y�� l=��� <�Iļ��Q=W�����'�<@F� �~;3�;��`���u=�6	=���;��m�x����vS=��O�+q=�+��Đ�;��<���@r=�yU�ںx����'�<�^�ҡD=�Q��?��b:=̖A��nI=d� �����Q!=o"d<��<�)+=V��H<�Y��B��W��Cq�r愽%��CV�<<�c�	ƼI�N�/8S��	m=���<9-�����K�A'�<蒿�ͅ�<'�2=sKH<l&��Q;�S[�P�
���3�<���Lk��{�$=s�[�ԵI=���<�@=�m =�0G��
\=��u��q#=ulw=�����
9��=�њ<B��;�'�J1�1���J=k�;��='�`���O=f5=��=�rI����<]V�		O=�D��I���>��!<�n�;�KK�8T�"e�<AEH�6�����x�<ո�<�Yf<������=%S$��r�Q{���c"=6�X<7�n��:2�ɽS��ʆ<(�z�T��;y)��%މ<�A���M=HM��qzp����<'�-��2�<���� �<��r=��=9��f�ϼ��<�;qA&={�c<��>=Wb��t<��"B=�� =��9<LG<٘<���<��
��	���.=A���n=H#
=�j���
�P஼���H���!~=U�5��e<;5=���5\�}�뼿q�<�`���u<�O�<��@%=�=���Z�6��Ι�P4=�ѩ�!;Z:p�<�)h<}�,=�g�#�HS=���<�]/�J�<���
�=�T_=��׼�K����<���J�p�稞<~�ڻ>�Y*=@;��� ��L�~a=�җ:q;<�<��bD=D������7�&��}c=6d�=��;<0	7=v3�<�稼:�y=92�<�� =��J��N��IqJ�W���V��B�;�G;�-X=\���!�N�H����g	�=�ؼ�0̺ĝ�<�j�<iI��e7=�Y�;�4=��&=������$�P�?�������:f!��`=��ݼ� )��
c=;L=�7=E�<�e�;A)�<�|5<M�����<v?�<2=K=�Ѹ;��<���<�E˼V� �9�"��?�p�9=��k;nL=�����<}o=�'ڼ R)=v�D<X�H�ȹ�<��0=��6=�:4=,iü���;���v�D��e�<M�?=�W����E4=
�������<�*���!/=�6�<��]=ZX�;,u�<+-=�����&J��-D<.q
=;]�4<�=��<�m�˅!�*�����ͼ>\�<YG����"=��=�*a<�p&�s��+��<�@�<'�<�o�1&���¼ś=�I'<t�;=92�!�f;���=�G���ð��o��� S��ZG<��<���<��o<��	���W�l8�L��<q�=�y�[�7^�*�~���u<��[<�ⅻ���=���n�I=���B<��<em(�!��:<{L��~���yq:0�q��q�GA"��E��\S���<���;7@�ieh�ڝ=Nk�OvL=X�Ŗ ��]S��-�K�]=�����G�@�#���zbj�x<�ȇ��߻�E��;x�<��f=vZ̻��Ի�
�<(���A��<�E��S+=g'���t=U4�<�<<�%<�	d�N�=�S<c��Iļx��eQ�� ��;��< �'=F���
<Ą��_�<���:�Hϼ��j�_D�<"��<�3S=|�^��"�s�=���c�!=�kV=*�^<8缱�	�@�c�F3�� �<�GR�).<�'[=�cļ
U�<( �<te���Y3w����/�)���ȑ
���;�Ge��-�m<C=���̾<E�N��<���<¿����sH���:=�i��� <C�<�R?�����;T�==���;oS�;��)=�����3��sn��2==e��@�=�FЊ�\��<«�<g*d�4��<:�<�t1=�)�d�=P)_�;�oP<��<=Uu�:ȼ!����Gm:�G���31�C�r�6���A=����5F=N��<> �<���e�M<��9=%���;Ǽ�/=>�'�;;&���H�[�>�9��ڼ�	���:�q�>J<@���*��^=7�j:[.x�$I�{Pü~kZ<�e=���;�cw��ye=��O�����l�<Kʜ�%#t=���r.=�����=�<^�k���1<;���W�O�=_�!�_`;�i����;�N=W��v��~s�<���<=� =@��<.X(��9u<'(��X��i�
=M�&��i=�=lJ)=Lvm�y�L�ep=�Z�
@P=˝�<��Z�	_�8IU���$=�e�<�+�<N��| 0��3@=عx<R�߻j�?�CӼƟ�Ӈ3�"�o=te �$��)���.�<�:�<�G;��O=rK=�<<���Tȼ�F=B�;=~	|:UH==m�`�'�<���T��.V�,�e��t���'[��>�<�
</y=�Ӎ;�>��%g=��MP�b/�j��<�󈼿�C=�8=�KK��&�ߥ�;��h�M+I�F�e=��E���%xV��ؚ<*���<��^��*�־�<b�"�sW=�z<8	���K=oD�;ш,=}�ȼ�=��������i=�OD;�7�<���<��='�t<c��f���4ɼ�3j�2����@=6g^<�J=����T�l���=��J��JܼD�N�[��:E33��G��=�NH<��M=j��w�7=��1ڐ�$��<��<]4=)&	=��r��=���:�_:<B�r�ܟ0����<��<�k>=7��<�t4=?=��Լ2�<=��3=y�g�ݕ=�	�;�z���;=8�y=>L�<��<�Y=�C��e�ܻ�����a���<F=��<=� �Y<���>�X˶�9��<B1��?���� <'��<�$=)�U?��ϔ���!=;�9K<��Y=aYK���<����/{�;�H=��S=�G<�W���^<�8�;i�D����%r�B� ;A՘���Ƽ��_m�<)�O��4�<ġ�<�����\�kչ<GT�<� ><y�:��N<_��;߄J<v;�<���<��{��2=!?��yN�� W�費�
0��������7�ڼp"+=�g	=��5�ٝ�<�<�R=��<<�������;�q��O�<|ƪ<�Z=��ܹZ?=s��2�A���<�M=,��;���O��O֎<��ZR<C��<��JI
�N�<�W���C��G�Rٺ`�F�98�)�<&�7��"|=�==��ʼ�t��a�����<�<�<��N��t==q�<�ܺA3��Ʃp�(�`=K�<��B<w�=����Ȃּ����3�DJ=8
�$���+�<l��;����q�2��A���a�=��%�����>̼T��?��<�Yļ��Z�U�<�	��K"�)��<.�a�F@�QLT==�+=`,����<@�	=���;5B��^����<�xn��g��.<G=�<L�D�(�U���k<�#=nhf���<�6���@2=XF=7�V<b��<���6>@=lbj;s����?Ӽ��h=�L*����:��==ᨲ�s�<�贻�;�<���<FN =���<�,��]<�!=pYV�����F�Lb���6=��R��K�<z��۸9�:ݹ=m}���s2���`=bf�=%�����=4=��`=#�����yp���K;=�#N�I�N������<��=\໖�^<v��� �Eه��p/=&�= m=N����㏼4	$���
�<V^��ټ��d�<�<Kt�~<�<N�<�I<�
=��=yo%=��Y�!=�0�<�>м� �=l�1�$��/ ;pLF��1�::��JGO��^ռ�L8�x)=�Z��e7=�F����4���1����<�{v���<A?�<}�<*⑼�	v�t��0�<�<ü�l ��^=6�<�;�p�9=��y<�z�<e�f����k�<{�S������ᗼ嘒����<X[�<��[=\V=�\��%��i}<5I <$������^¿�]��<�%$=��^30�C���4�<"P��92�<�@&=}:=�=� <���;T�u<��}=,��Ǿļ�_=d�%=F�?<� �JP��6�<� y�C=�<�p\�Q�^=���<)=��=a�м�$�=���^<���?�<��e�� Z��#�<%��<R�E<U�L;���ߵM=Q�E�?򗻨�H�Y�X�y��;I�#��ʈ���3=Ê=�g��={�dΰ;AT6��#=ۨ<��H=7?3<$�%= �<�O=������S�<�5��`�L<!-�.H�<5�=�b�<�%=�漂�Լ��o�����;�c ��ʼ���������<}�=1�*<�Ӂ�YR+=��1�6="ݒ<�Y=��x�V=��<<�碼��=s���a��!�<tc<L:_��'=���F=!�J���,\d��M�<R˿��P<'�����<=�qe�}ݶ��=s�ټot���g=Y2�����<��;0��)d;��ڹ=��8����:����k�o�<ė\�a������<`�N<{#R�ݜ����<�Un��Ѻ/��<�����<���i.��h;=4�=�É<�ք=K���'�dx�:Hr_�GA�;�՜;���<�|�<��<fJ;R�<ﱊ<�B�<�<�.=)��=�=��=��=���V@z<��ۼ��}�N�;��Z���0=LO��,�<��w=8pn<��6=���:�>c=�r=�D=��!<� =Ȝ�<�[< ~m=�Y㼦OJ�l�~=E�a=������<��	=K������|C��Խ<��
�I0���;�1��!=����V<�w>�粯<+'=�K��"=mjZ=9�B?A=��[=2岻<�<	�_=���<�{-�=��;�F�=���<�ӼV�ؼ9�����:�MH=���1�<A��<���;�Z3<5��V�n<���=3oz;�A=�Z��c?=�Y><�%%;T�U=v&j�w���W=�J<�K&;�Ё<��O���o=�[��+<��/=���ga%=ی����<��\��k���
�-�=�7мr�
��=y�<C�G�(�2=�_H���=|dZ���<�K����<w�8=���-}�<T���J�<�L��\�{�=hH����:�?{<b�^�{��;2=;��l+��>�$����&[=/��5����g;)�a<��/=(RH=
7���=5��;���%��]��<b?;�L��<ȧ���=`�Z<z��=�`������O����<߸�����:VAc;����-k��Xv���;t<8Id<���<�ۼR�Ժ��&�^2�}�T�;R��<>_Z=4MG=��0=2��	_����<�i�;�g3���f=%3���=�T�<�a=�9��;��6���n�b~3=7�lb=��=7ۼ���)B<�B?�� =mY=�Y��d8�����n��*��������<�h�~�ռ.kX<���vމ�_0��]��<4R<qh�\$J=>,�;�,�L=��)=<�]L<���<�L<6e��7�<�0=<�����3��H�<�cg=:2�<mmL=Co2�
�=�dY=�3?=���.�I=��=��<&�:�=�CR�9g=�<�4V=xѢ<'����1V<@����H;�H<�m��w~��<�^�=j�1sf�;�W<&JY��#=���XP)��B<���;�,k=v���J���P���x�<������^;sAa�D�5����<'�5��qQ=t��G~�<z�`��0�=^0 =ץ>�X��<1(�C�=�(�Z��aƠ<�^89�v%<i�<�K
=���G��<��(�;r4;��m=")�9h~;L
+=mk=8a���?=�D�:�e=\��C��o<��t=�����<-��2����;n�8�4����5=Jo!�c	;ô<��b=�W=�<=?H<�bM;m,=<�<���A=(�oI"��CO�IT�أ\=�=���<�Tk�w8%�\[;"�����,=��=/�	=a4m��Ď:�-�<�L���,=���9s�Ol���Ks�c�����l��<��/=�iz��&=I:�;��<vd�<*Ʌ<��*���ӻ|I=L�	���;�=)��JA=T�;�y��r���+M���e'�M�!�K!=�1����|<��?=���᫼�4��ޮ�5�m��%��O6��2]=����V���e=[vf���I�b�˼�W�<䭼<�x\=0��=pH=g����=���8s<�'�<�G�;7�t=�%��b�o��v��������o�E<_潼	(=�X=K��<il�F�n=��?=�<�E=$��
�<m@ɼ�H�Ig��AQ�j�A=׍�K��|p�[���cҼ��=�0I<ϭ�-�R����<�\i=�HR=��6<�춺�m��\�qv�<wƣ:�t�^�9�yJ�<Jb=�fi��c��D됼���<�f<{M��'���
����;»Ƽ���%Y=Ĕ�=@�����:�0=�1�i�2;j*E�3=���<)�\=�)��ߓ<��k_��(W�<�4㼔3���QȼN��;�'=88<>Ժ��;�;���<n&�&=D�`����&�><��@��A�1�G�?��<Ǽi�8�G=bfe�- <.;<O�ۼN�k���Y��+�D�m�
@]��?�򉾻�{<��I�T<�{L=�h=(?c=bK�xև=�\�<����p��|�ٳ����=Zt=�>0��:ȼ��ͼ:��<V��<~�|�b�&��E'=�R=�x�����)=s�$=�0E=�& �F�O��"�,Ag�\=y?ܼF(�޻�b��^=I�3�pG�i=�Ἱs4�������<�D�<�v	��t�x�:���
=�J��}��ö<h����1�|�#�XhH��f�����E=Q�W=bՔ�̱<X�f=��W_k��RR��tA�9�$<�S'<�2���`<]n*=D
=Eh��a���~��\�<p�,=*��7��8h2�)3�;s
�����<�a@=�?=�(6<=x���c<�V˼�=�d>=e#L=H��\ڼz,�6ݗ�%�=uy<�gP��m=��雼��ʼ�n$���<:���=�]_=-�缙A�i�l��;�dY<}J�:mK+=��:B�/����<JV=��=�5����Z��̼�㫼�U���=���<!.<�}��O�<�T<�<�=DM;�"=�~><;q����%�[e=�]4=��=F﷼���<��O�Eq�K1�<��<��5=�~%��f�<Qt.�,�<`�8<�9I��l<�)O��2=sꊻ`���<6���rp���=�	�A��I�<ۮ;��?=f��6+=K�R=��8Wt���8=G�ݼ���VV4���C���,�G.u<��h��AӼ�����0���,=F]���Í<�<��Z�e�y��S���\=�a�<%OI=��\=	t=w��f^ �V�Ӽ6=�1;U�=��]��lt;g"�<���<a�=�O<��g����<X�n=U��<R�L=u<�=�����<��Y�8��<+�^=Vh�<B]�<tiM=�<�����M��� =�k���;���%g�<������=�]-=�T=��h��<��=i̠<l�X��I�<
/��IX��Ll��g��+R���`=�B�<�(K�ݓ�<2=�=k�;�<�S��P�� ��ɻ�9���#<�P`���;���<�s?=?G�����ڼ�Ij�@k��E�H=���<0u�� 8m=�(,=��L��Q�;\=SD���`<]d1=2zV=}67=l˼*N#=ͣq��"=��Q=����PI¼�4�:܅�I=�{F�e�t�-�b���h���V=B�Q��k����,=_Ͳ;�=d����Q�-ꁼ�^t��:�|k�CKa���=n��s�ٰ$=�T=�H*=qCl;=r\�����i����<I��PO,��O=J�4=�}�<���E��'q�:G��7��R=�)��"�wa��*K=-WB;�]��*�(<�Ŷ<u E=��,���#<��V=��y<�G���:p=�j����<��W�6F��~_>��l	=��=��p<��<��c�-7=�D=	�;�D;�*�<����ϼa���=���[�W=����)W��^��!m	=�א��.=���"�'=��n�9=��g�b�#=eq9�(M:3�@��� =g�<8e��m�#< �m�C�1�朼�ӳ<+ǖ��N=��P<v�<{==�p�<>o�<�<<g��FM ����<�$�EŁ=h�X=~)�<r5�����U1�Ϭj���P=�tv<�N����(��w(��!�<Lv�<۹*=U�@<w��<S/=73_�����-���=4��$#���[=��ݼ+�w�u�Q=8�=Z�=kmW=̩V<傊�&lQ=�QX��~�>[�_��:�F�o]�{�s��du=�U���<���<v��<�<�9�<���¹ռ�p�<�*\<�K�W�w=�=�@=x�=J ��%=BN�Ǭ�<���<O�w��q�9)}M<0�(��A(��D�;�o6=%�@�\�=-�?����<St;�홡<8�<��<@b;=��/��|ϻ��<�����;
�P=� <n|�<(j���؛����f^���!=c�V���l���:���q�wN =P=���<n�U=2�꼉Ob�Ɍ�<�a�ÿF�U!X=��.�۽&�ЛY�Mk˼�?�:�(<�M6<�]ɼ�:�8M��;��Y�m�Eh���yX��G�<����~�:�N1�b=7<S��<���<�F=�$J�9P=~�g��%�<_�+=<N</]���R=s�:�z/=z8P;s�<�r&=D�=�h��/�ջu����<��&��V�;�U�<q~��r�a����<u��<o��f*�����<��9��==�pe���?���=;�����Kg=g3��r�:�\��]��-<�� =ǆB�vRA=�nG��(��J�:0�����#��o=ht���~4����μS�2�Y�=+:n=j�='LR<��ۼ&���'
��h�;O��<�HU�4n�;T��;��<��&O|:��4=3��!<�Bf=��Ȼ�B�;<�`�,�ʠ����~����;NI�^
���4��2X=2.����d�=�J+��&�=� <��K�y�����v��y���Ǽ`�����_��¼C ]=�9d��4�<�<�s��	�;�8ʼa�;��Ժ��*���5�����I���3#=mg��W����V�k�7���\<Y.<��=��D=x�^�vO&��{6=w�=��=�(O=�_<�����<�zq�˦<�ɲ��ni��a=�[�y��J =Z�=_�&�Hm�<\�˼�������l� <�+=W/=�/����c�ּ46<Y���,�μ
G/=���Q$z�22.�TK�<�A/�� 0�Y:��޼\h��+?7��.W�һ���=��3<���$><�S]�(�SDw��u3�=�Q=1<u�<��9�"����=����X�Z��CN�g6b��}�<n�=ӹ���H���<$Y
���<2C];�<ݼ��t���`��|ݻ���*̆=#f=ԕ=��<��4^T�c +=��G=�4�<�z?<R��-�꼄TE=	�<x�ź�8B=Lڼ|���BY_= aټ*=�<��U���ؼa@;��<��4='�X�.=[#%��CK�����4^Ҽ���<A�H=��;�� ;��o=w\=gi�<&=��^���9��<��p=U����>����<�y���G�</�:(�5=:�o��R�;�k����Z�<�<?[Y=���dG-<kYO��)���^;��޼v|��ɖ�/E�<��9<�a<.n��[,x=_z=θ�<�I�<;=�F�;�=&qϼ�1�<�=��O=ޫE=�iZ=i-4��ڼw2^=�l_<�����»�q*<���u=�NӼ�t�#�9=0���٘ ��۝�������]��P��9m=1�&��2�<�������U֋<35�<�]������YG<�G�;�~m�䘏��j~<�����/���4<UZ�H0޼c�=lO�<�y0<5<��L�����<9�n���5�����<=��l�=�<�<�=S=���<eS3=��K=s_=��X=������;��A<G��<�L�+`��8=�
ռ��<�9�*����F
;��O�����I�a%1������U��7=n=_.=��<X=�!;�O2��="�&�[�v{���~��=ڳۼ���� =xG��B �V�<틀=��d���=���<��Ѽ٥"=mg����!��P��CA2�������M�`E=b{�<���W6�E�G���<@6<��<��<�}:�h�S�<����s8B���a=Jq*=�=��:=��=��E��ڻf�;4�<C�
=��5<zK��3k�;_�D�Q�e<r3�;���%�_<�]=hË<�I������$=NJ�
�_�S%��D>=��<���� ȼp� �S�p=�-��m�=<��;R_�`�?�G�g=O�<u�����<JUe<{b�}IW;�0��V=��7=ӡμ��ؼ�̬�3����x��M8���D=�B�;��X=�WU�d]>���G=,�<1Z�<��<�3;������]�c��/q=1�=b��<n"�<,�<�	���f�ӥ�<��)��LX=?!�7�<qAW��z�����;��4=vQڼQ="l�:����uH)���Y��1=���S' ���ڼ+���J��<���<���{���i ==(�=�����7���&=)˛;miH=��;yR=�+���1=.�V��ch=� =�<ٮM��ᘼ{&=r=O=��?=��X�k��;=/Y?=��I=�m��p�it��"�2=��p<'�<�q�<L�v����<Ș��<����fȼ���J�����:�r3=�sE�5i= If��,=!��H�i=�a>=M� �G���Ҡ��z@��]0=L�	;#[-;�f	��G�<7�1�_Y�<rv��^t���==O�m=:8��(���L<���ΗƺL=�=���n���'�x�Q��~5=���;foy<C�|=[i<�{��N+<�g]=+�=��"��� =�!ӻ���OD-�]X/�=�_<�J��-Ⱦ��J�����<H�������ҽL=��=��W<�QT=R�T=a'�
5�F����;OM=��ۅϹ�] �rW=��ک���<��w��P;��?��3�<�ʼ#/<�Ѽ�߷<���J�û_��� �����	����7�<Y�B�!S�D�4�aʆ����<��=��<{A����+=�e=�~0��?q=��=p�p���2������`<��I��R��枻E��:8M3=؛=4n=��/=��;�0 F=QC�<�H�<�]�<��e��<�Yn��tm�E�w=�"(=�eC���ּ��<h�����<�x�<q[ ���1�B�.=.�Z=-&=�d����paq<I>��h=S��<屮Q��<� �Y�h���=���<�6D=Ȋ-:$[�� P=��Y;,�;�2ܼ��ʼ�-u�eߪ�{��]��\Ƽ	���@P��ԟ; �ɼ��L���<!�T=m��=�㼘c�<�]=���<iZ;<3[��=��
=8,�|�<�\=߄n=��=���e��#%=4�F=R^g=�X:\K	=-\���u�=У���� = �w<�1������8R���<�Z��vq���'<��'��Q���;E��<��=<�����c:�K��]�<�/��
��e�L=��'��<�]=XA�<��={gi�-�,<|W� �ϼ[I�ڥ�<I(=�x=� �s��s�D=-D��<���X�Ks�\F��ȏ&���I�\���AB=P�[�˶�<&��X����=���=\�I<�����+���(�!�=��x�D�<7�E=|�
�WM<ǰR=���<	�ֻ�C�����<�<������tQ�Y�3=&%��%�:�:$<�D��B�;�hM=M��<�xW�|������ 6�0��<�[���\=��mH��s�M���p�M�M=v��]�{�su�< "=;=ڍ<c��<��ܼ#�O���\<���v��<#��Vbƻ��;�M�+<��=$`�<'~��Lt��2�e=�"%�,*=ڣJ���<Z�^��O*=v�R���^� ��nV:=y	̺䲋�avh=C�^�Y�TѼDp�;�D��B�I���=(�=��
=��;��3=[S=�?=r%=�MY<ߜ��=�ʬ�D�<$)м�}l=���;N�<��������������6�2�L	=u=���ZP=e��49��ʪ<�^=���<tf=�S<E��<�O��[���=i=F��sV���
=ts��&=���l:Z�,�D��'�:���;��E���%�H�`�]Cr��D;�E3����;�s=ce�<n�=��z��=HN�:F�$=� =s�Ӽ#V=چ����<+F\<l~ =Y䛼g��;�g=����ֺ����/�<s=FQ�< ��</<���k���<�ѝ��1m�����~=��:8�;�d<�f<��;1<�<�"�<�(
=��s;syU��kü�D���*��@�%=m�|����<�T~=I�Y����\W��!�:��<U�#��L���-=)ґ���(�XHӻؔ<�.�Ɔ�ǟ=�Q8=�^=u:�D�(<���<�P�<��<���e�M������*��ȏ��kE<��Y<�$V�y� �H�H�P=z��<��M�PDm<z|�<cJ=��������vg�S���.��5)<f���$<[��<�տ���n=�lS��@<��z�KE#�թ;�T99;�/=rA溠��޸==�[�$#d=�[��5�:�+�<�9��<Rk����R�EG]<�<��6=�Dm�v��<�P���ǻ���<���<pFj�>�2�a�F�[[�<;|�<���<�%�K耽��x=��>=i"�?�~� �2�.�M���B=v
��	!��U=:O����+�Fn=/&=�J�<�N�ĔN�e��;����~��B�1=�"^�t����;]<���6=��1��+a=J�=���<�N��{�"=�@��d,=j�&�I(q<�4=i��<s�+=��,;����P6=�1���=�� �=6���$䂻�<�^<���z;(=��<s�=U�<
 ��Pw�<�D���+��Ћ;:@����U�/f2�u�<�9=��I<�����j8����
U�<�f�<�uI<j�<�� �46�l0���z=DJ���,�=�6����<�k����p�<4��;6?�4�<`%��=(�s���;�q����<.�T=&VH=�M��1><o��<�&<mb�;��-���=ҡ�
���G�F=��=�z��|�;1�T<f�o<��2�0��ߣ<�<~p=��B�����[�G~�<��K=!�� �<�S�р�>�:}�����<ֹO<wi=Iia<�=#��<?l�:
���=��<M�W=k��m(K=�w��+�H=h{5�mΈ;}0e=�����N��ѻ��<�z%<��+��Z��{�1=9Ѣ<���<��
<�5��:=g�z<���;c��l�Ԥܼ�����:��<T)N;=OXZ��bK����<S�xzݼ�G<��*E=��)�����=�<���;�m9��4��Bg�;��<p82�d�{�*=r�O<�/5=����s2;P���"����<�#p��D$�B K<h6�Ј;=Q�;n*���f=��<
�3�`'q��3=,=6�.�1%<wƤ��,l<�F�����.>=�=��`�0|�<��=�,�<�z�@"�i=#4T���+=/�����=��쉻�;8粀<v�Z�#��<<{w<o�Z�(�E�p�S�R��<:WW=�E�<�l��}�������
<��;jS�����<߬/<7C��_��<��߼�僺�a�<��;��h<��<|��=�WԻ>6=2�x��Ӯ<ʊ����v�!�	��DH��i=׍M;ѽR=�*=�]<�Oo��tE<�i����<��v��f����?<���E=�oD���'��[=�C�:#��;����c=�Ǝ��2X���=O�:t+p�������=�p�=�|�<�e����1$����H�I�s_߻G:=A+ϼ� z�$�	=-�7<v#==�����9:��3=W�=i=�<����N���	�pm=0���ò���Kȼ�p=�o���!=�'��F:+���n;;=�1�1 M;K? =W�;�?���;q���������e�����
�a=w4�=�K5����;Vjc=�?4<��,=���<=��y�c�{}=T�y�WL=��=�Q<����u��tY=zS�-<ӻ�Ԓ�@���=B.�A�C�\H������*���������<�`9=R�;������m�z<��;���<�:�<h�=z"P�RW�W�����<��p���3��)�;ė���N=��<����[=����y�����R=oi��'*�B�\��`,=^���<hi�@�l��<�8=�*ɻ2O=�J7=i��͇A9��������-���=�6=��>=6K3=��!=O�B<p3=�oP=�����ऻ�q�����<��m<�t�X��<Dq���,<g�/�%���5��<2|�/Q�<�<��<h���?���Pс�2�}="M̻�=}� [�<�񩼡3�������-��4���6퉻�';�Y5T=�P=!==��3^=��/�]ۼ��"<f�6=	�.�|�0��p�<m��:E�=�����#�<�mN�	/�_E��.=t.��I�I=��i<օ�<J_!�u�#=U�Z��[����:����8����;�M�<��>�1�ػ�{<�QI=��<��ּ+���9";��=��<�p~�y�K���E=+�˼��W�սμk�<�j\��'=i����v(ʻsx.=�	����9�!��=��B:���<��?`]��k=�Ή�[bD��E+��r=���=�I�<�]6=/S(���A��8�<�k8=����Ȇ�< �7=�/=zȼ_H?=�?�<�ѼE'><���<qC�<%�i�o�=S��<����e.=����(���&��I=�����D�(�=֭=G��ط=�b�<��=V@0����<:��<5qf�H�ٮ켢Գ�+F��ƛ<�A=�=��C={}r<?r+����yJ=$�=�P��!�Q�<�5�=�=�'=N"��=uk=�Rx<�萼h�;	��2�E=w�<��<&�3<�H =�F<V�D�<�d=k�μ)$����<ȇ��Gʼ{�<��a=��==BA��(.��0�<|�<µ�r׼�i�<}K�D&=.�G���L�p;���/ܼ�N<��#=�\=jB�<t�s[���P���l|����&<(9�<x�'�	�<�cѻ�w=|�=��"=E�3=,�#���	=s�_��=�a��u�<K�ݼ�M<���<QI ��1-�i�|<���;�ļ�T����>���xl<�
�<gmj=�Jz=���<�	<Af=��;��D=�Y���m�<��`=���<�͉�7��h��h9�S�7v(=1]�:-"���AX��M�<��Z��I=<վ��d�4��̃��g�V�=�[O=�x��X'=N�<��n���2P�^���,9�<]���Ttt���:�!�\=�
�<1�<�'E�K��2 =�,ۼ�`����C�Ȼ<�¼v������<�:=�Q$�*]��}y]=�4���i��`w=]JF���μ��=� �<.n>=�?f��#���"=cZ�<��t�n溻W0��II<5��<�_8��<�=,3"��p=�˻H����,=�ou��o�:@��;@a,��厼�?�<���n��e����Ӈ=e�%=r�+�ȫ�<ow�<�����=h�(=cC�<V�<�=?��<��O�<�xb�����G�:n���<�ݲ<T���;��=�K;=��l=�J.<��<�N��G<����:�˼�������ܟ<.S=�=#�����<��m��t�< ���4c%=m�Hv@��zz<:�;Yآ��L�:Ţ%=�>b<I��Lh�<vf�<C�A=�^�,\�C�_=�a`����<�;<7�)�0m׻3��=f�=r���VG+�ɔ=Nq><KK��<
�h�"=�"��u<<�����<�O����=AON�������:}W=(	4=O�G�T=�k3�np�<��K=��V<��;���臋<���O���@ټ������t+��6���~N�d�%��|G=z#������.�i8<>r��!�Dy<�v�<��m=H�n=B��l�.=�F�<���<}s=*nf=�v|=A�h�)�������8�x`P�l������ED;���'����:�/R�
�=H����r�<eoT<Ii�o{=��i;��@��`?�,�<|;�kɩ<��+=��4;�<=b��;O�=��F����<)?=����=����Z=�;�
=c	�<�%=��;�ۢ:%9:/��F=�g=��<jZ
�+l�<ρ�<)m"�HĐ<z�<��=���=iD�<� @<h��NN�`B���M���=X�A�g=Aq_=1[%=��9I�Q=w�X��+��꼚8�E�<\��<�P_���m;g��<��h<����^2���.��^�<��]�-�<��F���\�d�<<�J#=�ӱ�?f��r��::�0=��ռ��Ȼd0=�_=�.	<ʑB�g���T!���������}��sE�<�*����?<���<�T�]4=�&���}��n3��dB�-�r��?&�r�!;ߣǼ���V	�;�������������^�-=����t����Y�:���<�
,=)K<��U������ӥ;Ё�N=���<	O{;t�d����<�_i=�L�j�=��<K�s���<�	�<�)�<�P4=,�.=�n�$���M�	�5��[��x:�<*�0=z�B��z<?L��^=Y�{;�D9<e����p�;�� ��<��L)=�1;=%;±����a�<a�6�\%���f�[�;]����`a=����h�L<�c.=!QP<��7=�x��T.��j����<�S��
G=+ϼ칔�邦<=�@�����<w�Ѽ'�+=�ɼ�|��GN�yN�<�w�<�;I=Q�S�W��E%����t������=����6=��j��뎼4zW=���<wg��I^���<�O�� K�ht1�;w���(9�d@����`qg�>'I=�)��墼�|=�����C%=��]�=�+4�'-�<�R��H�u<�D<5�n=��*����<�l'==����D=C Ѽ5�@������#;�▸`N�>G$�g�=N���鷼&<K�(�|s=H";��m=;0;�6ּ�<��ۺ%$&���}���H<�?<�0A=YWҼ�'Ѽ,�a��mj�1�[L$<Jo��ϲ�<�v2=�\=$=��)H<�,�<�1�`Q=��<��S=��.����;Ťϼ���:�~<����=�Aݼ�/�<s�G<���;���<��[��*缬C;ET=1Rq<�&<� ��7#����vV=`_���T=P=fN�<9S�<&���x�쑫<�ѻ�6;=z��<��.���=HIX����D�
�v�=*7n�,��;m�L=�Y份�-�00�<�,=q���q=r4��䒻�/�<�(�ս�=��ϼn?�,)¼p2W�~*;E��&/ʼY
�<L;Y=���^`�<�Dr=6W��	Z��݆���y<�g <ž=P˼P�f=��c=
z��ka=b*B=��?=�L<mu��!9=�3-���<p�#=��#=�G¼T�S=t�� �<f;[�~ռ�~�;-�-=ش#��K�<�AF��5;�q���h���<ƇG=e'\=�2?��z<�DqU�3�=N��:��H= ~X<�����̼2��:URb<y�@=��;@=~�=^(	��	a��"��D�RPW�B�Ż��ʺ���ם�E�<<�W=�+��$�K�9<~K�;�u=���#=�Q �\=� %=�z4=�b���e�i�ͼ�6����<�LI;|���Q��m�J<k,=��[����<��3�a��X⼘X��Y�<<"xC�x�<�ʬ;]?<vd<�@�;�����֕<#g:=&�<�qT��ڮ�Ɋ1=�ޢ�<�]��
(��ݒ;a��<�p�xA�<�n��g8=�L�������R� �,+��D=�9%=֬^<h�u=���<[����<�=�o<z�<+hq=ۈ�f���:�cX=�x�<Y�<=(��;x�@�ںx��༷9_�z4���>�<�����(�c��-[r=N�B��:�<���<��]=B�P=�n&��ǃ=���<�Z���7=s̼��`���.�w
��T��KT�<�~/���^=����E�<��޼��Ӽ�3y��q¼Ow�lR-=v���5"�3h�<Ê�<RZv�L-@��v����<u���a)����\kq��==�4
��0x�ӹe=K%��1�/=Rc��B�<G-�<��<�kڻ7=.#>='P<�Fq=���A h�!f/�I:7�'�!�ۖ%��D�<`|�p�<�%J;Ugǻ�;=���%=��<�JU���;��<��A=�p<�����w|��z���<[�q<�Rg��4<��i9S���Լ���=�7=�Q��� �̀<��N<�h=�c�����7{� Y=�H="�O�E
]=(�D�[�#�!+�<��=��<�/�<g�=߷	�Ӌ
=�Z/��=%�F�<��,����g��<�𥼷q��
�<Hi���@�R�y�O�ļIG<U>�&1���,=��A�z�;ٶ=<��2��s#���%�)�<�!Q=�Չ<�����"<���:��#=�ɉ=�A=��B;�W=d���H.��9A��~<�*��K�8=EnQ����A���-	߼}��<k��:��'��Y.=֒=�"�c�I<&U��a2����<��W���<׍N=6#���\�:���9z�=��<��!��p�%<�g���wE;^�=#ۦ;)��%�<��μ�. =�&�5���=׳�:�p���m���<%C�9Ӣb<�rZ�R~R=�=N�F���n2�=꾠<׸��Jn=6fP�V�@=����=�b�E�=�@[�uO=�ŉ=K��D�<�л1+w<��)eR<�p9=<3�<���a=o�w�%�S����:��s=D�<yZ��(b�<D�6��1= �!=^Eڼ����H<�7�;��J=-I9��Mj<x�n�r->;��`�1���&�$�0�+#,���L=�����(N<'���_iƼz.-=��3<����<Q�-<���T�^�L#�<�����<#b�׃
�8�:�+�u�Ѽp\ϼ��l=J+O�y����VȬ<�r=%�;���:�=k��<hr�;���<x��<��-��ǣ;oq���Q�ܖ��댦�6��<�:=�/�;2襼[x	��D�<&nS=4�<H�,��"r=c]6=@�]=(����0�<眼�Y6���?9�Ӏ���~<V���g��Z�<ѝr;OJ@<��*��M=�#�#����w&<yMV=li��T�<�RP�ɝ�a;�;Y\Z=��<�P��
��
�<iu=yrɺa8������W@�<3���%=C-</��������<��G=��<���:HL9�3��?�;z�Z���<"n:=w=<�=��� 	T�D�F|=g臼�T=���<���<���<�Xb�ڞ���=��
��v�:E�v=T�����<ӏ�����
*�;_��<�/���.�B��aj=���;��U�g�5=C��U$=-\9����*����<�ѥ<P��;���</s�<�=�E7�:��<zMW����:7޼;�= �G=�-=���{uA� �e�:F��:=o�i=`H��g�<���?/=�5
�Me,=ƿ<h����ڡq=��6��K(=��<�= �ؼg����/�(2=`�<��*<�Z=�>��u<����ӄ<މ�&��<E�3���7=�j=ҸS�/S ��/W=VL#���!�T��:��D�����Z=�L�s6�<ڦe<�[=Gf)��I�<�p'<?�(�jE�<�69�o��|�k��V<�^��x�<�Z��M��!<����!$<!���8\=Ig:��"���<��<��#�q�!=��;j�=�!�<8@(����C��<��.=Fd��jl�\�ؼ4�˺#=�Lk=*�λ���-Qx�2�=*��<�쵼��&=7ؓ<1D�;.��\�:TJ�2�(���='��9�?�<x�;=�����W=�\==��Z=�6K=e�8=U~n=ہl=���<�Q�G��<��a���<O��Jf�<�5#�n}0����&3A�Nr,=}Y,���̼�MR<����a7��<X=y�.=>�[=KTm=���9�p�w*�<�y����Z���f�EU��hI=��Z�j�$=�+�<��<z4<����9=8fN��F�4.�:��`��#��폼�=s�X�7���Wi�@M=��=�ǻ�E�]�1=d2=�w��S�����L� =�g<���=]��I�M�4����;"��:���Н��g6�����M���;=S��<�.��fb6���^�H�H�{Ww;�9�;�46<�O%���O�%v㼇I=3E7=�VE�]���B=�(���5 ��D�<�K<$�@� �<d�Z=1ݻ��"�R��<Oٟ�71�<PF�e~Z���E= ܠ<��s<{�1���\��?�;��t�2�i=�IM��[�<qu���ds�%�_��s"����<�3=��Y!�<�^=g�3��������^�ػ��5���=�>N�� �<k5=x�M<�o9�м�Į<�_�<��=%��<�DR���$=�}D�jU\�.:�����RW9<Sۺ�)�<�F��ԉ=�HH�0�r<��@�"V�<��<t�o=�Mp�M&<ZS��L`��E�E޼�<��D=:���'ג<-)�\X=P���=�eh��qV=<�ܼ�[�<^l=�F<��<9��Zǈ�=��<�}%���<���<I&<�7�>l�<��^�[(�;&�Y=�n�;k<�Q���!F;+;=�=[H��ٻn�6=�$+<����hP���J�U��<���<~w=�׺��<^H5�,�K=`QU=Jα<��,=��@�_���i<�yj��C=�y�<�-̼U�<4'�; G�)y=���m�A��jw:����(�0�f=؄	=����\��_��<_:L=]@�9��Ļ��~� B�=�,�����]������ʳ<w2R���B=�����;n�<����#��<e�=�w7���f<[1T=��a�}uB=����&�E=�rk=��<�P=�>�'-�P�żR+=��C="4�. ���T��PJ��Ƽ���<\�f<�Ad�`C˻��,=��<�M� ?���<�n����=c@4=�I���rg=pG�<��Ҥ�� ���`�Jh;�<�Z]=/�l<-+���=-Xe=*��;�v=��S=Y��x�=�	{�~Q���H}6=#"L�N����O�F�0���j!�o�<Q����7�f��V4���i<�L�<�}��v�y=��<=��;�j���D�G���Z���H<Ը���<<���=E��;�%���A�X0�5�X�A+=�?H�_j]=��M=��ּWퟹ3N$�n<6�}�%i;9<<��P�L �<�=_�� ���:�S�JsW=�5��*)={\��1=�;��U���� �{=
�u=�ӹ�W��<BP=��Լ(�=��%��?��D�<��8c=��0=)�<C�2= ��Ƶ=b��w�9<���<^W����@=oT�<Pp�<�X=d�<�c���i���=.�&���p=���<XP�Z��F==2��<��<ƛټ��e�6��J2=�
'=��<��s;��<;�R伦U��M[6��O!�!1=�	���-��:<,�<�a���a<�
D=v��<Ԝ�<u��u���:��Rm=`<���<����fP�~$q�����Iz;}u;�@�93�z^==��)�4q �����t�Z 6�ua=��h=�ܿ<�����lE��=��%��Q��a$4���&�"��<��@���<Y?��'Ӻ'�%='U��7�F=�eμ��a=S=Y���mSh=�H�M=[��<���;�䄼v�<.,�<��f<��6=��G��M�<~T�81ü���<  `��_=L�_=� q�gE=������<��A;#<�R�<qŷ�4��N�����cM=H�)<Xa*=�h��|W�b͒<c�Z�ǘ��nM���;�Z�o޼������e� '�2k=r̰<@�~�|�=1r<00�=_ߘ���ļ���;�,D��"6� lH�
N=����<�G=�<D�=�V/�>�,=7��"��E�;�ͳ��`$�U�48=��3=#��g��<�F���V�N�;<����s�3=� %�9�;��*�x�,=V��;1\E=-��<L���%��5�a�=K1'�Ze�;0=�$��#B�<$ᗽ�e6=Q���P�:��8��>;է����<?ӌ�S92<���hZ�=���;�=�R��SB=IA=��$=���<��=�:�⑻9d=SļA�Vh���<AYy;�*Q��H�< ��<�Zl<��Ƽ,* ��s�n�<�d¼ y�<���<����6�S�0<cy=^�J=tV:��I��t�=�m"���)��줼�}=������<�D�<.)<����=��<��A�^�ϼ]\;�I�=� =�ѼB:��S"��
�5�J�@��U��<�}���R(=L�����[�;�p1��vZ<��=�=o�$�����y�-�{��<�]<b������;��,=�b:��&=�����)=����� �;�����I����T���=�{����</���Y�<���=b~V�p`����#�T՘��=S=+�c=�r=�f:=��@�S�@:7��<�
J����<��=J߼Zu=?k$<Qr<�� k=_��<���<��<-�X����n��������C���	I=0(>��A��k�d�<��;��߼=c#��n=։�<�쫼*�=EP�d"T=o��<�h��G3�2i����u=�����;%�(<��ۼ�����=(='_��n��8�<֟.�H�s=m"�@�=G�p=�H]����:���<��=\Z=ꙓ<Y�<��=ۘһ���<lHO=!/2=[!�^Rv<J�<~"�-�=�K=(��E��<+�k�<o
�<�6=�=�=�W=Rى��`��G�<j���FʼZ���<�Fk�-`�N
2������fv�Q 	=�9=�3s��Z=������u������T�<�=D�5��YK����<�0=F��;'�=��i�B��<���~�=(�!��׵�q����<��?5��1M���=y=���,H�<�A޻��;�K�<������s���ؼ�>D�JiN�J��W����<�Ǥ�W���mļވ.��*<I�p���9�n�*�>�=x�<�������E<46=�?��J�|=�=ES��\�=�5#=Q���Ʈ�o�����<v�C�j�+=|�;5/g�vW�2Y=Ķ���·=[EJ�7�i=C����=ՠ�<S�8<�{���Lû3�A=����;��x=;C<E�����=^>,<�/<��\<p;���	;`�$���W��à<�Ï<��C=���<�W�<㰳��#���<�|3<�J�ƈ��(@��ި����;�K���)<�z������B�A�P��X�<��%��h�T/a=�w7�;<@�<]���u?�f�<_�@������j<%�<-�Ӽ�7�B8���R=b�<�A�۵A=�q�8�=�\2����;��2=}a��`�L�;������WY���<˙u�m�����=hk�� :m�v=�.�;i�伲l���T<�H�^�=;�
=(�;=�^�u="��<#΀=�^�<F=���<%g=w�}��g��*����X�=���<{�C�Y ;=�@9��A�=}����0��O=�� �A��ڿ<�d���]�p�=���~��<�P����B��Mż9�l�Ԍ,=Rb�<tv�<f򻝡A�R;b�V��!"=���<����}�{��xB��C��x�6=_,��;���R<>=]r�d/�<���;C�;��Q=�7%;Y2\��D=��u��<<r;<�V]�U��eX=/=1�B=��_=�;<��&=��漖�=iXB�I�/=(�m�L=�!���;����<ia�<9�=$1f=n/.=X�;2�-=0 ��"�꼀��9��Z=�T=��@=zan=c�<S�輁�<�뜻�9C�h{ =�]=�������;ia����<�|�9���/�;���� r��Z1�<�/<�ؼ*�Y=0�<Lp=^�=�,�<���<�TG=0�<�?=��l�-jr���<���<���<������<�u���鼶>�@f��}�2Mȼ��T=�q�<`��:O����<��r��{=��B(���z�;l���.=����7�:�'=j <��;�ʀ;���<b2=E'�|N={a׻Ѓ=�,g=Mg"��w?�J���5�;�.=��{����;r!���,m<�n�a���Ή�꼺<�39="aE����<ɼOZ�<HŃ��F׼c�$�;���#�eP4���E��/�Ʊ�<�5�;i<�G�L;4=xj
���3˻��[=��;�US�nS��"�M�:��|�<����5�e=�ȼj��]��,@S����;-��<W���ƈƼ�C=�u1=Ֆ�Zn���=��U=c���F\ܼf��=�@�����|:Mz6�Q/7=��FL[���R===˕c��뉽q��b;�<��	��b�<#��<����f=�<g=�[��&��+ɼSn=/v����:�z*<��==���s��5��g���9�S;�<�cR=�=E���9=B�Y<c�
��_W��tm�K:�ܸv=�3������0�<M��;]���=<��5;N�Y=�Fռ��m=&:[���#��M뼀Ik����Y�����἗R.=ŧ0=�ԑ��F̼\��<�gE:�g<A�)=N|���sJ<�纝�v<M�`<K��<n�n���0��z;��N�c=S�&=����*���-%=n�e�� �+��<�eP=�����3�V;fر;lzH�e}��=鸦�I�����<zV+�㷼0Z���6����<e�=�=���	���X�<�\�v�P=�.=ק=uL��)��	�;K�#�M�ĺڙ�<�`�<�r�;![�%�$���<D
=�kY;��!=��+=2TN=��=6�q���A�o>==w���U;p���k��)��dD=ǃ'=I�0�״=<��i=�Cϻ�k=�po<Pqg�/u�<ΐ�<��L=$ �����^����<�W���%<yL�38i��?&�Q�ӻ|����ė�BP=w�B�8sc�,Qd=�{\<+#�,=-�Q<Fn=�I�<�������?!��`Z=\%b=�N�W	7<#!�<��{=o���w��37�=���<��<do�����<�B�<
����G����S�=`<Y�޼5�d��EK=&�X=�WM=s/�;���<�E<9�ȼ��o����<�)ܼUg���0=kxټ�&Y����y�C�e�է+� ��(¼]V�<�sK<ż@��H�T<���;P=#���<.�;s�?�7>==�ϋ��r��-`=��<�@+��˻�l6��0=�
=F��<�0�<����4��4׼�A�<Z�l�)�	�� ��)<(�)�
�ż\�<"'�0q4�W��<�ټ�7x�	v�:�F4=�^/=t��=�9������4�=�6<�K�:xt޼!��<�l�<à-=3���v�<�	<e�	=/q�����;�'�<�C�;v�Ǽ� Y���K�eR[�]�%�~<��=��<�R=n�$���'��ļ�Ӏ;+�κz��������H�=v�a<�N���<�Ze=z	m�6�&=�WH<M��;k$+=%�;o�T=��h=м<�1�<ߚs<�57��I=*���Ѽ ���܃�<��\��,V�@�H=p�v�V�O�L=��<wH'=��=#�A��=������ �g��4������@��^�<h�
<������}?8�Vm�<���f��<}<��=�&G<��=p��<��k�ݥ��+��<��A=�Y���<j��=�$���8<�Kü-A6��U<�03�w��<:3�;G<D��S���n=�=��g�y=�'���;�i ���V=-���0�ۋ���b���5���y�=w=z0=��l�we�<�O=��/=�	���s�:�2�H�<l�̼q<p�	�kN�X��C��?q=��g�����Q���<Q7�~�(����<�����m���I�ǼK�h=�k=�Â<��<��=ԱI=�2�臼�e�<������<{��=?�r=��:=tm��#�=�?D�%�����<�ؼ��,<&ٺ��yo��&��V��%�h=a�<)%!;��&;50�I�ϼ����z=_CA���<R?�����.=���b���{q=���Θ=6$��i�n;h:D<L��<�cm<G!<����-'���,��0�<a4����<�*�P�ּ=�>=��,=�I=��=���<�¼>ʮ;,�;x8=��ܻb�L=�ٸ��g�=IB�;/�-��\9�|LP�fW=S�����{Oe��Eʻ5}4=� =���<��(�փ�<ī<8�|���3��A<U�<=A����[=��<[D�=�<S������P=Z��<��J�Ť=v7��U3�=ν�;#����z���L���<=�ju�ɿ�;.��<��B�m^ܼ�!@�#B=�F�<~�=;}3=u���]��<�.���v=�,�3��=�o��])4����"<_:!���Z=����LbY<�=�����{�5=�w�<	���)=� �:��׼i$9�3*�<�H�<x@=��{=�9=k�{=�9��|;Z�K��}(=��9(V=��*��1C=u�������v$=��=oϼЈ=r�"<�Q=U4�<�T����$��<y(꼙�<��@=L =w蔽U1>��6�<L˩�ûu1=����Iл?�p�h��P���x_���mU�<;�$���
���=���<� ��<u�<��2��='=����M�=s��:���<Bϗ����FC��"�<�qo=_�<=p��;	�/<�>=X�P��Ǽe�I����<3ؼ5��
q����w�X=�*���h�JBD=�L����W�n!=��':���<m�=��e��$=���<Qf���X�<[�D<5�x<c =$��;�S��C0�<�;��5���Ϡ<�(=cN0=����]�-=�+7�
�s=Bqļ�G$�<?����g�($;�� <���<��;�X���QI��1N= (�虼��'<���&#@��#¼���<�ц�?���@4�x)<��S�;�%<u4
=�(�<L�޼��t�LL�IM����!��n��jX=*&���<�E=�Z =�]�<2�?����[^������d7�t�=�Z�<�=���:�M��Ȧ��f$<a<L�G�;��3=�U�<
� ��3�<���;��=�Z�<)=�l��	���x���=�$=�u\<
�4�(�J<�Y�H��:t�<��?=�==3�<<�;�<4��� 2,� P=��=x\켟_��༼�m�;��<yR�<��-��7����v�#=	!��F1p��y�<�9����;� =L.;��'�|�<����k���Nj;�f�;�d"��;�m�A�^=���yN<�*|;�� �b�.=�*���}=�5�f��qX^��2F=?1w=��d�<5E=%��1�6�$;�6	��&���
�<G�����%<��0=q�:DQ�&n��
�:O)�.�P9��)=rt���<�.<�����<����al=G���T���m�TF��uKN���H=�=!r��h*���_y;�H_=#�<�}<8�Ӽ�J�<����1 �}�6�Nr;}�!��]�_.�<s�v<��b=�[�g̱��ৼz�X<lg߻u3����Y;�7��<V"�"�<�н���<*m����<�`�<�m�N�(=�	�<��<��(=���:�<s �Q�D��={W=<�y=�֟���6��bN�lʍ�]1y��=�<�!�<�S:��Ӝ�	��<�N?=L��<*F�7�=J!=�@л55o��Gz���������@���4�z���߼�"=�s��S"�������;I%�<�}�<c�;=n�:<DH)���;̂T=�䏼r���L�"�(=Ʌ<7[�:N=٦�<��=��a������{6����&=t =+@A=x� �ݼ�<��<&@ü��'�U=k���
�9+X=ݼ�����`�@�-#C�K�^=LZ\=��X=������:_a��<�Q/�<**ǻP2�<����ev	=�=�/�{�W��R����;�/��f�<m��<��*���ڻ$r�����^=���t��	f�0����u4��M�<R����������x4=(����;OL���3�<
H<�*����<��=,:~=��.<��(=�f)��=�^��L/-��%c�x�n���<-��<O����S��OI�=�d9{�i=Іf�So�Lo�y�G�8<=�+=v\����<���;6.=@�.=�2H��S]�1�==2�缚и�����Lܲ���k�[� �	���>w!�G/F=�T��p�;o����%�;��=�_=ѼI��_6����Ҿ�<�k�<��<��<D�G=S�;*�,�3p���=[0��X�A���;�D/=��1=1�\��q��* L�<��<nѼ\|R=�d8=2�<����.y���
=o���&&�?��<����O;�t#*=+o��G=�O�����p�j����:K�'��`��EX0�`�G=�5|��qJ�)3��j=a�;Ҕ0=�@=vf0��!�qs��y��������d�f�����=�P5<X��<��6=�L��]�;ݼ���i�=�ib��P�<�ټ��q==Ni�&n�<9��<3��;��󼅁�;̓=�\U=Y�:;�Rj���Ӽ@zJ�A��C�h�S��=~f=�Yq��O�;�櫼�zS=K��<=3R�DK�<��4�<i��q��<�~:��|1��8�<�����-��h��=v|1<�]*=i�<]�;<���Y���x�owO=#x/=fC=!`�<�\<�!=.s*=��<�Ո:��ĺb!�<�R��݊���I��r<�.���<︴�;<�J����@=��=iߧ���2��X��'�<{1��Rl=D�<aQ*=$��<��v�Dy����<�{�3�=����5�$����=]� =8�����,<���;y{l=\+����<,'�<	�E�^��<��;ɋ<�Ώ�Z�`�n9T<���<Pk=��̺^a�BJ�;q�:�)�@/=3�F�*<��+O�(��<�Km=��
=�����4=�v}��5�<�j<X�a�����t��<�|��(/i���ɼ�=0b==2��=nUz;���<�p���L�X|�c�1�Ǉ=�E��~���=2x$��T4�-��o�	���Q;��~<�#=N�8�gվ<ї�<�Q�x�U��Xc�����:�:֛�<�o<""��7p<���;�UU=���=	�
�Mg���=�9����{�-=I��:J&=T��<�Cp�GD��?N�<�0�;]�S=��=Ð�	�<�~�9)N���_<+�+�ZL�w�Ha;g�p��bR�\��G��<׋��$c=n�=���<9p`<
�;=�J{<)�,=��i�'S�=�m=�v�<x(<�8=��мҏ����[=�fp:S�=c'=T
=�>/�ޠU<\+��03h=��6=xD�;��U=�99�Q��c��e�,������#>�Y��U�<S#�{�$L	=]Qc������R���U�a=\&=�0='O�k�TG=��f��"�:�)��s=��[���<@�߻H�ּ�"X��+���Kc��8�	G��M�Z�z���d�aO<,�&=�20=	G��#J=V� ���=dH=5�<�@�<e���(]�	C񼥼z=�>�:�ޟ�?@&<Y)=�׮;l+�< K���f�<|�^�s�5�<��7������!;�=�c���f�6���J}��B�;���>�; ������=A�����=�^μ�q弍�\=���߻�<��>��J��0=�\？+P��v<��-����[&=�х;�����Y�zꆼ3$H�|2;������<�������<ڃ<�-H��h9=����==�K
=�0���N��S=�5"�&=F<�%=�l(=1�Լ���<�0�Q�=ToI=o�<��m��Bû�6<-0���!=�֧<���<�=�(S=b�ʼ�w�NM�<���<��D��~�<Q�5<�iZ=�!;Q�8<԰a=X�q=K��s�o]�<�W�<k�0=H�ټ��j���{=��ߺ��b=W�׻A�i= *��˩d��}�m�=�	'=�f�:!�����6/<_	˼�����<bDȻ�>=��h�n=0-=|��<��=,M���R�IѾ�d�-<Fcn=�)�<�)$=��$�Ut=e���=��;�8N=�]G�"��;�p;��%= +ɼ���w��<������<>�ؼw'�<�!�;K��;�]�1=�:�<��=5;�<!w�<�Z�<e�(�8�];]V@�e�ɮ2<*�D=�9$;�<{�@=$�t�����a���t=�'$��ݻ ���N���<ټ��8�1�<Tٻ6ȼ��m�2r��PJ=Xs����A;ǼP'\�dٶ<��=�i�<�S*��B=j�漋��;��ļ�㼻��<��.=�@�<{ҍ<����E�<xO[<B��<%/<U^�<9M=��Ļ�1��Ah����9L�����:�m9 �<I=�I=,�<l�<���5	m<�U����r���I�:j'=�jϼ`a����k=9�0�� �;r<�u���I��a�ֱ�2=d=����1��9<3�I,a�-%,�#
�� 6;.�_=�r�;�1W=��}<w�[=J�t������O�\:��<=�I�<���-e?��eT=M�Ի;� �I�D��q�<oqY<J���W�C��_��g��q�V�T���Ѫ�e�K=TDG��,=,�<)?��c�k9���+=�-�p0���� =-65�F/<���Η7=�c=��<@��<�9�?��<���O�<yn�= a�O4��M�<A������8NK[�󨒼�=�s*=6�z�x۸����=��1���#�~�<d܍���<��/<*��<]�ٹ���<�zW=F�L=R|?;jU=�� �K�=�=�8���<�q=�H���5�Wt�m	<=2�����1�<� ��Q��<Ps����<������@dZ=t"�,�Ǽ�&�����k�4<�o�<�(*<E(k��q�;�u�<ֶ�<���<��=f��;$M�UL=Qa=�\��4�B�i���N�6q*����Ck<�o	=L�`<+C�<���<`�+�>�<r?��P��� %=�-E=d�<�Ny;B;��"d<[���쬼�N����B<�4=^�=.���k�Wn<������V�<2���
�缬�?<�*�<�>���<���;9��H&�0��x^)�:d8���~<�5����~��z<�g`=nWN���b��:t�v=��A��I��T�*=��l����}v�]���-���͞_�:����,;,(�������x���P<إ1���/��q6�w0����X��߼j�P=���=����� ��P=7��5hY���v;z�����<�=�5T=�mO;WԼ����I����=x�f���q=�%�<�J�=�Q�{H�<��<�g���!=f5�<���X=)��7�1<%�K=hL�S�&=����4,=�x�<ϱ&�b�;;�Y=�+=�hy�"�v=�v��"6=n���Gj���<��E�m��_y�< ��;:@d���ӼwS!=	�ۡռJR�<I+E�+5D;C	M�\��<�����s̼�`�<��<;=~�= <g�ռf~���K�U_��h�;%=���=u�Y�z��pB=����G=~-�Z~��NH�a\@��4Ҽ��0� g�<~>��?r��0<�0c<�6���d<�9l����~d�V�����2�=FW�Jt =,�v=��<c�;�i}3<|�T��$����e��q��q�=/7���$�׏����=�{D;d��J�E�����>O��"��Y�7�=���j�:�\�<�9�9�-?=̳=;\�;�u<y8#���<���<El?=t�輛�<F>;��=d	=T=�`q=
	c�6�޼��]=�臼C}���m5��@q�>U�����N>h=�ي��>=�~�<�u������A=%�=ˀ4�6�6��-$=t�n=N|s=)UB=dTx�GXZ<�5P�9qz<�/�<�%A��Q ���$=�H��6Y=u8������ʼk'���S=aZ5�c�<r��<�j�sW�c�R�Y��<���;IB�<��<=b=�l��=6Q��>%�A�n=/-y��:།zr��E�<�L�<@μ���<@s�<{H=� <N\+�Qz�<1�<������&�2�w=�f�<��S�V�߅���.��x&=<p-=��<t�t:�����i�h&=�js</=���"=��*=(�=����"o��7"�\8;�^	��m�	r=tِ9�ؗ�0�9=JB=��Y�y�E=�X�<b� <wx<?'�<�<i�p�5���<���<OJ�;���{1�;��ԹD���f=D���Ü�,�[�����gb=LɼB�z<,���s	=~�
�$Z��Z������G�;��/�+�i�$Z�<
)i��r�;��;8��<�	-=e�D��E2�j���R=��;j���
7h���E�2����O!=/����_�'����ɼܣ�M�ڼb���T���<A���T�<x��蠚��&{<�*=w�<Ǘ�<O�E�d
_����<c=��H�"��T/����Pu=�lƼBs=����h���ぱ�=�=v#��w�a<x�Z�K��#���x��5���Հ�=a�p�2�	�5<��<���+�S��y��'T=����MqN�O��<F��<w�Y=�Լ�%L��g�9]E�<x�H;w&�<���<�J�<>�<A>C�2�L�Xp=��e����c��'�;?*p�x�(=P���/�48�<�<���<)@�� =� 	��fI=���4��<7�)=��=]<�:�[���A=��_;-�a�G
P�0OB�g>=f?;���ּ�c��M�<���<R����ɼA`|<7�<�~=��!=2�%���L��T=<�3����Ѓ���\�:����v�<��W=��=�ۼh^޼af��ug��.k<������M�0ձ�-0Һ��c��=��=j�ɼ+fG��I=i�N�4���S̼d1�<&�=�b�:�KG<�}�;*"���S=M6(=�3�A�'�������=��ʼXMV=�7�<̄Ҽ/�0�칚���<�r��F�;��2�/�Y�'P�Jna;�#�;5�#=W�<	[=�/�<{�m��2�����7��;��B�b�{<'���W�_��C�N�m���r��a-�Z!U�oD<�{=�V"<a.��ۼ9�m�Ҽ%�?��: f�<.�A<�
ҼW��<�b����?=�Ŗ��kA��r���g`�d9	�&.Z<V��<|���m�������J�qoǺL/a<��)=w6)=�OɻL��G��� F����<�|'��]�"3<�M_�~��ҍ��ե�=v7=�<t��ϓ<D���"��g=�}�;XZ-�e2���ߩ����<��E=��+�����&3��:��%
����K2R���Z�����b�<���=pN�<��<>WL=d��P�>�����[���t=�б�TE%�7ɼ�`,=q|���G;�O�<��%=�A=��I=i�<8�9=Z���U8�<	,���1?�QKA=��,=��.�+d5=b,^�}gH�QL<����;���L��q]�U���Ω<�������`�=e@�hj���}�;�]�;G;�D������<A���2�<��'=<�;ǝ=���<��[�v\�;�����9L��,=vv�<�*�z�ϼ'@�E�M=�,-=J*<=fM'�p4M=����⺼�n=z3���=�*=�n;�\Ks�z�<��<.�<?�
�N�e��.=9XN=���<�3ڼ��r;�K�<]2�����f�N4#���<bTF�zy*=a���,F<���</=�<�Z{�>[Ӽ��&=F
���U��o��!��U=�����/����=|Q����=� �<�����B���^|�����j����W�	�=D�LL.�c0=(�����u�jU=%�R=6u�£7=��=�/׼<+�<�w�;kCX�P0 <�ݟ:�<��<q0���8r�6��;%�/��Y�e�0��E=��C<F �<C=OE@��t�>ʆ<�ۼQ��;�g�<0 @= m���r���r=ۓl�0����U(<o����-2:�'#=��=�6z����<�t9=��<�����P'��+�<�1ܼT�=yn7�q��<�=e�.��Ļv�h��IV=��T�������<d�<b57��*������z�O��<ȋL���#=�G<'�:��a@=��<� b���e=�@d�>��<f�=a�n�޿�mY�'5^��@=#����I�{6��vS=D�/�+����G=�!�Jh=i�=�m=��ɂ=��P=זm�Q`��t�"<!=W�}�M�+���6�87<�|��<����r�����<���<FV��N�=�¯<���<��j=�p�<�;�>ͺ��e�6;5�G�s�O�<�G<%�;=צ<�[��sH���5=�?=���dᘼ�|;p�<�M��U$���=���;T�]�"n%=�;��d�}�T~�<d�̼�@�3����;h�b<8�<\ڼ.:l�!s�<�M=�������Z�VSV�B=Q$��<�6�<�Ǽ�0��O�G2�5�=�h[=�T�B3�,�=>)S=�_g=���;e�:��9�°�<T��=n��,�ϼ�9����&��&5=��`=�mq�<�B=���<)6#�����~��O��<�,>����j_��;�<�褼mN���><�=�<�2=w��<g�}R5=7.�<T�e��>����-*��X�<ؚ6���׼�[��O�� L<�߼�_�<V�=9@����<�"=�j\=M�G=C�*�1�x2�<��:==�<K`��@�d �<��:����;0=�*�oC���==�����'�4
=�Wm��;�=��=��q=�#=Ը1=ũ�<��b=)m;y���<�����S[�
$R����[��;H	J���_=�$=�1*��!�і��@����<_	��a��x$<��i=V�T��Ha=�#w���g�JME<xڋ��H=r��;B
��Zp��u=~ټ�	�m=.��<��:��<��ӻ�<c�S�M��C�P�;���;خ7=|�n;�7���R|�;���d�����lP�'`j�5,=�==}=o2(�W��< J���;�z�<g(��7�<��-=Zc�<���a<�%�<�<�9=eRh���&�p���Ql�<8�^=(�!=��~9���O�k����e<��̼�v=�ߚ���3=�y��[(=�ZԼ�ҳ;�(p���"=BO(=!��p���P\��21�b������=��E=0t���=9̐��P�<�'=o�X��v<�����9=�<�~ؼ�.<5IP=�\�j�<!B�T��`�WL�<\��<7Z�<@��I{ϼS��({�;��h=M��<��<3@�<�jK=�=伦R=a(!�ݷ3=`4�<p#F;��8=V�	=�x<�=<�V2�J�˼�>�+6L=�]9=�Nm=�RռM|f;!� ����<�C��NP�<Y{+��1=��lTG=(�;κ�8Yt�8�<�y�<��B=8���q�5�.H�<�_,=��"�.<��:��j��={�=*s�;zN�����h��x�
<��<Q��<��;tS�����V=���<�$�;��B��ڑ<������tY;P����uD=	��:<+�<X� =��=&!����<�x��vC=\�9����G=^�\�"���w q��QO�"��8Q��5���=���|߼�;n'��m�ʘ�<��z;�̻��߼���<ڑ=��>=����EH=�'<����E�=L��<���<�Z=V�P�[s"���{;�T�<�Ε<۾�<�: ���_=����&�T�=���<�(��Y�M<��N�P?�������<͑8��s�;�=���<w�3��&;����=��=(�=�G�:��ȼ��M�[R=�'9��M=sɸ<`�=��s<􇻾�=Ī,=�U�=i��;I�+�	k7���跀<��>�M�<���<��j�<
.�j/�<BL=��7=�3)��+e��黊��;���<vI=���<z����<x$����L;�΁
<�N��au��3&��%u��nU��\���F��9�<=wT=��<"J	=U'A������*�.�5=9��=#�<}_,=z�=���<�$����<�.:=݃u<ȁ�<f|Ǽ�l�����P�y=��=�co��~U=��"�I��<z-=� J��Fi<�e/��,};5�;�A=��e;m����<��<t�3=�@��;U��<�X�<Ew69�Ӷ�+�������aTI=���6�y�N%L�ջ�<o����n��;������M��Լľ�<l��<u@=U�;�wϼ�_=!&��DS����O=G���C�:J�5<eǲ<��N�.���><Gnj�M1"=M��������-=��üμ<V�[��_�<�I!<�()�4���ż��=���;����no������W�4��ڡ�5<|���vt)<�gR<9��k�{��y&=}e=]�B��4��b�0����<R��dG<i���߼�L�<H[\=\�g,<�Mw�}8 ����?����;^�)=)6h�O�f��<����=����5<K~[=�<�d��z����<X�E=Y��;/c��%�O����<8=�FR=��r<r���Ǚ<S2=7��<ltf�T�;�<�I���<=ዻ����~����+U�a	����t��m=#<TC=l�a<m�=�<�,�<����,q7=�7��bc?��X*:��]<�'<�Ě�b}D=�Z�<�Ҁ��`=$:�����μ��F�P�%<J=&u���o;�?��D����$���:m���������6<I��;r�=�=��P=?|��ք@�J�&=F$�<.I�,RǼ
�/=)vS�K�f���<\A=���<6绻U˫��|���?��p�/	��������<�5o=����h�U�ǼI�P��Ū<���ڻ�<���H�b=�,K<}J���W�� ?=���g	k=n�3��ɂ�s�`�9fC=�f��E׻F�������o=+\޼z�==L����0T=�4��F���7���_=!�h�W���n�#<��<*��<:�U���=u>a�8ϼFQ"<����n��_I�������-=J�"<]�=���<����A��F�<�y�F�;-��=�\ < ᄼ��F=��!�/_=�B=��(���;`�*����sP;�у<X_r�+���Ӽ��j�7r̼x���dR<3L�V��Yts;GK�V��܈4����)h�<�l2<�'=I�<N#��?UA�Rn/=�*ٻx_�G�7��(.=P���V=�od=e�*=��X=����1�=)ۼ��u����<_����`��A�'<C�<�q�ྤ;/⢼y*�l�H=~�<;�����ؼ�ݼ,�Ժ�,q<�<s=��@�$>e;��z<X�+=^)9�T��<���<@�|��nJ�Ÿf<b�<�G=/E=6�=���𐱼e8(=��;S`;D��઼�����\���	��!�<�3=��ܼ�3�!��8W孺ğN=m������o'=��/=6҅�6=���<@����&?=���B������1��<�0�=��=���<��8<�H�<:kQ=/J�eX*�{�O=�u==&�4=R[��aF=�9�<c�=��V��/��^ƛ<4��<�A-=�oû���Q��<�Z߼�&�HWN=b�R�8]��Q�#�U���)��2?=�E�-C�<�/�<��>�)��<�Ů�騜=�\<�<���b�M_2=&����3=Z�7<ϧ�<J =	fn�#��������=&ځ�R�t=D�Y=9&�R���	��p�ۻܼ���*j���<[|�<toL��Q ��L�<+T_�n�<�C6�cI�;�aK��K��~];�_2�~���:�Z��Y7�<�X+���!<���&=�����JX��,3����=�)��Ř����	����<��1�3�7=BD��Ƞ�<���g��<�`��4�<ғ9�Xz���<�>��R�����</2�(�:=Rg�Nu>=yGC=�m)=���<g6��Nw<r2+=2=K[=#���"N� ==�%�:%��;R)�;a�9�J��xb=�/=Z+�<1���!T&='o�"'=��;�t�<�xS<�4=�9����BE_��7�5�=9��<瞅�=�Q��{�:���x��:腃<˫��!�f��{�<��lOR�V��0��;�~�U����M��1���'�;�%=��=9��<*���6d;����'����<c\=��V4;�*$=�r7=a�q=$�ƻu�<�2���VF���1=���<���<PN<҂Ǽ�����e=*�Q�]�h;t�E���<dy��@���X=(<W�ۼCB�<F�／�P=�w��<B�Y=<C#�GCX=1|R=:�=��P=f�"�n��^�=)�<L�`=��[��)�:�"��6�	�i\v�V:�<�o_<7�g=��|���3=�^��F�ּ{�61H=��v=�q;Eك<hw�<�L�����=��켫��;K�Q<�r�;�!W�BLe�9 �"��<9�����>���/g�<��������1�b��< �>�}��<�3	�sx=M��;�>�;����>I�������]�zM�<H��:���<�
���&�d��:�v;�i��y?�<U�=���ΈѼ�+�<�U�A#�<i�R=��:<r9=e���7=�><�Q=�s��y�<��J�6؍�)2��;hQ���H<�D�;����=��q�|$6����7�p=+�>=��_�$�3��p�;i��<-��`B=��<���;f<_�u�K���\�𔚼"�Z��<Ёܼj{�=�S�s�h'=�]�<��P=",<��	=1�y�s
�;U��<�u�<u|����dF���J<I;�;��=���N� ��</-H=򲡽��<�V@=�΋:�`B���;�7=�\9='������;�=�yŸ��=�"=}�,��]���<�T��.\ �g��<R���;�<�c�<��:��n��2�<m�����&?Լ�6s�J��f��H&���5�Ը�<�{���=����XY=F� �xH;dIQ=U�	=���]��<�$��'�<C�<_�=.�"=��Q<ϙ����$<��׼^qy=���(�=[�T�y]i;���� �;�?��j&�9���È��$�k�=W�<�e�����<�w�~eM=��=�A=���<��Z�CX<Y)O=L�!=V��<��H==��0l��=�ͅ��A�<��<��=����GV�g�q���@�=���������#����<�=C�Z=�I=A-��N)� I�<�f1=a���bs�<�D�mм�޵<�tF=�S��Q�<��+;��=ɤ�;��<=9H�����7,<N=�4�I��}�Ƽ��4=�ǡ<���<��=٩
=Gaq�P9o���<[�-�%!�;�r����������m�SP=tב<+\A<��K�7�<�y=�m=�]:=Jq�<r��#=��P��3_=�պ�tq=��_�<�	=�Ud��%=��k=�c�<t�f=��t=��<�����TڼEDF��u�<4�$<#<T��{=ǁ)��G���n��]_<ғ��~R=�'���T��o��{Cc=2 ���7��뗼k׼3?�X�
=a>ؼ�F�zg=�0ۼ	m
<E��|���	cs���1=d�-=nR�V��8�<���cij���m=�{n�U�=P��<�S��iC���޼��F=���;�;`z"=ѼT��<��=΂�<%�_���"�=Z��@�Z�T�<������<+_��/���zCZ=H<<�ld=�-l=U�G�u�ĕ����L�f:��B/�jK=閣�].�<~���<
״<��E=�=ת= ��<HG=؆���ټ��(=l�,�_܀<q	��J�<������.��h<��X=�����L�,ۦ<�St=��Ӽf��<�W=�"=<��.=�O���j�����<W�F=�-�<<��j��=y��t=�=8n;��5='�E=������;>P�<����R����;�<�hF<m-�<�x��%>=�ZX9J!0=�5���E�uD;p���Bѻ疹�wGM���<Nux��!��=�J=n��<	w3�J��<�]�<8�3=��)= 4��Qj*�5J�%C^���&��|d=�H���j���X���<1��n)�<d0y=cV���[�/f=}��!�R����<��T=zRg=A]*=࿀=*��bc�<Փ��d�"=�=`=6\=�D=�7='�<H2=����Tռ:V����H�ma#���t�=;f=W�C<�Q�<=ą<l ���f��ܼye<��༴�<e3�<�.G���F�/{��=�d:��=<�;=�su���==	��<f��J#B=x�F=&���n�'=k=k����J�o�;��;J��;n�/�fJ�כ�Rn�<��d��:o�������L=��<���<�c/<�~���0�����:[�wvu��q�H�T��u^���E�+�0�Լ��;=J^<�~�;
�D��[=J&
�����
�=H�1���ڻ��<�h��f��;�O�<b�N�؁=���t���ſ<��W�\��<�<�B�I�vϩ����P�-�d 4��ְ���;<����'=��E��Ώ<����<��)�%e�z���s�*�1���Ϛ��	�:|LJ=�"�f�J��T<D�z<�F¼�,�� u�;��׺����u�5�X�һ��r9=�xd=�3��X{&=�����=��</L�<9�;�D9�Z)=��Y=�'8=�~=0�^��8�<GS�Z8O=�:=ilJ�R�P=�36<���v��W=��;�bG»b�,=ڒ<�h�G��<eӼU0���7��/
���Z=0�=�M���<'"�W�=�n<�ꅼ�����<f	=�0�B�Z�����u�;"�A=�ң<&���w�V����F�<X5�<�J5=�2��ؾ<�:=s붼Lo(=	dE=S�`=���;�T�VP=��<[(üʻ�<����q١;�,��<M�"�<�C�F����<h�(<��=��λ�����
�f��;<+��	ؼ��x=�L.=�7c�n�,��|�B�A<b�v=i�G��_2����<b�	��؈�d�<��5=�N�'�Z=�h��mq<gx�Ĺ@=a�=�d�<���<����
`�w���g	t�s��<��s�9	=�$?<*E.���r�+�u����{�W�J$�<��;j�м���<h�=�y<��T<R>_=��ȼ�#�T
�<�Z==�?��8_�H=d�U�6G��=Z��N2<��c=� <�����Z;�c����ؼ�M<�,<�qH�ӡ#=j��<�_�Hi6=�b=i����O=�+�|	4���^�:�Ln<2C�� ���"�<�O�	w��_�+��S!=C�b;������N�F�5���4�դU�K�<$:���<�����<�B=�`>�^?��=bG���VB=�0=�)f���<BE�<��u�����M�����<R2��S�vX��UR4���<?�7=غ�<J�B����TO�<�v
<�Eͼ���X������U�;a�	=���J����u=��=l4H�Q�Y=W60=��B����ټ�M�����<X��=	Y=��0�iH�;梴<^0G;��<n5�:s�<^��<g�K�?[@=��:ܭO����<8 ;�MG;�kR=�t�< :D=�����X8=�<\��ڊ3�am�;j׻=S��FI��t<��<�a���8=W�1=���<�;��j�"=,OT<>���'4��"<�ML�� �<|����V)����&o�j�o��kY�;!��<�Ѽ�=_�J=4�������M-=�R=_'�:q�=�=�=�q�<H��<�๻�%]��m6;]��<(�O���z=W]�+5�_�n=,���mV�ʷ�����ʼ�<=B���+<����r�Es��qC��ć�f��;���<�5�<�����#=;IU���J=(�"�n�AɄ<U�<�kV�%�<0���:����O	���޼��7=|R�<1r5����<R_�<&���*��;����$=�)_��Χ<�U,���h��[�z㌼u�(�E��sA=����!��<�-�r �6E=������y��~x�<υj<��K��#���Z���=C�<)�j���<\���Q=��<�j�<'P�Q��<�ʻ9&=0Fa�a=�l�;s�=7�}<�m�=��ż��I=�(�b����|@=n�=��L�FT=��<*P=�B�<�}���I��6����<	C{�������7,�<Mj=������U=T��5_�<:=��=�=�BX=ZNȼ�Q�<����8�<l'<<��<N�>=Nl =��ͼQ=�R=|�*=�`<����E�+H��+r9i�<�o��@[=ϴ�:��]=�
t;˚�9!n�<��<��R;!�j�1��0�»�_=ַ�3�?ˀ=Y��<�;=2���e�n���<aS�?�(���D��"��q-��x����oD=-е;�O@;��=hi�<ҝ�<��Y��V?=�T��}吼x.�<�"<�Y=7\�4�<��
����<M�_=;����K���9%m=�:<�b�jz���Q=�J��8��p*�<�yh<��T�����r��;�<]&=��<�����M=�`=�k�<��w<B)��Z�z�s<��N�=�t=�,j����<���;��2����$=]m�<|��<O�Ҽ�=��&=�b����<`��<Ӣܼ��=vͼ��x=�TS=�#E=Y�'�t:��2��tB���=.0�$c<�:��\-��:��;KW5=�"?��a��=�:�Oa<�>�=#�<�sh������Ǽ.�:��Ӽ��:=^!g�OFܼ�P
�AC�d�?=WuW���Q=+F���4 �5?�O^�<�L<���;�D绕�;BZ�=މ<>��;V5� �<�^�<�%�<���s���瘹�]��ؠ��=�R���4=҉c=`rX=|H=��Q=0��:<�.=	�;�G�FO�&��8�/�;�g����<_�<�j�%\=��K<zC��-Mt��B1�^C� X�< O�>\��u�)�EQa<�~���h=�i?�0�$�M����3=�^=�Q5=�)#�;�i;fA=B�.=�(�<�p3=��<Κ;\T߹(�J����
�y%������<��*=� <��%=u�:��2;49U�>�4�r�a<.:v<*�<��F=ş	=j*��7&�<N���K֧��(<��e��5X�w���M�m=\�I��|�;+�V�t.�<rL=C5
��5���4�rxX=��m<� =َ?�c=����<�7Ƽq�<����tмX�S��%(=�B��
;�<K�D<��<��}��<��$��.�B\<C=�Q�<l7C=	�n�6=��=V�=�왼��<�U����<B�xT���&Ȫ<e�P��R����+@+���J=+�=޿���V^=��<'l˻��5==ݛ<�C=<\=H=�.�<�E�<�"��pp��[�1����<�cJ�h��s�컚;�:�Ӽ��9=E��4W=�%=��jҀ����S>=��༏�����c=B��<%JW=�k��h�4ѱ/=\*(��;�<��t�>�����MS1�F��;<�0�N�;�j&=���;�N/�o{���;�T=U�F���ļ6c=�:�<��{==O}=F1�T�y="�#���q�b �<Gw���4�$���\?=a�\<��Y<o1=T�t=��=�ʼ0�<���;�{|�e�=��u�y�z�3g��s��V_4�K�G�$;μT�Q=�8�>�<�Y<ݻ)<�9ۼ�V?�Ps<��,<a=V���H�ռ�y�a�|�����<����@��='��<O����i@���=�<������/��<[�:�ż&m���w�6ڼ���<� �#�<$��<q�;�^��\MG��J=Z���k�3��<�Ѩ���_��qR�y�
���U=&8�W�c=����Ƙ�VE���������f=~I������<"����=�;l<�)(=����u���K4=d��<�fY= H<E����\N=�m��Dt�<�ս���c=�^�NDX=�.5<����T=y�J<�0V<�3��!�v�}���λB���(�b=�kU<s�{z	���Gl�<-=��:��]��I��(=���������3���P<��=��B=Q�F��m�;�>=�O�G����J��|(���:�ļ�N�<��/�>���j�ӵIB=��<ȝ}≠`=Yx�<�@ļ2��<��)�����6�k�7=�
X�f���9=�N���h1�Ƈ;�l=�P!�"��<pw;��<����g7	�<9=�ĺ<�,���}��/}-=K)c=@&�<n��1�)�kV�{26<���;�gϼ�d-=�m����<s��<Io��_Lz<�L�C�3�+51=	R�������Kj=��J=��=_�5=�%p;��J�O�����غd�<�i�<aֹ��N�,�*<,���cA=��Ҽl���L=j�P=��<9��;�_�-��;��G<p��Yၽk'$��)��d����Q<����6�Y��<��<�i�;g`޼�5^�_�<���<2�`�j��
o��S"��U����<�o<f��<�@��M����KE=�����ԛ<L��:"�[���ջ<���;���<��=N�=��u�و����<�>+��@7;2��<�&�<]G�5��<��V�q�=�����;v�=-��<إ�<]�9П�<�@=9FӼ��|�9�ϼɋ���=>�<�!��;*S�;Cܘ��9L��� =��X=5��� K<=nq%������N�4�<{�0��;ׄ�<�_L=�=;Z=-y�<~���J^����<�w�<�̀�ዽ�m�<r�)������r/=Q���{r=�?I=��;��	=��=��
��f;����P=�RV�*�<�LL��.>=�	���#=�K�4�P�1�<Q���{��;���<Yi�<���ӳ/=��̼����G�=&�E=q���NX�;I��<4��;X��;�6�<��=-=h�,�<=;�;����6�����~<�ҙ=EB=>=�ak���O��b<��T���N;�\X�f�W;	u8<HP=Q��<Z;�<]=W�<`=l=�м𩕹[��<�*P�)s!=�� ;Mo���ໝx�Ts��G�<��,=��Y=z�q�>K =��<�#P�wZ8����<Ǽ�T'»(�(;Z-�E�/����.P�<^͈=�_��z|=TX����<����Cjo<�P+9ֻ�y�<���<��<�X<E�L���v;�ү�`�x<U��2$�;�	-�D�O<1�:�p$��U�<��8���<��<~�\�}܅��Z=PMw�)�̼�+���n�=
�4�������I=�!=-��<�������޼?��<ǗP����~��:�Dg=��<��J�d�<~B������v/=�e�<�3=�%�����<�=�����=n����ݻS�{��H�<<�<$���)=�tt<�TY<@Δ��� :R��λ�< �����s=n�=Y�g���j;�.�<�r<�E=S�=Vk���)輖a=� i=��; C���U<���9=��<��l���=W�Ǽ�W��+�<<�"$�g Ҽ ==��47�<��󼭣K������\��1@��IN�c�&���m<�<vY�<�=��X�%��:�}%="�D�qv+��!�s��<
�P��[=�t���Q=����a9��<�w<:�<�"=ɹ�<���P�.<*)��_�<@����%j�ZE� �;b�=*��j�3=�H9��B=q�7��+P��{<a�!��5<;<'�N�Gq����� � ���~9��=�E=�ܔ�%C��׼d=4<C�0�6�<���;,A��>�j���	�º�<h�!�9(=����=�	�<tiC=��=;	�,=j��(�S=�������4���<�9=��O=>#=�B�W�R=N����m=����tI@�gA5�D�:o��<�qH<���<�����
Ƽ�`=�	�1=�_˻9zl=����=��5=�y��Qq�;�s:=�ݰ<�;A=x�*���>��9�<��μ��'=�D��H�y��]�1��J���k�o�{#�)A�<(�}:�>�/�<��7=Y����&Ǽ˅�<"�����<#��<��E='E=�K�����?F���R<���<��߼Վ��C�=��<h�u��ٻ�[��+�/=��%=�XӼ� �<*�:��R�0�<�Rۼ稭�<L<��`;��<^�r=9��YN<�f=qV=���<�|�)n�]�=�� <J_,=��o���<9s���ܤ���"��O]���+<�%�Ȯ�;.
�<j�<��7��į���D��x9=TH=H2�?�7��η<Lr���%=;��Y=��e�=�o�<��:���<��켁�=cAx�"3p=2E=���<Ť3=V0k�7}һʥ��?� =R3M���H=購�0:��:,	-��V{���=O�3��o����<���<L^��\�<v>:;�$��<]�<.��2_=�f�;�KB�-�k��pm=�'�� N��=����է!=H�p�^� <�ì�t�Y=K��|L=�F<�89��_-���œq=�d�Z6<�7=u�=�s�:�  =��<��-=ND�<�!���</,G:."�<#�;�3�(��5�<\� =z�'��F�<-gg=7�;��0=�R�=�`=[Ui;��<�Ѽ�!� ���K�<IV���E��\&�	M�<\�?<	�N�i"z<p/;��r���a=��K=��<���<r��|Ⱥ�6mW;�X�>�=V)|<�/ټ�G\���3����<tՈ<�P�<���;�<�f�s�b�[�M<�,w�+d�<�_==�S=��D=����n�li�<��`=��a=d���Vλ<�N���K=V$���T<�t1��N�<E�
=}��H둼~�9;.yM=C�ʂ�<�=4ﻼ-�Ի��<?1:����<�^]=��M=��=DC�����y��<QG=h�l=��d��8�^S@=qb4��T=�Ӱ�U׺mjM:�Z=_�[���!����'�a��:h�<���[�Q���շ�J���<��#�g��<��0=��h��Y�M����*=����̉��A���ຽ��<�%��.���&O=�Ӳ���#�1�x%D=1��<;P8�p�y=�ʳ<F6���)ڼ�:�;�Ay<� ���x=1�#<ס��
2U�%|�<I��x]<w�&<+<^@=�F;Z��<�'6�gym���O='�v=Sa��C=������1�k��}=��<�/F=v�<��Z=b��<G����g�A=��=�Tѻ2���?~ =��k=� �M֫;wV=Cl���m,�f��<��=���,��k�*=E֭�3<�QQ=7�:�n���=����擼�'��8$�Q��<��`=�3=���<�x�����vD=���<w=8s)=�%���<���|�I<�D<9�Z;s�7=��S=�� <�2H���}�%'=��E=0B%�ļ���=�zf��ۻ�?3=͒�<�89ֻ����:� ;û�<�DP=��
���b<¼5��o�<^�<Q��:��;��<gѐ��k��B���=�����`=�ê<�t����=�R�=�6C� (�4U=����9<=�= ���x� �}�%="�w;,|��[�<�^�<��0��<<�cn;��<z��^��g����M�7�E�����J=��κ�T ��^�<��༓�q���`�X�=�%�.����<~x�<x@�7?U=HS¼�k��L=*d�L��<�`T�l��;È���U�:�����d>��ց� JV=-]9��$0����<��`=�7g<[�X<?�<�Xɼ���<�N�<m�C=�j��ޒv�m3<u��Y�¼[?3�s{���=��=Ҫ�<מ)=iO�<�qL��$üBc�]��<��ż��=�6\��<�<UE׻��<�K$=:?�<�
$�=�s��ۼ=����>�X;�<��-=4����W=q�;^�<�+ݻ�	�6�<x(	���=4=A�T=���<�6=g�	=���<;=��|�0��m�9�6=�	*=�8�o�=k��;�H��x=���<H�<�V=�oO�����zz�1�$��9���<A=:����<V�i=�ㄽ�k���S�
=���<���<<�����V<&D���C�;#V��������h����_4���)<��(<�nͼ���;[���W̃�#$p��3N<z����n=���ysR<�U�<2�P<��(;����*	��*�]=X�J��5Q=��J����@ry��Z=�몼S�V=���<,Y�J?'=Q�=6P�<XԔ�aE[=P�T�	�ɼ�]=<dʻ�q���ƻ����l����m�=) +��u[;�ź�\
=����T@=�:Z�+P�<WX=�d�;�W���Q<�m=�|1��s������=��8<_=�=�<��<ϲ<b*�<+�1=��<<5����=-�<PM��5�&
=�w�<(=EzX��ߋ;���<ݬ�������ڻ|�ü|��,�n���m���\=I@�;!�<��\��
�<V?=���=��=�k���Q ;�Z����<�.G<&��<�\�w�߼FQ��j$���,��)����6���f=(=F�=�!�:<���;��]�Xة9@P�o�u#�JD4;���<2W��o��S�Z�z���#=���uvK���=�x=��u<,"p=#��<6�,=?H�$4
� �P�=�o�� �:];ɶT=~�<�@�;�������<�\&��]�;*导����z�!�n���b =�k�<$'=�;��0�<�U$=��ƻ%����E<;lT���,��O/��I�<�E =L��<`~=�q=z�<
����
�=ڊ�<�*�<љ��E<���RaQ<!��<p�i�:<�������/_=�b<��z<G=w=w�
=�,�>\�6���k��;���r=ޚV=x�i=�G>�ӳ�N��;����*�>=n��;i�=7����d���<	]��ϟ��Ο<��g=Cc=���<�G2='�I��g�<>�˼�&�;.?������=��J���<<i��(P�0j!��mӻv��f�} $���<�>=	���D�;$%E:R���ۻo[*=e#�<.e�<#����s;Ĭ=<,7��;<��<k0
<C̻�I��uy��)�<�= j����<&w�����,\ �34=���<���<���F�`����<�D���B=Ժ���#=V$���<��v
��Bi�<B�8=��]=�mL=�T=)
�:�[Ǽ����=�l��a��;N��5����<3��<�B=��{=�3�z|d���~<�|<d�1����<r:���TټФk=�{���+T���;9����Y����Ӻ�L4<�=����"�n���2`=�D=\���C��G�
=mKw�'J��}$=:=�Wr=�K%=�x$=~^����<?�<vM�<���<h�&���*��D�<c@����89%��� =G�'<�� �[��<I�p=w	�V?;�E��~���v=�$�<�̒:T�<\�_=�rn�����s�<��=�x=":?��Z��i=�⑼���rW=Tr�<��<7�=>mt�_W�)B�:J�)����<rW�{_�9l��j�u<�=�WR��	=n<��ƻ:��<�m<�=I7@�p��<�0J<}.=�Z��f��]+����,���׼��W��ͷ<0�V<�����!�;��1�g�X=�F���һ+D=ؚU���r=�z'�m	�)�üż�<ʚ���=��=݁Ҽ؁-=�f�<葕;��J=B�9=�B��l_���4�������<���;��>p�=�g��F��E�<1�)<���<�������O=>��<i�);�X���T!���1=K�߼4���9;C�&=�L0=[Z�1$�<h�=��m�]��=��2=�U:���e<�$�"l<��6+;݄��Qc==s�<A'�����෼��~<|�u=68R=��>=cB�<!�����<=8���H@=�Y�<��Q���<鰒����|Q�W�H���<�� c��}�<�� �ێ=S!c<,;6�Y���2?;�|;�j��<VE�����<f<z���<��T�G�<�!=��L<��:=��$=����4O��[�;��O��_�;��<�7��Q��'$]={
=�l1=,Xb:�ݢ:�cT<	e⼺'%�R=ș��f_��wm��=���<n�y�7�;�_=�J����֚d<��O�P%<���gY��?�<%^���~�2�+=���<��<w|�;�����i�<ixB���=�`�h=݂�<��:�8�$�=%@=:,Y=�̎;��=�\=aP��<=ޗ/���ȼ6|%��'N��H��6j=�=;���)�T�x���ى<#�4���)=jEf<=�"��q(=Ѝ=C�R=���<ɈN=��9=����sKF:�3=a�5=��<���Pߖ�I��Ӭ�<8�߼]��<	x[�;=���<��9=�<�;=��<AA�<�}�;��C�?7]���!F7=��z=o�;l,�	�*�@���?�*=?�$��
=��.R���8=���;������);4Q�)K������)��26=ͧ�<q��<���(i�{׼��<�2蕽�c;���<��h=��P=�5;e=v*=�A1�ǧ%�»��M=�#7���<u��;ݙ+=� ���o;�ּnK<�\";��h=\��u�
�V�<���<�Ӗ=�ۓ��a=pQ<�{=��㼷���K=���Լ�\ȼ���;l_���}��<=j<`</�D�˰s;1�?=qi�<����t�@�G/��Z�Y=�Ų<��޻�`=�?=�aB=�� �^%]=i����P�HD�Xk=�m2=�g�@Aڼ|NM=���`$�dk=�B$=�0����;af�<n���?�w��,=9�v�،���:�2q<N�=�	K<��r=�}F�ةT�m�9��8��t9��;�<��<����ќE=p�;�0�:��� )7��N<p�0:��l=,��:�h�e��;��r=��=ۂ�<��2��U����<���;��:/��K =�j�q#���\w<_y?���=��D�ꗼ<Pȼ/�=f�� O�<ե+�H+�<t����ü�Y�:���<�ע<*�7=�˕<��:$9��R��A$>=<1к�8=�9M=}�O�ݦ<�J��p=cLa�L�w=�n=6���D��
Zټ���<h!���R�! �A˂�U�GF*=�Mc=���F�ԺQ�S=�H�<.����\<|�ȼv)W=j�;�ְ;kt!���<�e7<!�=M�9�V�=渓�W#�<C�D=?*(�}��<4�*=��:*ۂ�Yј���@���ػr^��?8=)�������?=�p=޺S<�(/=�F�<�]�e�w�=�8:{<*�&�/�e�_<�
�9�E=�zݼ�!B���IQ���:=�?�;s=9���I���-�;�W=3�1=�+i�^Lʼ7;<���<s�=f����EL<���<�D=-tu;c�{=�I=�)=
�,��ء<�P=��Ҽc�@�T�.=GGm��J�8��s<D�}=I�2jܼ^��< I�<-�WtU=�b=��ǻ��<��)=�m���<��,�b1�=;�=��;��=�o�<�ko88�s��K���	=� ��f=y��<�^_<:�d��ܶ�܀=�"=���/m�v˺�O'�u�N<)s"��X4��a�<����8t���Լ�ջ<��1�x��;>d<�e#�-qY�K�T���<�6$: r%=C*���I=��+=SEi=P$��z���2��<4���UH=�<W=�D=�9D��%¼g(��&J�3�ĺo�k�U�众�����<�&��a�<3z��H]=�(=XGO�p�2<�@:��<R��o#����;�����2*�� *�C�.=�4���<vS-���<=�e�aN9���Q��"�<g=�,]<ъ ��>�<��Y�NV+�?��� ���H��-v��~=q� =�g=?��
x��p�V��=�
�=ڟL�Yc0=;j?:p�=r��<C�=�c+=��.=�i=��z��w�<s�T�g�_�w�k���;ƐI�;�M����[7=��Z=�tH=��5��]�<�];�,=+��<Z��'�=; G�;�N�<�9"��`5=��a��_�<`��<��"��5���;nj��fI�Y�N=Y�<ΪQ�;�<2v�<�'=b�><����=1�X=�8=s�U�=J<)j�\�<0��1���(J�\Qﺎ}K=^��;����<+<�M�<(�;��;��j=�=!���*�x��,I�=ݷ=Y2�;;�,=o�=v���|<\�;=��L���=�2�<���<�b�*e��^��x��0b�<�8�<|�<�V4�����Tz:^���4�=O�,��q�;zM=&<��i�dVk�� ��c���=�8��;�[<�sǻs�0=-Ձ<L[��m(<�95�B� �AH=և�<=S+��I:=8�,��N����:P�E;h������N�=�5W;{�!�$E
���`���<=�+=���yEμ+U����x�7��<)�>=�=T��;��r<Q�T��;���O��|]�I>����S9�������b;u�	�_� ���E:;=��9��R=�TU=�o:=��L=M�I�ln�<�=��=C+=F�<ua:�7=����:="B�<��=Ô=��J=���<*=ߋ'�?���T=V ���>E��gk;F�������=����=0�$=���@����]���Ҽ0j<�B]���1����1�;���<CA�<�?<#�P�S�0=@C=0�==�t}��sI=�;�;�3	=l'8��9��#�:��H���B=�S�:EJU��;[=*���Ϛz��G>�O�<�O�z��1\���p����<������{r���<;;jJ���<$8���|���������[=�mA�R�m��)M��)��a<`��<(�i<�=yy��/�B���D�[<�ʠ�����OüOX��u��:��&�>����;��k����
��;�۰<\�c���t=L�O=׵м�j�=���bv�������`�[i#=�m����;2�{=f�=�Pi=�[C=o�:F-�<6�Q�V�b=�V%=ޠ黁5�<;��l=�*�\IZ<��d���=�)����<foD�J,N�J��<�y�<���<��=��=؅7=�	`�^�C����;k�#�S�:�`s���M�E�n�?�:�G��<��*��2�"��WD\��A�<Q�\=���M�
�0w%��a6<��E=v�~�\�p�L׻M��<	�'�^L�<�=��7=��h<� ۼ�4��V=&B!=�W��Gj����T�=ô��8�Լ
%T����6��V=�"5�.=aG�Y⼼��׼;2�<u�T���<���;aB�;�N=	�\<D�8<?#0;kC�����G=�9�< ��$����rۼG��/�<��<rW=G���LZ1�-.=(��<��=q�<�ل<�K�<�4�9�5=aȼz�<�^�<-s<�<��7���"�ٵ =�O<=)��<���3O3=���;J�<��ؼK-=��@��J"=~;�[�6*���C�<�/=��;=ȟ=y#���"=M;=q9;��<��3��a=���/�dG�ۿ�;(Ij;(y
��0�<�������<��߼H�<��=Ū{:�^�;c�<fm��Z�˼w�=ed��YW�<�ż�w =٤O��$R��Q'=���b5]�rN�����W1=<�>O�[�J��@����᲼v��<�`����=�H=�����һ���<�D<��ݼ�#��?=�eu=:_��4&=E�k�����_K��a7��N��qK=J(��rM=>Ng=�*.�=�S��<�|�<#��a��<L�n�HX<����<u�9�Լ|e%���I��n�������hI=��E=�;=��-=0Q��)f��_G=�Q�<�<g��<��D=u�7��s������9��<��#=8T<�׼<�@F�D'v�?�6�;�m�<�%k��/=(�="�w;Eن<\65=�uw��V�<)�':��<v��<���4�<��A���a<=�C��ç<��=v[��)����(=/e=L�[���&<��0��2����<��T<�=��螼<������;n�2��{\<��=��$<r�<�+D����<8R	=f;������!;��
�����!=/je=f��;	6��*=ȁ=�?W�D�p���;�*=T%h��Qg=�~<HM�<d��QK=}�<&!���`����P='�M8�z6���=��<R�#<�_5={l�<�R`�<9λ/�H=�?=���N�(w����Q=��@=N⻷ު<�hм� =�_�������<�T�<�N��l���E<���;8�)�O~;=�
=�����X=Tu=E���{p��&C�?� =V�N���5���<9�=%I�<��=�*N���b�!����&<I�S=��I��>+=��*=5v=+R���N!��)�<��X==x��F�����<��;u�o�q���
1Ի�L���%=zч�ː��c�b�ử3`�d�+=�ȼ1Y���o;Z1P� �ʼ��S���o=���<'9ۻ�-;����ռ.�Q�[Xܼ]	C�	�><�N�<�m�gd����Ǽ���<l����p�&#�-�=���<��E�>M4={�< ���~���y&%=ݬ��b�¬%�����	�\>���z�C}���B=׎>=i�L<�v0<*�v=��<�	=�a%�̴;�&h=��<@9=���;���<�嗼�'=�"|�*ʓ�t$����(=
ư<<�<��e�o:i��i;����53<�?=9,�<�-�</K
�DV�<n�%=>}>��Α=Ա���F�����wἣ$��Z�=�D陼�aT��Y%=�>=���;/+���n���$�<˩/���6�IUżK��;�D*��B��#<>Yk��6�<�=$Ȇ<0R0�J��#u8���g���n<���;�"�|`<'x<��!�7���T&v<J���$W��J�Q�ɞ�</B=�(�3�a=rPμㇶ;~Sc��<}0h��_��ZV���E4�J�?=6*S=�(�<�j=�c��Z5�<i=&;��r<�i��==���<*��;��_=?��K�$�����M<r�Ѽ��U=kQ=��s�_��:�;@
�<���.��<�]߼��
=.,����H�g��<�2^��$D=��<�`�o�=� ;��;�U6�f�i�=�j��~=�f���ӻ�1B����<wf�;ߝ����<�ś��==�HI�sq��;>w����j)=��X�z�<��j=��:��"�s�v�!���`�=�"��ټ*��<�<��G�_;iQ(=��&=a�[�o	<LL��Jd������<f��<@Ϊ��a�<�d�a:%�K�I=P�=�e]���<�S)=�xF=�����=��}��q�<���Z�<Cb�"�2��!�<�r@����;��:=Q��E#N�d���RV<�B?����;acg���<Y��6�d=�Q[���f=Qip���;\z=���\{0=>;!��<:C<�|�^$�<x�\��!=���w;h���=��%:���<� d�e����<��Ư�T 
=�k�;fu%��Y<�V9=z�6=Iъ=XGK<ܢ� ?R=k� =��� �=AF���2=�H5=�{\���<CB1=��Z�F%L��A�)�߼���;�I=���<���<}��<������^��RT<p44�dl�0�2=oi�j =EU�<��M=s��gh+=��1=0(�;��==ެY�঵���G��M=�����;�!=M�==#8�;)�Q�;���<lB=�
���}�f*x<|��;�;�ξ��C;=�ۼ?t=�ý��IH��Լix�;��=��߼4�=�R�:�Z=�Jj�����A=�Rϼ�(c<���ļ�~���U=�  �ntV����o��<���<у
=V;���Ǻ�g�<PH=���;�/"='8�<����-�<����O�E�l;/��Z<��O<�>V�w�G<X�Ǽ��s�#+�R�A�M=h�m<�Cr=�'�<'�=�b��G�><w>���o=k׼�W=�A�Z�=��b�"�><��Y=��<��׼2)��\���;�,��&��~5=���O�re-=d����(P�Դ&=Y;_�#<C��:��E�Fk�Re�| |�a�'��(�<K��<x8���=�lC<㽼=�ֻ��l<Am�<�%Լ#�a��M=�}���<>�%�Q��<r��<�E߼�TB�s������<��l=؁3=� !��W��8ټT���l��5!��f*=>c��2��$���B�<1�$��ȴ��3κ�U��4lS:56�\�{�o��<�Ő<a��I�<tSf�t�ռ5./=��b<�[=(ċ<k+���"3��>%=A=k��a,���!=�#=�	�;�-L=�+;K16=.<���a=�W_�84;4vO<A�ļZK=�j��Ǉw<�T�<�Ϻd3�<���8RU=��=�[<�t!� �:��y;f;�<]�z<�d=���=�@*��0=�.'=���<[���u<[-=R5�:{�'=�h�许<<'��c=�<p�F�4	4���y=��u�;�6<�:��UX��,'=�(����=m̼���X�=�|���Ҽv!?=R�O�6��6���3=�1���|<�V=2�<A.�<@)�<b�=`���'Z=X]�<�￻H�%<��<<)`j���s=���<߿<p�K=v:=����t =67�9Xfk=����M��P8�G�V����:L�-=t�X�T���P����=ko�;�I<�� ��=�'�Gj<��S�0l�X�=sՆ�Bd�����\�U<�zv;��X=��I�j ��}�u=�@���޲;�Ll�=�<�n(�h�&�eo`�0���X�r��<�	^;Նo<��W�/�	=�=W�뎼�F�U
A�	@!�ɬ�]Wy<K༴�=5�B�l����<��#=�*~�)l�<.<<Q噼!w���(d=1"=M~[=��H=�|	����Oe�<�`=d-L��p�<	�#��ũ�<4���7��:�n�L�Z���<��<�2�})�<�KD=k|v��.=���<f�!=�b�<�np=�K�;;m�ٞ���5=�L�cv�<�
�X�<�.D;�屼���<'�Z�yk%=w��;%v=A�����G<����ƞ<V@�."�<vぺ~���8�.�2=��;g锻�����:o/�0�i�87=�r���i����ף<��K�T�3���6=n3��o��zn=ё��m>�:�=�?�<�x/�K���6g=T#Y=ڨ�<�޼|_�a7ʼ����Jڭ<�<��Z�(��<�;�<kx=�ؘ�m��<����Ի�'�#<B�l=$�s��<0���	���`=kґ��[Ƽ�s =�=,�F�(����Mȼ�:T;�l�<;�J�~<��<��[=�b4=�<w9{iL=뷌=��ĸ��{��-�	�W��V�<\�B=�ڼ��=$��:�o<��� �=-��<k߈<a��n0�����������ϻ�֧�c��;���9�ޣ<�!�<�_<=��<w1=!L+<l�j�A�=��7=Ly{<��8=���;h8���J�nR¼|�=�I=�e"=t��np�<]o�f ���_=����[�+�,�T��==ʤ9=��6�T��;��*�<[y�<Tп:�Q�<)e}<�Rx=V�=�K;(}�;WV'=.��9'3�!`��ڼɽ�<"=q=�W�u��<�ļ,�^�sc�$Q�$�A<
ہ=gGK�w8<wǢ<���<�1O��=)>K�J"��_ 1=4�q�S�<#�K=(�*��}�;�-�M����?���
<Ǭ�;��O��z�5/g�h�<��<�<RVW�".U�j����=�>�-��C)=]�*<������K�j="�meE��u<4ـ= `�<�
%=X�[��g��^;1=,=����OC��芻��=�
�<z�%�,��;��;m�"=���,;�3p�}�L�!#=H���?s<�;f=r�Q�?�(=J�8��}-=Y�G<�A<�:<�_*=<T"=Ev�9����?�/��y�C���=�Ȼ*�!���<\D/���5;E<K.�=�<>P�_N���)<�eQ=�%�<bρ<M!�<&H�Y�:=tg3<�����Mr�%ځ=0�=�մ<h�ɼ9͇��o�a��b�!=�ns=`k0=�!T�o�;Ed�L�y<O�#����;+;v�Q1�<�e�<g��Լ�;�@=���x�5�f軻+J���~2������t	<Z��5P�q��=�?=�#=�A�<O��<PQ�g
�=Ӣ���=��?ʼ�"�s��<�:<�k�;�{=����<���s<���<����LH<;�d��[�x=č,=��?�B����2
�׾M=�n=��
==Md��}	�<�żv(=C��7&i�׀=�;V	<nd<O2j�3��<ǯ���=�B�<��<�z0����<�0Q��b��D-��*=��%=�G<�d����,4<Oo6<�o�<4�=�AD��I^<5�^��}꼷/.=
�=pN�<�K��)-;�у<O�;��<Yh��_���<(b<�м<+9w;`B���M=;�E�2`ڼUv�:rT��`E=��<a��k��Tq<��<Re2<��K;�h=D'�=�xW=�7=��+=�@[�
�:���k�W�1<�׼u��<��;�,=Ӑ�����g��쿼�<��-��^�;WZM=��u�kk3��[<�N=�w�<5���<�����I;h|N=�N�<pI>=5/K=nk�<����@gB�,�=S�<�kq<��0<-=RnJ=�����Q=btE�6����=�7�X�<��`=�";j�4<E�g�j=��l�(�<d�_�(<�M��H�������=:�!���F�PW=��:<*���c8=;�8;,$����<?P7��j�<�1���O=tli=8Lj=�"�lt#�VӼ�l��9�="���<�����&=�<���5M<m�v=]c4=9Հ��~伦!<ߝ%��4�c�i=f�n= �S���m; "=RE��ȫ¼Р����<�d��V��<���<�Ճ��U�<Vd���2�<O��������<�A=��<�5�<YNo;��/��A2���.��S���	���1=K��=����==��n����e=$<�C���+@=��&�����<�:�Ƒ��-�=�9�?-=����$�"<�w���߼��;��x<EC�<�0=ZQ�7�(�	_�<�'=a��=b(;=�6�$8<;�༦�==��=(�G=�y�<բҼ��<�F��̮���<�����$9=6���BX�G�m=[(4=|%߻�D=)󬻼�=��"<{<wg����qo��d+=n"�<�	�����m���J���/�k'�SD�;RJJ�%d�P^=����t�u�<���<��5<���s�2=nh=V!=Q��	����:��W=��<�2�mۅ�"S%��<��u������"�v�I�"I=�;镨<r�ļt��<[=��k������b=j��#�"=��d�S��T�;~6༕c�e��<�w�S�x��q�;��W��J=�C��ݰ��k�G=o�!�m_T=TQa=)��y��<��%���R�WQ�z,��W=l�a=A���6=T�<�#�������Y�A����1��J%�gP�<�<���<��T=a�T=�0W=xi���ؒ�ޏ��O�s"=尢<V䒼��=΋/=[�缂�,=\����)=07/���ܼ!Q�;&'q�W�{������=�	���P=�I=�������<����(�̈<0+S�O�<J/=�8��)�}�b�<=�Fj=�O%�YX��i���[(=�~�</�<�dE=�H��̔<�#�E ��뛼�I��w3�VD6�J���S?�<3I)=��5=�ѹ<�s>��Vi=�pW=� ļhm<�24="I��Iُ�9�<zl"�E*��L�<=�v�<∸<!�o�f��<Q��= �=-_�<�5/��o�<X��<X<��/;f �<�g=qtV=<_<=��j~��ѣ���G=K������8��J��<��<_�	�G6��ϻ�� ��@=���<~W�#���i���)��җ!��ǟ��� =�պe�"��!8=�>,�4�`����<fr3�X����2����}M*;݂1��3(��%V=#5�1��B{=hT��*�<P ���4��G˼�c�{`
�J=���i:�=2�}<��_��+�iݔ�@>��y7<!0=H�H�Ga ����6UC<؍��)C��&�<4�o�u7�<:;=#�=�濼��d<�����9P��P�{�X�;e�<8t��c��<@Oú��\=��Ⱥ��3=��o��A=T��=��!�(;�<x����v��7�<�A��:��o꼀F��&C=/W���F�L�=��#���`=��!:e{����m� ��:Bf=񲍼�s&���y�1��������o� !�<�(漛H�<3�n<���� ��<�0-��-=\ul���B=��<�5���g�;�=���t��?�<t��<6��<E�l=���;aTc;d$��Qt=�g1=0�=����;/������T<]��='+�=��*=��-��@+�� �A!<=��[;��<����c)C=Y{=k9!�R���� =Co=Gv�<�Ne�����,��<�=
�c����/��1,=B�<�$��*^.��5?=<� ��6���Q=�홻o��a�zk����<E(d=0{'<;=�|�p���*���=�pK�����=�<�
I�a��<R=mS��(Z;�f��Lˀ���d�=���<ɋH=-�=ƹ�<>?�;���<�x��h�����<rS��0	>��(�<�C=k��;}H���@�;α5��@$=Y�:=<P;^�`��ۻ<8�b� TN=�*�;,)G;��üM�;)7<S)
�P��<K��;�齼��J�h��Ѽ�<�Dz;�R���;<��κD��u!������L��U=����	�<� =���=�$����3�4x�3(<b�"=_aV�����d����F<(���K�<�~3=��.��<��<�S���^�|{=�<<=a��Dz��PZx=�	����b=�dD=*I���H�<{\8<�v'<:II=y���/��H�����/^6=�;7�5��F��5����S=9X��TW=M�3=�?,=�z�<���;C�;~K*� !�uC�=�B�7ka�(c��������R�{h@;�[�<S�=�@5<Sn+�]=߼�~<���K�Keu<5�
=-.��;���X��u�aA���l3��
=\�1�)�ɻU�<��a�o�R���<ذ�<�;2�LT�g�����;C~�<_L�<�=��l:k����鐻=u�؇(=�c����B�L��<�%��N=}�IK=�6&����;}�8����<:B�<\y`����<�|ռ��<��F�L�=d�}=�Z=�o=���<�����
�"?�����;��Ʀ��Oj���:Ӥ��Z�=�X=vh =����ó=>%����6����Xq=�<�ۼ-w�<�ټr-����	�tշ:e\���I�<҂�#�;�b��o�S����<jy��R�0��3=�NA=��)=p-L=��=�[;���q7��	�;��<a��O�s�a�ȻȻd�W��47=��2=��I<�g=Vq|�徬<$Q�3k��� �61=:�)�4<D��|I��O==���g���1����(�;mǼ�IB�F�)=��6=�te=34���-a��0��]Z���6-�<�΅��	:U�%=�;���c�:�#=*\7;�㤻�+g<�H�:��U�z�<s�(=��%�˽ �;L�;� ��Y�6��U�i=��ܼ���<$}_=��!�U�5�K9=Y��3U���@;�$�K��<�\˻QǑ</+ȼ���R�ؼ����d5˻\�<Q��<Ug뼖@`=Z�$�\3�<jĒ����+@ݻ^H��o]�~TM��З<�<O���ʼ/|d8�k��ı==��	=r-1�M�<�����O��z��=[R��]��y=&=_�s<�IA=��_=y�Q<R�:��<���\0#�3�S��yV=m�<r�N���)���s+��,л������D�<�"=��*=\P�+;3���<����D�%=��<*lN;��#=�N�< ]=�&�����A�<i�_=�y�:�Z̼�&���@���Q=1QT=>�&��H)�T�Ҽ�<8\O�o[��lB��>%���T=��������U��eɼ��H=C�<yK���R=�PM=(��<b<V���T��8�k�T6$�t?��jؼ�;�iѼ�z�<�����L��>��,e=�CQ��al=g�B�u[��km.��j`���4<��*�9���{}s;�`�(�}=u=.��8�=V�2���:��O��+S�[���	N�o-м�) ���;��x�;-�1���<}v�oWI=�`;=o#����{��"=b�̻J�<L�� ��0%�b9ܼ��5�%��<�E�<6$\=Gpo���<=Z`���$�>=�O=,�{���2��q%�GD9=���
H�<DF;�j&��9���&���"<;=�'<=
B=���<U�h��?��q=�_�; F)�(5=�j�<���ko�<�	����
�`�<_�<O�λ�2v�!$�HM��M���=k�%���~=�O�<W+���:=����>S<eK�<�p�»\=�U���j�:<M<��5��l��뿼�R����Լ��4;F��::7�@�;��f;)A���84<Jb�[�:*����z=���='ܫ<��T��2�N�J=�`Ӽ�jf�N�'='�&��L�<�dy=Pc<P��l๼����=5ف;%���("=��U=O�l=��T�
>=�������6���H=,�<����π�1"�(�$�����?1=	��<�]�?�9�&0��n/=��ػ>k=��B;��:����<'�D��R9�x�g<4͊<��k�k�B=|8!�!�&��>�;&�[�4�Ȼ<�W̼B�<�4k��[<����u�I<���<�3=I�$�8m輳l9<s�ݻ�ͼ@}��iU4�q��:=_Z='�=9��<j �F.�=�wi=��Pp�%�<d=[�Q=�!��+��*��1=g=L�{�,:��;�v��I�<t�<K�x=~�'��D�CNϼӆ<�~�<s2J=�XF=��J=�!�Js���*��!Z�;pC|<w�<�v4=�мxe����<��h��_=EM༿I��N�=�5� ;'k;�4_�F�'�����'�=�=>;�{@=���*,-=]䀼�H��I=�&(�^LZ�40���.���=�O9�ҩ ���v���8��W]��.�A����$=Ԙ<5���IU=��߻�����{�ANe���<�Њ;��C=��<<+�ݼ��o��(���{�=��<h�%�ۙ<%�&=EѼ���<�F=P:=����7�7�+6:��5=�ͼ<l;�O�!A	�ws���m<����s�S=T�P�Z�c�i=Nbw=oTw<��Y:)?<@J����L.ƼP�=<#U=o��`�`��0��W�x��E�<ޫb�,ӱ;R[X<�U�����u��"B<��eq�;Pd��%~=^D:��y��-
c��K�<"�W��04=��=5����8�����B	��B�<]+6�'��<%�3=� <���'�AƉ��Uϼ�p׼VN�<jΖ<�R=����ࣽ�p/=7G��4���?��R=���;��=�a��ӑG�I�&==F;��~;�"<X�f��ɮ<8F��u!<xݣ��<�>=IH�<ΣR�`�<����=��!�n�I�|��:�����=�Q�<�Z�;�@�<�"+��>S<��T����<4�;}�<Q���yNa��E�<��L=Y=GP;�0A=�h���<�.=)�B�s��<�e=���<V����2�:�u�<١M�Z�/�Y��<��=�yp=U���GJ��v,>�>�L��ռP
8�(;�6��p
�<�<a�R�u8{��80���=����<��>=� ںP0q=f��=��<���<eG;�P<m���%;���;�i<z!��op=B��:��U=��.=/�z�+�=Q=���++�c��=D��.�����<�_�;��7�W�*��<:˂�֋���t����M��Ў����G�D�q�@<:hD���Ի2�W�	��K�<��i=F���������<:\���^=��#=��E=k֎;��<�}���H.=*��<����;Q�{��<M���P=�󍼋=��
�e�w=�B=n��<�'=�V_<�D2=w;�N'=����N�U	���t�v�(��̭;G�A���<�\= �=�~�����̛<��;�D=� 3�NhN<U���B'�� 4=�qY�3�
��L�<�FV�����n�;-pT�m����Ѷ�����^e;�;�<��5���C=�Ṽ�rR���<�E޼��m�_H�,�p�g =��	�.�!��&�X�ۼ�8�`�7���8<&wA�w!S�#M
�Q˹<��#=���_�K����;������r�}�V��C��.�1�g��<��<F��<fv�.Q;=-�-�Vp�:q�X�ά�<�i=�8�<��L<wAż|8=�ʺҮ��5�¼�C�_�?���5\=����o6��E5��ϲ��PG=��<�*��h���=m���RL����<;��a�(=�|�<�S<x!�!��;�����<�B	�H5=�7; =� ��t���zY�M�������
�ּ�����G=�wں"�@���J�#�G=^I�5T=J��<�t.�|��<��@�<�F�E��<��<�큽��3�ռf�e=J(�!��<�[=7RQ<�5t:��/��t-��<=��P�=�ً=�7��z��L��<.��h�=�G(=���<&qD�y�ټO�k<�G?��;V��f���'=v��B�=r�%=A�!�;.��U����<�
��� ��ʣ�p�&��&�����<_-�Js�[`#�nYb=�y�;�hT=��)=-���"&��P��ES=�������<�Dռ;���<���<�d!=�Z�������=
�G=ۗ=��a<��*=v�;�e-J=�zC�9:@=�q��j��y;ǉl=%2׻���_=��<��I<��ZHG=�=m􋼇�D<k;q8�����;S�b����;�0�~7�<a�ּב� ڞ<����I����<;b<ٻ'��G�<��D=��a<Ox=���;`7��Z�<���<<�&��)M���<L�Q��׻�� �+���z�<fva�j J����O���9���#=�=�@�kĂ=�U%�|�J����<��<q4P=�L:76=�.��;�k���!<Є5=��9=�a��)=uĂ�GN"��tJ=n�8��z��K0=��<w�<��W=n����m<`ސ�r<��q~�<��F�h0=+�o��l���]=�^�<?E�<Za�<	�c�c,<��G=��0=L-!=��2�5��M:�UI��v�����ĻּUH!=�u��피30/<������9=�*�:�_��� <�48=nP�=`�=�c�$�{��EG=�z_�J]r�)��擎�G��<�c<��O�c�ry˼���<�Y=.����XQ=I꼨��RM=(�ɼ���:C1=*���<(=�h=ܼ==A=_Y�9�u�V��<As3�	9I�u��)u�?V=
���gW@�f<����IS��TM=х� 1R���M��-���v�}ν;j�<ɟ<�]�r| ���T�.>=�ɼ�1k�p��3�_��-z=C��=�'==/n0=֏��Vΐ<<�����<<�b=�ď<D�
=�h�=ߝf���L=�$n=tS+=��5=��]=�<��5=���<�35��0l<b̼�BS<�T9��G� J9���,=
=<�4�1�<�P'=�$B<7#.��-��J����q�<=*<���G_ �e�<���U�o�<����=0	�f�<;�@<���=�����>���	��IL=�5g<�h��u�<&���I�'<��k���=��#=(�#I��1]����<��/=�I1= T�~ki��)�?l��� ���<�R��E��]u<�1���/=�����Fa= �E<2Z<w���h����C%�������b�\� c�</��<� ^�����Ƞ=+�������<�3��<�<��;=��?=F?�M�?=K`=w�@��=��2�&,�=iL�<d�y<]�(=z<=ŏ/;Nz�<e�O�?��<�r?��"^���_=%�:��p��Y�?�<o>Y=l<���t���=o=K*u����:�h�<����/��<���<�"S=�m��\�	�=�݆<S7=�R=.9�;h�=]E-���;=6�}<��S��>=t@�=�5<8a�����<)rs=�|Q��M�� T=���<� ��2;8}T�P�������S�U�+���<���<vYZ=�.~=��7<�8=���<1�����&���D����<��<<����R<y�=�.鼗gX�!��7=���>=�=�:#[���G]=��Cu<$�9=K
Z���<�=?*�[�l=}����Q�����弟��K|;�l���a�:�,�N�y<:i��Q}=r7ӻ͊=�D"=hG=ja�<:�0���N�rv<bn�'�������=s���mؼ�=�M�=tg>�؃�:�ڼ�`�/�~=���<L�&狼���ߛ�&�W=����o�X���PS�
�ؼP�=~��<!��Z�R=�o3<F.�L�a��S�=$-0���ռ�$]���ڼ��i=l=H4Z=G�w�h�h=�h�< ��;H|o�:.G;?�t���r<f�<�"�<=�<�a=�b'=��
<�n2�L*J=nT=ψ=�\1=?&7;6�Y|��><�P:��w��d���I��|�b��[�]&���*���,=/
=MN�<�o�:�l�<�y7�b�?J�<A8]����`�<eO�<6,���:=��<�)n��?��=��\<�$;��q����<"6��}P+=u�<=��.=�	f=�}���: N	<�O���
��[=�G��m�=U%f='c�()���I�+|��}F�<�zN���h��#<�i3=Ҡ���E�f��<&������X�=�N��-=�#�ِB���]��C�`�ҟ:1���16��յ�FP���<�C�=�)�F�<V�@=W��r�L=�~��q������ �%�c<U=�]����ټ�C��=����65��1�<Ӑ�`� =)%=Rv�n
�<5;<��n=�C�~��ֽ'�Ĭ<���<�K=��=<�U=�
@��K�==�A���h=�1�;э=�h�nOt����;�0y�f|�<�T�(�-<���<���<������Ҽ�Y���o�|q������=`�����m+���J5=�<B�=�|�<��=IKV=-�a=j�O=%��<��˼�ڍ;��\����<.Q�<�j$H=g�续�=Й<hm):f����ȻP�ݣ��Ǡ����f��B���T
�-/=b7n��٫�nh�>�<g,=�N���t�G�R�F�<�4�<�;�������=���O�����;�s[�X��<��#<?�M<zpK;��c;�OR���K=�B����:k-�������=NA�;�!+=�>\<��;�0������:od��7����Z=@��<�Ҡ<L&�=t�S�/\���n�<o9_=��Q���<�b�<N_;�3Q=��`=���;=ZZ=z��<K�����������n7¼.�=Mfȼ �E���$<q�Z�l�;h5,�{n=+l���W<��<�<=�H�<U�+�n�#=�۩���;�5�����zq�<x�:=Z�k=NV=�v�<[�P�<5��3�7=�
V��T<��M��|̼ol�<�7*�����,,=�1=
0���z�!x ���Y=��x��Lƻ��ül5�<gy��I,)=E�S��q���<�<�#&<}rc�\ʻ����� <�=��0=���:��@=���<?��ilG����<\�:�-��7=��6=��8=��g=�1���;z"�;"8�����;���p�y<1#8=6��;�Z�<~;��h�<!�
=nAc=�>F=ǳ�<�CD��񧼏􁼲+����LO���ͼlt<=���<8:1=C�=�%W=��I���<�b=��<p��<4x���9�⡼���9e�<f>K�͇�r����\[=��J=��';�^i�n���c).=0gr=��<�#l��*HV=i���8���;0a�<��=�낽����0��=I0=�6;=�V�>:V<��D=�x�<��E<^=��(=� ;���<r�<����(<���<p���h=��<����7���`�*<l=�f�� 0=B��;-<�`�j�1�@?��M?y�ӳ'=<�y�s��;�G��>=Օ�;{9+�9�V�	�$�:=����-��˼�ZA=8�T=.�3=t�&=3m-=�rG����N`�����Q��cj��h-=�-���<��=�c�<�`�<�t��"�T��Y<��<��:�<�G;R�<���`=��5<�c��d,�<�	!=;:]ڼ���u�$=A��::�C�
��<�y�e|W�\��<�ۦ�#�(�3;���<sZR�$.������^<�Ѹ�jLC�4"�<�>R=��=���<��'=�^�������<��<P4;M�ǼՅ�ǋ{�LVȼ[�=kr=�k��y��� �:���=��mt��lD=�j=��F=��>7s�2ъ�����#�+�W�1�A������Cn[=F.����*T�r��<���;X�<:��`=Z�<��F�j�� �^=,X=t���3��� ���g�Y�9<j���S�k����u����_�<oq�<~Yj=�"�<j9� ;T;�yX=�g���`<��-���<BT=�N0;0�
=M軼iw��؀��|�м{ı<Y⟼F�+<m�<kk5���O=��#�����k�<�<�7:i�&=w�<W�<3ļ�q�<���<H�C<E���V���κ3ߣ<m���P<	TB=S�=��=�r�<Z�<Nv�����D��Z�<�,�<��&=��=�����M<J�<�X�:��q<2	T=Z0=��R��8=�P⼭��u=�%�<#�M=E�}=�俻@5�<\yj=q�l;F(z=W�c<I\<��<��J=��=�=bGr�hI�<i�z�F�<{3>�� =1cռk1 =z�	��Z;�˲<1E�;{�<���^J����<	p�O��<&�*����<>�������<�����T�<W.f=��U=����a�� �="L	=��;=�A�<
�=cR*=�d�<�j-=A���<�#a<l�/�Z'8�o9T=���yW���t=X�G=#o�<����<���.?7�)v����=�Z�����G�<E�=d�A�����kГ��=���ƥ<�3\������%��*���¼�wC<�㸤���r����<sF�=���=(Uv<B�=���D�;I=�H��j�<l;�<t�M����`�<�' ���;���4<׫>=G`%=�
ϻe�=s��j����=KD�<�'<��b�[�:KE��<��;���;�mf���4�qx,���3;�4n=��㼧G���t�ؕ����[����3=�"=k���B�<��뼻0x��:=xWD=��.<�3=�e�'�������M=��M=Ľ��e%=*�,��o���l<[�l���=��*�'��S=1q�!���5
<C�=�f�����P����`=���UQL�Ђ�I׿�[��������k�򢺻	Ң<�c���O=�+Y���=M����[���p=�gp=�0�����$=4����w�5^=��{���=���
 s=D����ſ<d���
��d��<��=�z=fw���������J{<*�p=��0��6�:e�b�/=��F�W�A=X��<4�O=���<Ε�?s�G�<p-�X*̼(q=+�/��TH��"�߇3=)F�?G!����ﺼ�����;x`��A���ň��<m�x5=Å�<�#�<�C@�`�<���h^�	�<�����o<!���,�o)>��[=���<_J=��6���E=��#<8�����<)٢<P�����p`<�_<��.=$"�-\'�"�P=�v?<�Va��b#��U��[M=�v�<,���B=�|�;�<>�x��Lw��=��6<^f%;lp���" <6&W��0����=�X-�X�F��k����L�R��8=���;h���W
=��I�Y�2=qKH=�P;��3=0��*�
=�U�����<�1n=��U���<x5������6����R=~<S#O����}�����r=��@�Wt�<V13=��4eq;� H=�߼��=�콼1���ܺ$u"=}+��$B�<x3G���ܻA��9=�҈99����9<(D�<�+�d��=�Cj:�^$=*��<�p}=j,p<��2<�tw�p�-=�q+�{R6�2G���<�q��xL�=��<��e<�dͻ/ٻ��=\��<��;�vӼnf�����!�;H?�<�n���;f19�?X���<��μۍ_=�-=~=�<�D����C]�x?����I��1�<0���<J�<)|$�|P�<��-<
@)�2q>�UZ��2l=uA=�Q�/Ts�����8<�F:�9�=�F =��<򁰼CL������Vq(=1�,:/��:Jem=!5I��i�ԙ��W��;=��<��=�n������/@��U=�!�R
�<�>�6�3�d�7����<N�8�i��<7W_=���;�����A=<ei=0��<ψ�9u>_�)�<�m<��<�c���1�NA��;@=��<e�r=��g�=��=����M=x�:n�:�st<�h�<G!���<=�(.��8�<7B=��K��N��A��;��<liN��>�eAw�a/�"�`=,�<d<��:��fb�N�ټ*V���u�Y%6<c2+�Bb3� �=��ҼF�A=���}~=_�ƺ�r7��\=�*����<"�O=�=���7R=��<=2n<�y>�;`L��{I=�Ք;�L�]�8����<ȣ��+v;;J�<.ȼ�5�[[G;/,=�k.�gr7��ɼ��8=|a�<˳�;.���b��	Y=R����s�]��M$=�;���>2=��$$���a�;`X8��5��1�<Z[=:���ۅ�R�@�᯼�-�D=��{=�ꓽ�\=%N���"<y�{�En?=[F=��<{Κ;��</9�<TJ��@�<��ػ�=�dKмQ�*=<c =�1/�'u༻.C� %=ށA=��S��<}}��|��<p�=�->=������=$=��<��<<h=����,������/=��E��=��2��ݣ����<�a"=�E6����T01=�����C��_Ϲ]����<��7�dE��g7⼛T����v��D�g�n��"=��<Г=�A�#]�;�z ����<��l=<ⶼ0g;�X<�Ǽ��/=�m�<;鯼mm�NV3==Ӛ:�	4�#2�����=g9=����]����<z�<������<9%�Q��<#�=X9μJ������%9��*ܻJa�=|]=(�<�U=��[;�׀=�-=��v<��==>��<:�+��<��c<=w����t��7{��)�;��E=� =���<��ּ����H"�H`3=���S<�
;=;��<.yS=z^@<\1:=�`L<I�.=�c�j��ZN(��v"�x
=������<�I�<�4�;v��:Sݪ;ʾL=_qs<!�#�4㑽��-�t�Q=�n�;G.7=�3=
�	<�<l�<�R=Z�e<���0�[��;6O�:��t���r�r�μA���W(=��#;^��(��<�ȼk�U<�)D�"o�L�<���ɼR�q<=�y�rD=���=-ݏ;$�a�I
����P;�%-=ֲE;��U=�B���m弳j�=�v��ꈃ<��;F��Fl=S�;���<��(<Xϼ��
�<r����(=���:��3�M��Z)��~:��n<�z�<��ۻ?)�;�A�<��r<��:�H=�&мg;!<��T<ޤ?�#�3��D�<P��;�.�:`�G���;��V�<�oM��1<��O�<��<s
�<�e�(*=�<B�:������`�<_=�CV<�)=�Gh=�U<y�����&=��;`����ܐ���<�u�<��ּ2s=�=L�]���G4��C=�GZ�o�'�
)�<�'0=��'�oL&=�	�<Z�=�z3�WVp<�XȻ{)=Ѯ����<�(�V�4= I�=�A�(�\����<0��'([�	$Y������ş��=�=��#=���;����Qc�<�ᆽ�ړ���������[=����t3���M��D=�uH=�6�Tm	=KG��.�="Q=���<��%���<���<�;�;k�<�s�<m��<��� �{?����F=���<1�,�P< �<j�6=�h�;�3}�g��c�<=�ʻ��;Q�=۳ûUki=��7<���k�"��F���V���k<xh#=�m���낽8 �9�T=�K�Y�=?W;4�m<y�u�۸��ʯw<t��J}=�o�F��<�<��0:�-=:�<AFм�Ce�F)���H��}�sG=�<D�g�m־�79<��I��g�<KA=�����;���<�g=����a:��SZ9�!B<����:<=RQ�=���`m�q�=���;��%=}=:�<�Y��<��k��
)��WH�lsV��;��n�;�G<�׶�𮃼➀=921=]D�<��=1v=�q�Zue�ݴ�<�2G<�,= �2=��	<�oZ��U�w=Y �:ؒ�<~�
��*V=����N==z<�}k�+"�IHJ��λ<)n=-=d�`��<�?�;i��<A�Z=\b�N	)��O�:l���%,=�h׼&y��+���"X��f=�;c�V�� ���<��<�F2��.���<�<�<E�<¯.</3�<�ٝ�߮=�
`��:D=��/=X�C��+-=X�<�9���+=5h���<�̟���ܻ7�D�����-��w=ds���<�>/8�a�<)g ���=��T�l�L=��?���g�� �&Y�MT�<���<Z>��j><�=�Ff�p*;��F����<H'��dk=3.L=�K=��=O��Ο=K�2<��W=y��::�=��vwY��#�+8���\ ��?�<&�⼨@0=� ��dx�<r��<b�w�Ra����<���Hzn�;}�=��ļ����a=���8$,��{�=p�<_[<&�A�4>���ür�޼��[<�����A=OH�D������<ٿ���k<6~?�'C ���<y(�;L����y��=Ђ���o=�m����.<�j(=#f���<��<�VF=�[f=��L=N|;�1#=w
8=�𼖿�<r� ;|���	=��=�=�Q�(�¼&]=�zQ�y�'�T_�:7tl��<�"��ԑ�;���</��f:	�(=!<�2C�Tu|�v}��wz<%�;T=�_�;�?V�(+��g���ؼ�\M�Y&�&��O��9EC=$��φ��+�;�= "g�߰�=�2Q=`7b<�d����!��<e�ݼG���@<�W����1�/=Sq=�����KQ�;۱��~�8���=�I��b�>��
<�X���^ܼwb=�'���<�����H=� ��o�h<:	�<^�<�|�;�
��fN�T�<���o����;��j=X�k<��g<�[=t�(<T<���Y=�Nq�J4�[���G/��+1�W��<�,��+�:��_�t��@�T=�S���r;�C���݇<�w�l������<�Q�<'I>�c��p�<ì,���Ӽ��$)V��kx�F�	<W/�<�!��F=�����������lS�<�iy=�z�;W/��N�ĐQ���?=}�A=t�'��s�<�FK=�N�<?/=ȃ��"f:;+ ;%|x�� =���AF ����|�P=��<������@L���V���=c�[�����AA��U� |�<"=�L<�ĺ<Ll?=��߼���κS=�H#�g��H�Ҽ͕����=���<�*��X&��U�<թ�>�S��<�ɻ�'�<o��V��<��F<&��;x	�`�ü#9�O�ȼŝ�<���se-�����Ѳ<�����G��w��/@�%�����*=k��;��[9<M�<��<�&��lt��$k��+=����<v�ί�<�b5��o���;���G�/�<Png<��B���5<��<��2�.�;s0º�J�<�.S���������<���<��P<l�<���<��<,�/�����E�ż�d�j�%<^3-���>=��Nk ���f;Q��<à=.&�Q7�{�+=�a�:�z"�O��}�H=�2�<��g�@�Lf0=IJ�<�<�6�k�c��_ѼnUV< �*=B}�E�r=�9=���<F�J=�Q���_ټ�p=M�Լm�1=XD���mA<[�Q=���<Ltc=��̞.���*�!b�<�����#�( �!�i���3<\����<畽<�]�<?�0���[�ߴ�Sea���;ka2="ޏ��Y� �3���ip><\3=&�<`�H���=x2=Sh;=;<�=�U��vu�;����T�=�H�<��< /�H�<N�t=�Q�;�5;?�����;=��R=*�,=\h�.�x���1��Ƿ; j��E��<��Ƽ�S�;�qv���J��'����(}��e�i��;=��r;h=��L<�N=ѕ<=ځt��T�?3�8hD=u�w�>�
���`�ü��Ѽ�<�.L=�-��� �<wH�;&_j=ɸ<�9�W9>���/��`�<�6=�=���<[ht��Q <Z҃�3A�<AX`=�=�}�<��<]>ټ;�9=A_k��w���==-�=�t?=���<;ټNv����%<蒅��!_�_�	=c�=��A�K.�<Fd���o=�eԼK�=M���}�=2e<I(f�!���`�B�_�b=�J��d=��u���F=��<VU:;��;�J?����G�7��'�N�<.q��Y�<�4K<�j���k=�U<���Sg��U�<^�<�r!���Ҽ=������[b=F>��L����9>0�Y�ü�;,��0O��ȩ���J=��z���'�� k=�AJ���q=�=�ϡ}<��;U��<Q�	=�|�g.3� �4;�ȕ<�P�;"u=�<��O�<�70��);�,X��z8<�x{�4����=8r���ػ�ҡ���<bI�<�J�sp.��e&<�1;�K�<>��<T�<� <.<Q�ڼ_7e��Τ��A	��A!;T��<�o):KT�<C�(=ט<��<
璼�6��l����=���T=�T������\�<��1<ܱi�	U�<�fl=ٹ��IJ��켻,Y��ˋ�7p����:�7�<�RC��N�9��q����!��HQ2�F����s��1D=� <b�U��<���E��<���<ڙ��o���g����ڸ<�.8=�X[��o��u꼁>���%=�m=�7�X0�;��ݼ��=�Ԩ<������ڼY2]=�
(=v�I=(�;r���_�[�;A&d=�����1E<��<��X�����lx� %=�KC�x�Z=��0�k>�A!��~���/D��:1=�i�)S=bD����X�%�m;k�.��E3=M��<�:3=��=�Ec�����E=�f;a	Q=N�v��O�y�=��<�������<�����s�Q(O�װ$=�|B��^�v�¼��g=3���!O�^�5;�v<�?��|=�; 4ȹԇ�&v�<$L�<���;���<���f)Y��f=�#���
��ǽY=��; �:���B��z��=/g;U/<����/�sV��_�;���5�;C�<����Z&G=��.��ip;��+�ŉ�;W.�t�6�L+=���<pT���1P=i��u1=�)=�X���<��>=�6ǻ�DL�3V!��Փ=�7��&�}=��;��K=#�X<��r�bu~;@�b=`�<'��<\$g�]2Z�oE�<�L���y���즻����2 ���>��[��D>==�q=l��<�I����<�׼Q7�5��9�<�lu��#�<��;EPr�~�*�s	$=�e9�[̼�<�e�<Tg'=��G��';����#A�<;/=�* =j�4��2üX�;=��r����%��,�;$&Y=��0��1�<�P=ܵY����<�d���=�f�=l+== .�<���.ϼ8�J=K���p�}C�F[ =�sL�yʦ<��L=�ۚ<�#��Ô�;$��<#C�<p��<�ʼH�H�x���F�͘�<C�	�1�=B<m�q����� ��C�9��=Rg�j��<m��I��z�-��:i��!=a
��-ٻ���;Q������;K��<�o`���i=���<�Ց�7�a�,�߼`Q=��8������< �==����G��l����<��!�<fY껝;v;BEb<)�y��)t:����zM�=�PP���j=�4�;��O=P�M�˻�i�<�Q�<�s�<�:\;6�X=h�A�v��;���<�X��;ۻ`%Ѽ��#�vk<r��)P=:k��R�<�Qg=L� =��Ｌ�N=������x�e*k�R�v<9�g�<�;D��ټSV�<_Ab=0��k ���>�=5	ɼފi;�Щ<���<�샺`}n=�_E;z�=|H����)��*<���<�v����24��p=�R�E)�<�}��j=;�=%=,����ѼB4�<꜉���9=��#=�晻�=��;�ӻR�{��<!�M�=qva<πb��V�<j��^_-�Q�T<��C�F?�I�仿E����Df=�kE=�~�}�<��t!=�e�����b}=���:�8��=�<�_��H<�.5=�Ni=e�=j�T�R���^_=�G��c��3O<�*]�(�l<����QC&<>**<���;��=T2=������=$}O=�R~����<�»�&=�/��Ew���c�۴���dO��3���:�-ݺY�:����=�^�3�+�������U6=��<�Z==%�<�yN=pЌ�g�=���� 5�;^�<"�=���,��+=ׅ�<�*�<sG_<�e���)���<1;�<L�N=fR�<��
�4sF=Q.�;U=}0�<"[*�D]<Ё�do#=�*�C��Vp�=�7s�0�m=��~<5�<*=	=B�<�2A��uX�A�C=�o�<S�*��%=U�>�����n;�Y!==Y���<��F��
<\[`�Yf�<�:7<M�ռ��0=l<=$���$��=�_�;��`���$=^ <��2=�f/;�QR=�uW=�{�<o@̼<R�<v"�T-==�W׼�a.<� <?j�;s6�<8=��-���0<��)=};��Tg��܉;�@=>aL�G/=��I�@�K�,5�:�����4=���J�b=qX=~L=s�@�ϮP�:ٶ��OD�#�z=�q;�1�μ���;U=2�<qv�<]\��(�Jp�D~ߺ,���,=�Mȼ���<�:��Y	=g-x�<#=pG]=��(=2�[=�`�<տ5��h�2?=�+�ɞ�<��*<�~�<�_��=�}�<�j_�lH�</0�����<�X�<��G��g��K7-:�!.���J=r泼ވP<$r�A�pʼE0<�"�;�"�<��;��Ϟ<����#�<�Q�;K�D=JÆ<�#�jCL<~)�< B=r��L�<��+��-=��;^'=���o���M��<BL���$?=T%=R	��'��E�<:�;<Ɯ]=��"��q/�{X;=C�<�;�4p��� q=�M=��1��o�^��<�ů�����ͺv�N=���7����_�_=��f��NԼr�R=�3Լ�C��rq'��.a=�XD��L���@�I��L�ӈ�<|�0<(؇=)/���4�<ܱ<x�%��O	���F�	��;&��<�6���`Ҽzg��,=����<�E�<r#�<h3�gN���=� �<C��;�52=v��H �<U��+:	<��r=�¼�-���E�$<�<GG����<�D��^-=C�e;���;}���9g�yIA��Z1��<i��<e�4�<�Z=�o��`S�AwT�BW=;�мfU�<��<&w���:�<6�<�.<ZA��=����~��k��N��d�z��B�<߄�;|UY����;�f��I�g�pe"�>	��,j��UF=�4��=	B=�߼�,��ag�<R����&U��')�g�*�L5=���<y��<M�(��\ ��s=��;�@�<wb�oC��} =��Y��3=�k=��<&̹�dS�<e��<-9���W���=��r=A�~<,=��;0k"���׻g>=~�=42��I= g=��"ü�P]=��G��Y�<�@4���i��=�*���=�r�<�K���;��ļ��e�nc<�vzR�#�N�xl���=��;t�P=i��<�(_�� J=Bu�5G�� �a��1�%��<��c�3�3�;�l=�u�<k���<�<�j1=Er�<~�Q��C�ǰ�=	Hؼ�>�<$#J=�;�$�=.�<�TZ��ya� �a=M�� <��ӳi�ޅ��_s��V"���;=0o[��SG��*�<
`4=w�����e=�=!|`=V��<��<ڵ�<�ۑ< g<�%�<�5s��z����=�x���<�u�"=�U�:�tP=�<t�<l�4=Fn��f6Z�wM=�a�tH8�A=�68=_�ּ�Q.�e��;��P�A{�<��0=�8��v�$q
=>=_<c��\�=�=�X-��K��A;���TҼ���t�P�F��<��y=����8��s5��5=�d������@�V���ػ
�'<���<E.���#�B�Y=ZO���J���^=�X�<���:�<�?=��0=y��=��!=�C����c�D��p����5=��>���
=�<`�J�
��<��y<�o��<&=c4�<2�%=���4r�<��9;��J=���<��"�l����k�<K{p=��,���H=��3=��м!Φ< � =�$/=�m@� �R���=w:�<$?:�Y�\<U��<��F����Y��z�=��a<���<�E#�O'Ի�9�;�U��e=��=K�ڼ�}f<��)�>G�ڼ/�A���e<����h=���Ǳ�<z��8^�ڋ<i盼 c6<�r����0<��F�3�=.u0=JV=�=��	=�B5=�3�g�E�?�����>=��:�)���`��ŷ<���;�J<�$���;ݍ�;4�8�E�E�ҏڼ�R7<oҼ�L ��׏\��L <�;�<�Z�<nx_=N������ؠ�;L����$=�=V �;�lm=L�1=c����lg=���<�xd�Y]�<"���1�\�0�rsǻV>U�!w�<�y=�'������GY��?��t�;���<���<���̬�<.Wy��=B�������;
(�<`$9@W=�1�<L�b��|=��O<��=�� =�?7��U=6��<n��;��zӊ�~�k��-=�Qм�E4�?�<A�O��k����;��;�|;C��7 =�8=<�٨�*��<�4�<�0N����Og(�=���b�⻞i~�s�3�;le�H��}!=����#H(�'����p�#��L\���O��h�=	�:�
S�+����x^��
�<8=��$��s��z�ι�������Tl��Z;���E����J}��v�<)a�1=�ȉ<�Vw=��F��/�;��<�s��T)��	=��=q��=z�D��z7�9�=W�<��a-=�fG=]���2?�<u�<n�ͼ:��q�<�{`�;��<y*� ������=�*��C
=	n=$�`����<�dN=�ʹ��-�ӶH=^��;��&=2F(<Ѵ>��0��8�<䗁��K=�8������r伧�L=R7����<�1�;�2�<8�,=���Ҳ<[Qu�-�p=s���q�u�.�Dqh=�?����XQ��ܼ�U ��=oу��=�f�<+�=W2��/�=9u)�����)�<�e�8�;)=ᩎ���{�I�E�׻����P=��<�Z���=�G��!ޢ<\e��4P�<ӌ=f�<��]���<s#��S�<0v7=ȸ���r��×�M*�����<�����c�
�[�Γ;nL;�I�0�w�w�b�c�[@�ᐚ�Kx�<����Ā���Ǽa�<���=
�=}5�<1�"=e���}��;���:��<�<�C��r�<-|��A;c�ٝ=_]"�'6���S�����R�{�*:=� �܍=��%=q�z.<�~|�5�=�P�<�����=)�n{�:N�g���;�"k���W�}J�|=�u8=�mA=�(ӻ <�઼�l=�,=/�u�`�<��ٺ�ƅ�X�����]�I���)�
=b���@
5=��[���=���n��\B�<�����=�(����=Q;ѻ�T��9��B7=<�;=tV�)'�<�y��@��{>�;�� =<��˂=�[����;�x�=��<��	�}](�����gj<�K~<�"�GtQ=%K!��r=����`t<�=���:=
����;b�L���u;Z4<���<Yk��nWX=�I��͠f��m�<�02<ưk�ni��&�_=A�����<����Ǵ=��<S	�<*1f�{�ڼ�E8�`&=��b<�V�<IԌ<�K2��=�f��=3�;�<�#���#U<��w<z�#=u�,={�'-"��»ᕽ|<��=`0�<V�i<|���Q���R==?�=|�7��|�<��=�����7<��c��g=G�;��q��=��<�bԼ�1:=ٟ
��]�:�6�;�����7�~�G� =�a�h�V=�;<�v=�J����<I:�;(r�<V=f���\\��ƈ=�u�;(F�=�C�hk_=b�:~l�;2�s��<r�3=���<�SD�NIu<�/W=��� =P6�=7,�9����Z=K��;�7�:��O	9�+򻡭�<
YǼHw;��x<Gż#�o=U�<6�'=#�E���A=]���7���aJ=�<W�3=P���fS�$����`��G3��3�=�3��WS=��'=�2[��b�
Z���Թ�� ��q<���I���*��<�q�t�r�C�޼�d�<�G�"
=�M��\S�@%=P�Q���λ�=���b�
��<�EQ8=�
��.�<�q=�7��P�<z]��(��9U=���y?���#��B�<��]�G	=����������q;�9�?��'�����;n�s<M<�x=�N7��y�;��W�	"9�'9$=�!���i�<�1�<z�C<������#=2�=�ݼ���:Jv;N1F=6�M=�J���9�E��A;�<��%=T �<��h=��=�}5�n冻�1m<�Q�eB=��*��\=�~$��a>�=��d�U����]����u<���<M���^�<p�=o!���@��l��<��T=���;�Z�<2�F��XM<��g�0?^=���r<}40��0��Nv���)=W�N�$�<�g=1z�4���R=�D:��$��#n�B'=*J�<�S�q��<!�O=��a<<m��E�Ļ+D=�K����9�<���K<�_�<�c��;�0Z��Γ��8����	<|�%=A���C8=l�.��h(=9˟<W�g��tG:T�H=G�=OC�<���<�h����;�32��m <�ۖ<�ϐ��Oົ���I��=�|<� <�=�G<�L�vv�zH�;���<9w'�(��<Y��txw�>7�<��!9���<�,<+�S����F�<���#=�Ѓ=�TL�bHм�]/=��W<e��<x�%�!�P7����[=ʔN<?�x��F�<�0F�|�<$��s�<N\�<��ʼ	�V:mf�,-^����6��K�N=#�����:J?��z�=��_=���=�
���A�Q�V<X}<�����U��x������<��I=M��hE$�8���T�:��-=V4<�=]r.���=)o:=r�9=F;ʼ�
���u=]�=���a��	<[Ѽ�=:W�<֓�V�;U5��kV�|�
=p�M���&��?�<CQ<���<�����u='���Q�7<ֻ�=|1�������<z���]����u"<{=�A�X�J �W��D�n=�`:<���;�a�<!s�h�<!�w���5=�=����=��;�%�<�¦� X<�A��$%G=w��<�4��NHX�;�M=1*�<O#U=��=���f�=��$='�=N����i�<��D��<�b5=.�I�q���`f=�ex��B=�QJ�A+�<m�=��=x}���T=,[r�3R/�M���5!�<��=&/<���=���B�?����s�9����<�U������T�O=0O��Ƈ��(y~=N�=��<��x�6��%=#r�rf��=6�5�� =G���dI���=r�q=��A<��&=4�r��^Q��Ӵ���w=*v��q�)���W��<+o3=��5=m�<@�q�j�����;�o����<�sʼe�:�M������=`Ƽ�)T���|;߇���=��<�d=��q������0ȼ�����e=1��ݗ<�)߼s&B�"&=`˙<0Ţ�1��45��n���н(<"�׼��-=�A<ngU=a��;Z]�<�*�=w�[=��=}p��x{��B=���;�u:=�d =�=�Q��9���
�(��o��+�|�B�1I��3��<������<��̼5��QD&<�rM�O4!=��3=A
�<l��<n3=&��<��/=LI�?S<��"�L�U�>�@���7�i�7�g7<��=��js���9�=��_t,��y�\�����2��-���%�i�T63��u<�%�@L*�ޒ_=L�2=�h=t�=V��o �E����;.H�=(����%=a�<��;���O�D�א=��K0��(�<1�)=��V�k5=�5��ѣ���?�;�K�(�%��B������8�<=t�j�9o�;���<���Z�ن�=��<Y>�<��0<˕������l�&�I��:_�+=�/W����8=�F����<��w<DA�������<d����1�i���"��<s9<���� <U��<[7=�K���
q������'=	��?^2������W;�f<���<���<́=If�@=��F<��d=-=��=��R;&�ջ���<:J�џ����=ψмՌ�<��x�	K��#�<�=Ǖ���)=q�������=��L��U���>=�U�Թ���NT<�����<�ݼB���?�����N=~ie��<x�޻��<p�=����P�;��3� �'<��<�\e�G��<����< ��<��4�"Յ�� "=�(�nE<I(s<|;�;�3<��<�����`J�R�<���<���;_n4=�e�<��z���B�l�9��y;0O��Q|���4�Z`&=��6���!a/<���xg#=4m-=L�K��"��L��<��"��=��l�|�f��!�Hj�;S�=a^=a�ѻU�k��nƼ#O�;6U=NOb�F�<QQ�o�,��Y����<��W�`�Y����k�;��<n��%M��S=E�a=o���<tG=����B�
��
:=̀I=d=���<�
=�<m:�Z���FX��U�e>�6MW= 0=kZ�Y�<[;P<�%v�|K6��Z/�Շ4=!���|��0����<d�=~��E.����:�ex|=IƼ+b[<���߁=��<��<l{y�����G=���<�6<C��<�f;=�췻z��J�K����<�`����9�y�<��7�B�<�<�9�b댻jA�<s	Q=�-k���g=Dif�𳨼,�<���zc������)���<ޥ&=흄<u�<:D�=��O��P8=�#\���$�dq�<�Ҽ\��;�s�A��<�=2 �<4�:m�����,��:)�<P$=��lȼ�fM�����N=�fe�3�G�?����@��c=ОS�W�oq�;��=�+��\g<;g�<���  &<4z�uq<�Z�����<��9��犻�9=�L�=��<.�ݻH�V=�)='R����O���3�@�n[-��~@�h~r=цG���<&!�q��<EY�<Ӄ�<��l=��T=�W�<[�?<�'����~=AV�Ov<��S=`ͱ��"���<!�I���=��<9�<��<c�퇄<��;�v�<��<i�ݼ�@j�;�� ��9��`=@�;��@=Tg�<����Y�Z<`�<}��;Z�,r�<�KR=Y`��$QI=�⼨f(�P�/=������;�v�:0�1��p�:1���Z><5A��G��Dټ�<X=�d,==c�<��.;��@�o��b=]n�<ؕV=�u��a.�<e��<�>C�,�P<�M�� ��ҳ�<dͻ�vx=p�g=|�S=�v�Cћ;�!k����<��G�&l.���7�+�=�#=�4=�_=�/�@@C��Y�<�@H=��2������<Y�_=��O}!=Ш=OO-��(�<(~C��B���y���K�'@=�0�<��i�����D<�J5=F-=9#B<�=�z���Z��nO�����<�'>=nX�<��R���μ��=��`=���<}Ć<�]��:�<��<��d��P���;=�|��.��j�F�I�$�Ԛ���EU=�b<x	x;A1b��t��h�9<�E���Ҽޒl��4l;����=�GǼfW��<rl��ryU<�c=O�D�#<}�� Y<�楫��G=���<��(��Q=�!<F!��)%�7o���$=)l�<�W�s(-��FM�#�T���]F=M�Ȼ?�a;ཀ<�Q�������Fμ��E���Z�Yjg=��;���<�:�<
ig:�C�m|=A�d={�<<�j��N���l��=�=�S#��f�F��<g����Ž�y�w<� ;Dc��kFּ,�4�ȴ ;y&d=3����ֻ'N�<���;fs�P��<a����A�!gU���p=yc={�<�b7<m�=��=��2�Y��<"65=f�/�D�F���5�܈=�<��
=�c<��=��U=�<��7=�����+=����H^=��>�x]�<FcO�P�"�w���a|�����<9}�1�a�=Uj��T�h<(l��c�̼P=zlȼ��������{&�T���!6�M|[=�$(=�<�<)H:���!���=�|:�� d���I=�(=z?=�<>�<��3��6�96=S!=�ne;�T�K�Ƽ�sü�oM=�+�]�<�`<��[=G�D����;�B��j��$j,;���<�8�\�<��G=gzO�x弖��j<iC9���<T�#<`}�慦�b�{<x딻!�`����:�n<�x*�<ӎ<qY=�S���~=�`�5;5�"<ּ�s=�S<��u�� 	���<�G����������=��A=L�O=�o;��m��6�L=ѣ���;����h���w�4ƃ=�,W<_`�v�X=�TW=&�<��I���B���)��
���?���6<[>����{���3���»��D�7-@� -U�ei�*R�<7V�/>=N�=B�a=I�f���=%����:=�}�<��I=#��<"p]=.����������=m=�I?<u����8��HO�Z��z4j=�)q<{�k�ܻ=3˷:����מ==�w�J6���4P'�� �O9=�Fr�x�W=$��<T�T=X==7�4�gk(����m}=�7�u˄;�ab� fJ��qg���޼�v;�v0�kP����<=�:b�޼��Y�6�R<zL��Y��<zzϼm���s97=}��<�Vϻ��5<�ګ�.+�<�KR<���5��������{�o�<?��Kw,���=g'�ZxF= �;�O���4?=C�4=��)=�Z<oE���4`�P$�<�g�<��7<�k<`4�<�я��Oż}/��\ay;"<$�Oiy<���s�`<źF�Z�^=,Z<0񩺙��;M�O��^��劻�e�<[�����E	���<���S]~<!}5�n]�7P���[A=&]⼁ܷ��w%��l	���Q�Ⱦ�<9Τ�F`< X�<�4;��<�RH�AŘ�����A=MyQ=� ��C�5�[+<��Z����;��n<��<�Dz;�p=C�<ת=�7�<���<�6=��<����<,h=P�'h?�����=��g%<u�f<0!���6���7=N㒺��z=�u�;Yi�<�<
=p`0���7=_'B=,���f�0=^�@=<�=��=�P9�Qq6=����?/<�@=�ټ[��#���
/v<��<M��mA=p��WD��[/���S�<�	=�F<]	�;{�U=w��u[U��'I�<�<�;Ҕ���<�}/�t_�=�/=��ջ������=�gj=�~-���U�"AS=Xg��91���W=�d��@g��u��GY:�y�<�Z=�g�T��W�<���4�U���v�5�C���=�=8�W�M�������O8F=7<������؈<��5�[;�|�y<H?�<�{ȼ(�;��>��C�<��w���&=��������<�50���<��=��z<G~ =%�"=<�J<p�Q=%x���K:=�����뼐,K��%�<T�6�خ���<3�.=i�A��:M�j�<��]����<%e,=���Aqּw�-���z�pRͼ�$�<to�<m&�񤼈��<mDX=�:�S�=��~�|�u�q8<�h=�6�]�� =oJ=�]���)��\�Q��f����=��L�l��<�#�<-*���ɼ���<�g�*=w*`<��=}�<�Bۼ�ie=Li�:J�;��M�D_A<?��<dO���9�¢w<t���"R�n�[< �x�ػ2<�$����<��V��t���� =P�)=������� �< �I���i�O�M=�/i<�����<��޼U�2�hwW=��><]�������8=R=��׼CF��V�<W�+�7*=f(���D�m�:��ͬ<���<�kK=#  ��ƹ�-�̼eҼ�z=6�d�+qm=�*$�Ȼ����-���7�l�*�B���K���ٿ�=��0���L��!=�D@��D�<��<���=��\��C+O�֜H����:c�IeS�h=>`��(D�uQۼ�	�;3��~ӂ;e���:z�<��L<}�_���B<�C�2��<��ڤ&<X���̎:=P߀�/�\=By�<�A��2����=T�鼷�<vʰ<;��<E�C=g-5�T3�k�g�E<p\���M< ���k<9�����=���;��<M�p��S�<
<��=��k;��P<Қ �Y�3=�v��*5!��F09�!R�h�G= �<}�>�(��T�c=�͋�=�=v���ve�<�}#�x��D�;){����v=��19��+=}�l����	9��g�_���l��[�`. =>�f=�&T��&��Ax=�żd�"<C��RL��E ��"�;�;�<#��;����m=���<)'��h�:=�C7=�G@���<@����	����O<���<�c�M�;M��:P��N=�������	��9";�q�<nHe�:6X=�K=]��'S=��	����ӼMa����żu{=_��}��<��5=H�T<�I��w]�Ո����g<�iO��%^��qż���p(���,�o�j=R7=4b��N���G=s��<���U��r��5\v= �A=o�h��]R��C��p�^=���T�,=�n���]=KgҼ0�(=��.=G�<����9�T=�M
==E;.z�</R)=w=>�h�$[��w����߻�o=����j<x F<Se&��)�K�3<��I��<x�ʼ�c������A`<ҡ=��1��;���-��9�+m��t�]�	�v�P=8���.�δ���<WWD=�p�Xp<aqu=�lŻ@��<8�+�H��<�
��=�<�II���� �W�O�=��<
��B� �8�<'�<�y����;���j��&O=��v<�=��6�����=�|�<�o=��e=�<�ԗ�>�H<+/=�o(=�Y=�8���7<��:�<����=�]
=�Gs�;�<��
=�𳻙����k��è<��<%���k�o_��SX�: <�.g��Z��3�=��<k��=��r=x=��E��<X��<��@=��缛G1�>&�<*�;���\=��5=ߚ��+����d���6���g�QTＣ =Af!�8#F<��X=�r�}<�w�<t_��!=ue�`s<=b�g<�� =BM��8H-=��9=5����$=b�[�~n�<�&X<�%=�[s=���<�y<�v=�	]��Mf=Hb�X�-���=6� ;&�<�<)�W='|�;8C7�$����;������X=R�X���r=�Tj���q;.0N�A�4��M���X�:t�&k?=k��%:�<��	=+��Oe��9�=��Y�Sq������μ�Ҽå� K�<rջ_�:t���,=�{<����=>=XG���V;���<E�^=s�!=�=W
�w���%�<dx=�.=��=��i;��)��� =�\����<�*�Y=h��<�s&���Y=&�`����2.�;T4Y�La=
����:�G=��<��Z���U��=�����b<��N=��=�6.��83�76_<�H��F=�:Z�f��<�`E�z��;�x9�e��z�k��<�ؼ��}=�l$=r�W�dE<g��; ��-�:�;��8=���z��<�ބ=��<�Ļ�1+{;�x'=�$�j#(=�5<�-�WS�9|���;��O=�
��{Ǽ��=@����¼u�*=Pjf=��@=�=�>D=S��<�4�%����X���<�lR�XE�**-�7@��G=�,�M =K��˨�=�J	=tbY�^¼�p��@9�<��>=�wh����~�<�;J?�:`M��.��ύ��X��@��BĆ<B�����(�Ǽ��X�˟=V�T�|��<�y7<����/�F���_���h��;�9��	��;�t;<��8:�92��$<�F�х%=� =dO
=ڝJ=�X=��G��k=xX�<�=[d0�eU=�n;��ƃ�|�<�p� !=�6�<����< &=t��<.��<����<]�A�����)=G��<Q�Z=^��<�ż����I=ϩ�;���<V3V=���<�]|;�=���<��+���8<j|=��O=��ļ�����<̎�<����R/=��L�:91=a�����<��=1Y=�:<������G=�U�<���ZA��_���gJ;T�[<�~<�He�^n<mZ,��#�<6���U:�9c��W=�O�<�@!=V�M�?g�<��:�X*�@�м���<H� G���ܼ��l=��=�<,=�V����ܼ<�����I�����X�o=+��<dO��(=�;+<Š ��⋻�I�<�nѼ&,=7^<���~=��,<dӼ��+��+]�<��<R��<��<��Ƽe-^�ǻT=E0�<U����j^=��Ż�zx<�y��ު����/���ؼjJ�<��<��<9���G=F���.�����<�mV;�e<]��<y�=�b<ydX<�����"=4`�<��<�Nt�E�=p�8��q��-��:e���;����<6�׼�=\��<d�	=�a��d�»�%=�t���7���<��\���;=M�=P�<�����P�ȁ_=������u6=��R����<�n�< < ��
��@;,��J=+�&=��F��i,��I�<��;�$=�5߼�=%=\�W��(���O�&d^<��P�t�Ǽ*J�����خ�8���<�;s!�s�[=�����	��fּj�k=�~=mIE=��E�M��(�<s�t�{�w<�ۈ���L=ⱥ��A=l@)=���<Q�ͻ'�y=�d=P%�;B��o�J<:�F�h���&`=lf2=f��<�57��}��/��_j���K�qJE=ec�<!�<h: ���h;N�<�^{�*y|;
\:<���<��4�`!�;����
��v���-=kW�<f8D=����b:6yS<4 Ǽ�X�<�T�ڃJ=[��9���<�Q=F��P�<�E=�$$�\M�b�����<|����U�<$x&�4�c��<5,���=�z�:w*�(6d=(8�[���]$=���<��=I���μF�<�{�; "<؁=ȻI���=Q刼�f<쐟�5Qa�g������C��ǁ�<Iߠ�֛����L=_}�<���r:	��0����u1�G8n�/�J�s�G=�PD<��#���;n<N�s���=
��=��:�7����ϼ�J�<�}'=ߩ��R=H�7���=N�I=��"���?���#<�<.��<��g���<*zy<�Z�&�3<C�b;���;P��Όc���7�C(T=�n	��	��d��K?����<��<<�<8��<f�q�PGE=�=-V����=��(��p�<t#=�F=c����<���W�l= E廚��f��<Y�S�"�<�K�<np�<���<(��=e�ּ4cB<A��Pjt=fy+�������!<V&&=���xh���%;ӂ}���w=3;x��=^8=� *=�t=z�L��od�ϖ5=��O;W�����!=��3�}��B�6�A[�<f<x)z<m��$����M�u���x�$�%-'���켻����<~b=��8�h9���$�=�<�d�/<��G<�G���ѷ�B�;���<��$=�����)��uH������(9<��=�/�;�.�(�=����V<,񓼂&��'0�<ٵ�;˨X:��.�aՀ�1�<d�n�?�~����P=gѐ;�\<���"�UQ����ͼ�6U=�bR=́��;�$<5�e��L��=�Wһ�R<��F=��*���#=Y�H�m8(=��<�>=���c�8�D�@;4� ���;:��<�ĺ[�k�;�~һ7�K<�c=U�)=�$ʻq򂼋2>��6=n�6=at����=Aļ������<`��<ѷF�3��K\ʻ�~k=>(��W=F�d�@�"=f��n�*����kջ~�.��m4=��Z<DCϼZ���'A=7�P=�<{����^k�Lk4=�9�&{�;ހ��v���$��,<�q =�ߗ�>�<^-�<�==7�����2�=\	�]�;�5�<�7:�K�=FZM<]��n�C<�]_=������ڼ��R�j�����=�w4=A�1�y�ӻ�)I�;��<�?���=N����ٻ��v�Sv=�)����<�r<�N�μS缪Z�<��L���=�4�<�'c��NF�����G����)<	�7=&-�����;�;�c�<�o�<�\:<M��<�4��a=+n"��`=��<��U�!�j�8�_<�@=�$\�]�W;�B��E#�Q�)=Ǧ.���;�V��:�Ѓ=�UB�VK_=����2���y�<����ţf���-=K##�� E=ź��,S`="27=0M߼�z�����.�5��`=+�"=�,�����<�W_=yn�<n 
��<���a��j$�N�<���=�(=�0�<9�,�����b�Q�&p�<�.=�q<��ͼ
%5=�l<r���a>=Bߝ<��:=h�x<��h�vdY=�Tx=y�p�e�:=�������<�/����<��)=�؋��͋=��I��Y��Ò�P�K=t�P;���<W3.<�kk��O�)ZO=�ʮ<�1���p��g	�S�k�*�z�<�$�<>������4���[���=c�!���l=���<��<t��<>��;Z	�<
�ѻ���<��< tS=l�l��b8�t��<�S"=g0����F8�<a�%=��b�k½<�C=lH��BT=���<�޼�_"<���<j4�<ZtS=hz==�#��=3�����<B��N�&�O��m�I�m�0��L���n����<�8=���Q�g=�������<'�6=��8�uw(=|�[��s���V�<PTM�U�<�[�<�[��i^=?:&Ӆ���W=�Se�Ww8�����kA����0.<������Xd=�a3;�#�9'ٻ��&<�ʒ=��J=$Ah�bgb=^w<O.ݻ?YF��NR��9\;���Q��<��<��9=u�V�F^O=��X;�󴼆]c<wi:���;��2<I��<�ܴ<�[2=kߔ<���<�R2=����3s=�\H�3gV=�Z=n \��H=�L<�w��O�T=iE���K�R�`�����nP<&�H7}<��T=�`��g|<��G���/��Ւ��2M�ɏռOY+<T�j��ʋ��b; �v��G)�;>���F����Bd�<<��;d�Ai��xM�<b��<�5����:=fu�v�̻G� ��L=Q���k�>r=9)=οB=`/C=�
��l=*R��}+X�$�:��3}<K.=? e=�4F�y��;<��<�*�;�~���Z�W�=8�i=#��`$=�����.�o-#�N�1=�}�<U�.=*|6;���X�=+�˼#D��.=��<�qV<��<"�g;���=�d=�J�8h�<�2�=
�=ȴ#�L5.<����ES�?�;�; s;�`,5� �E���z=z=�	3��	+=b�;�$=�����2���U=�+żf�U�jg��tń<<>=$��`�F=RD����<��Q�]=��m=F�=��<�\=ǎ^<B�f��V'�P��<���I�����<sE�b�<�1�͆ =*'��T+&=FC��>�A�,<;/���e�;�}?��'Z=WM�8޺�p�<:ޙ<Ǯϼ���<5���E=q_+<&�<�(�;� T�_7<��q�;Cy�E�h��~@��'< ���b1�)E_��=M����=h�F=%x=��L;c��<˅%��S=�M[<��;�*,=i/�ӻR�H(\���J�������=co=>H	��Xڼ�t��̼�o����s=�A=�S�=Z�<�+4=�W�[h=u�Nl�<����'r=�K,=�w`=��߸�Y����A�"=���o3�`�n���.�5Eg=	�<@j�,�o�o:M���m='O=�5!���s:�HϹ+G:�d���<#l�<���DC�w�2=�k";�)h=��=��^�
kf<�|�=$��/
��==��M��XӼ(����82���-ļg�$=I8>��:����/=�C��K��<ڭ=j=D.����;��<�O=�8¼�O_�������<�n��V�==��6��R=�f=Ӻ�5==$=��:��/B=�º<"��<a$=�a��1=5��z8�[(�|�c<5;BĻ<�7=� ���R�<aN���I=u>^�Y=�����T>��;��<b��*h�;eP༠�3��<�F��M�=�^f���m<ℼ��<�.�������˻�9��Sд�n"伧9=��<E�a��:I�ܼy�=��e�*0 <X��<
��D� ��g�;�"��8c�=�=�7=r�F�o�K���(=OAN<�}{9>�.�"��;t|(=G��:k8��7�\<�m=|1ݼ�p���%��=�?�	�����X�&8&�^�R=�t�<  ��3�5;,{�8�-=�1�;�6'�uK�<��%=����
<=�><1Ɨ<��6=��;��]J=U���;�n=3���g��<{�����E=����;L[H�ȕ�<��ļ/�a�9H&=��<��<��:�)V���d���-<�<eV=u5=r[��{o;��;�����B� ��\�:�J�,<��#=X���}-�;f �;��PM<ml��)�Q���<t�=|=�<��i=w�ȻZ74<�&�u��!n=X0<�NI	=���<�����2���2���K�?���I;�A��<?@=v�<n""���)=8�V=sa��G�s��P!������a=�~غ��-��9�<t��<��x<dQ=o�i�Y��;�#��4=����9�4�$X����;���M;��
�&_�<<��;�)<g;��<�v�s^��w�;!"	=S:���~����<α�,Y@��(<��KhW��1�����=���FO$=�-2�P-D=V��:΍߼�{*=S:���;�ё�<1A��\=��<n.���|���s<��K=���<f��<|x�����<��<��)�HV��S=��%=IL#=(���ˏ���ؼ��z�d=_�y<t��6�[=G����!=qI&=6C�;�-=;B�V%&�k�=��������!���.�%=��"�8�#������n+�Em��򇽭HG���=}]=� ���=y�<<�3={�<<>�d��5<"�6���H=$F�;jǼ��:l�;�s��/ۼ8y�:�P�F/=��!=��;w��<�4*�[NK�=�9�
�U=ӣ/�A=Ϙͻ��=`4ԻĦ���μ��;��M=���<�=K��<�[�A�g=��"��}��.�=<7���k�+�<���<��
�C�����9<X=g�<���<�O�<:lE��=N-L=��t�ȼ��<vS�;�	���5=-������O�-<���Q=Xt�=�,<X�f�=&\=�r=�Oi���M���.=*}��%�<H{?=��<�t�8A=�Ln<��6����Ay���f<<.�;���<�3=r��e�;3�n=kN$<�Em�m�E=������3�&�֓;�K
�a=Ǔ��ݛ�<-�����ۻ�RH=|��<��M��\C�%WC��� =K���@<bm���"׼��L<��W=N@�<��0=<��!j�<h,H����9�&�;���1W"���<G�<ywڹY�<�;��[�N_ۼ=Y�:M�߼~A=�@�:�o=��r;�s����޼�9=|tH=m} 9�,����<��~�
��</4l��l�J��aC�T�u='�W=1�=��<A0��˫<�c�����<��!��r=-h=X����xj=\�!�������ܰļ�Q='���<�<&�W��`ݼ�Z��Õ��D�[^;�c�=&A=��X:ﻓ�زN���b�����=y� �����'������)F�Tc�<��.�B�p����;5E�H۰<Xd��\s�Fg=�A<w����=�3���*���<l�9��Au;?���I�=N^��\��<�e��|��?\R���<�i��o��� H=T��<Н��#-����;ڡ��8N��<�8O=�-=Kİ<�YQ����<6�=5]�-n�<�)=b��;֊<q8z=2<�r�&�k����<>����<f2��ڰc=�C�<W��<(|�uɻ-����ۻC���#��mie=��]=<7L<��<��D���=�I}��E=�w �V&�<�`=񬉼6���`���i/<b�M=N�/�Z=�y#�p�G=!�,=�%n<V����<9+�e <�U�=��== ��U0_=�Wʼ$R=�ES<U�X��f�<:�<9�f�OE<�X�<�#=�q=��Egʻ;0���<�P�<6��<�4�<^M:�8�b;�����O=�<���'�<5�<���<�	׼��8w%��i�W=dg��+�;k�;*X=���:=}+y�4��;��o<���]t����=�!����_=!�Ǽ.|���0��3�m�o�T�a��.T$=��Y=]=��;���d�.���ǐ��� �׻$3Լq䕺�-=��<���<�\��+����<��~��-=������V=�= H���g;A�����^=�J`�?�����:���ʡS;�𒼃�a<}�庠ʻ�=I-=�(.=iZ2=�D�g�I�z���<5��2�?�G������<5�ּ�X�gA�~�<c<I��5�u���C=�ף<�H����=�|���8%�Xܻs�<�~�<��g<	�Ѽ7	 =Kk����'<�]w�M�Q�3�ＯZ��U;�{=���=m�C��<��-=�F��{$&=�x=%Pu=�dûm�1;�dּ��= w`<�$<g�6<��ɼ�ө����:���<���]���{�=�]E�y�=�H���;=��=����R�-�C���a�e+i=٪r=db+=A��Y�<��‘;n�"=��:=��l#�<���<�� ����Pi=�= �<SO�8>/[;Gq��!3=8B=a/���;��;XX�H�q;�+�m��<�j=��j�=���<�f���;�(=���]�+=1�;S�A=z3,�l5��'��b9<�6��:�D=|G=�l�<k=�B��a�����=�d,��Ӂ=�+� ,�<#ܺ;��uμ�B��5-�<�3�{�7=$6&; ���g=��+��a�<���;8=��?���=R�P�ӢZ=�dż�x,�8c˻zs�=גE�1xN=ܵD=N+L�n3�<q\"=��<i��I>����<qH��x�紆�����r;���;{�<�.�<h�*=���.<�IƼ�R=��g.��.��ә<�/<=N�j:~b=�d]=<	л^��;��<=<��<���<=�<W=+;�;*����a��A��=�<.��<�h<Wc��WD=��"=�w&=":¼y� =$Pd��>�<���<��߼�#�;Ī��K��%�B��(/�[f�䥚���8��A�C�.=4
���5�����9`ѼK��H�5N=��O���	�vM=�q�=?YX=�Q���y��O�剚<�X-�
<ҾO=�r=0袼J�U=� 1�O�	�f�2�)=�a��=�iP��.��B�$=�'n=!�H<��:�Y�=P��jx:��ؼU��<���߼�����N�<h8Ƽڄ�����dk=�e��]�N<��@�&\A�Yt1���Z=��Ż��=<��t=�Ŷ<�28<�&d<�/!�|q�;d�%�*a��7��Q�<�4�=Ƽ;`i<7ƅ���<�y<�P��=�Zv<����k�ȗ#<v5���Ń��s=��y<���l�<a�e�,�=����;�g
9(jy��S=U��h+�;�μ��F<�l����Y���=M O<�[
=��;�_�<��?�3Ք;<����#=!�|<���!������+���3
����<��=���<������:�Q��,=xͦ<�G��������+=��=�*���?����=��;�㼶+����ӼP�<=(�мT���t=8�d�e��<�Վ<H�.��TR<����+|��7�<N�c=j�3������A<	�Y<�E!=s�A=�׭<x�aD"=�'< 5��ȸP=p��<���<�]���;L�
q�q��U�,=��<Ԅ�;[��<�+��y>�kX�h=�u-=�I���~=���_ƼuD���a���{��-�0l���lY�=�N�2=���;#��=!��/?�<��:�X����<��;��y�N�����;i�b�!6�K�<��U�n�l=������<+\�<��h��Ph=N22=���<�9����;Q-�¤O������=x�<h��<$�)=��P=�5���<~��f��<� �D��<W^��J�*��9i��ȼ��<v]Ҽ}�= K�<���/�s���
����<dR��͗w���<	VB=��=��)=�U:���;�(=��Ҽ*᷻�����Dۻ��a���=?��<ub=�Y`<�>=B-f=�A�;8�$t�<+���Q�L=Cpf=m/=<�;Nk�|�$<�lk��=�
=��]=���<�����p=91��� ��8���_���������"�~��<��,=���;��S�ؼ��<�Ǽ[��<c <�;'=!�?�w8�W3|�<k.�\�<E�{<�<�<�3z�*V��_�"UH=b�M=l~��f[=����"oM��:/�=�<r��9w���S=�cI�F��t];r`�<�ހ�پ :T��;�{=�Oռ��'�!4�\f=4�Q=�x���鰻�#4��L�<S��Y���	�p���nN�u]��B��Z�Y=Ǆ�<�� =o߶�9�<��	������!=b�/��ȕ��1��-��E�<�rٻ��7�Sv�<Y"л&Cؼ�3�o��C��V?����)�=Q��~F��;��������üu�t=Wp'����#g��#�.<pX��*��<"���	�<w!�<"]�;�@;,]L<,g/<AQ��>�N�ù�p�m<��*I����#�ǽ�<KtѼר<���<L�=�>��!����<}T=���;,�<�]<q���c/;�W�<����}�^=�}`=��U�0|/�@ǐ�+�'=��_<žT��<c=»]=���<��C=G �<^*��&͵����D#�0��W�U�KX��:�;̄2<v^f;�[=���~�;+7=�68�s��;����D=��=�ℼ� =�I='��<��*���=�}9���!�M0��f��H�C��/��P:!��t;�)�<U�'��=����t�<�_�&��4=��e=�;�<:���<�[=����ټ���<�{��Pf%=�6=���px�<��=�-K=F�<�7 ���f=��1�::�e���!��?����L=�לּiB�<�:�Zd=?�="�<���<	^0�!S �>$����I<�=F�����=�YN��S>=��%�N���>���=�v�<&��<�z��֮��0X��������C>�"Q���	c�P=��=���<�XϺ��Y=�[���=�[�<Pk����=�F�<ػ���;���Q+#=�DZ;f�=�=���<�Sq<'z�<
x��M�&�	������(?� KԼ�$���}<�u��4[��t=/�H�z,T�x�<o�<g��Ѵ��r[�<��<3���ŕ��
�@=�QL=8������� ��{�=�6���=ߋ�<}a�Q��<�<���;=Mq;�3��:����O�"�K�,�=r�r<��+��+�<fS�;5�x�f;��=&W`<Ŵ�7pF=-�޼I���e���<��'=>�=l�мFR�g��<�Y��
�<n�:�o�+���,�f7=���J�; !Ӽ�/�<�Op=�˼�y=�`��m�<���<8�}�s-�;v�-�����¿<�;�`(��c2=V�0�<qi���7=�;j&=�k-=n	���1��~����/�+\�<x�p=/�(<P��9㢼��";��F�>b��|�S�>=�t������;[�<#�L=� ����:��1=#�=|�
�E���!�.�j��0�`:t���=��|<H���o�i��NE=��B�0���C|�p_=��_=��<�>�<��3=A9I���<�#.�^˼�4u<�C�<����o��:��;�8Q=sk_�b��P��<�Y=�&;��P<;�=�ۇ�9��V<%|�;,r���d�Z
��fx=����0=�i�e�<w7=��=iߌ�s<��v�'�ϼ�d��b�!;��[�;�(���}=�9"��&G���,�$��<@ȥ�nJj=�=��<�u=�Y�<�k�:#J[�e�<[)�������<
�=&��M�M��a�C�~�=�7=)"�Փ̼�ze���b=\x��k=qJ�<��;|`=�w�<)� =0"�`hV=�&O9ш��P�u
I;^���=\&�����hc�kr��mP���e`��߂9�I^��B�����wґ���; N��腺.�<��9s+�!k
=6Ї</^�</8�����<[FI<?�U��D�9nT=�{e<^Q��E=^:�=IF�����PiڼeC��+��[�<�G�;��;��=�H܌�r��}�,�*���_�=9O�2c�1썽&�(=}�r=��9Y&�������=^���Z������;y��<��
=�/:'�@�p�fP=�H��⧦��@�<^�t��:I=O�1���������[T=�;3=gb6=s�k=��;w�ؼ�J=J�C�~<$��=��$�3����<Z<I�-g=�#2�
8�����<c�8=�q<#��<�덼������=�;9;zx<竔��IY�e�=�v.<ԑ==zP�k�;�?��^�<U+=2>A�'�H���x<�?������:��<��<6Iu��i9=Cm;�:�<U�����<�g�<��t<9�b<���Υ�<�
Q=��=���<ډ'=�.��D{=�=���=�X<S�w�;�l=/3��K<�R� J�/w<�?�gzx=��C<��3=�5�V̰<����	7���1����#<�b����|=*�;C��<yQ8����;ƃ�|�*<�ы<���	���<?�ϼ��2<!��/7s=�<���;�/Q���<�߼m�<���<Lt�UM��ȅ���7��ة<�UO���?=V^�;"&л�쨼"��%��bp<<�>=�-�<:�ÿ�<;�⼵\|=�B=�^�<ܟ=5cȹ�i<L	=�7=��߼�:����<���<c< =^׸��S+�����2~=%(<�#%�dN";=*+�Z#��s�<_�3=Yi���8�<��[=j{K���a;��߼�.�<�̼]58=0ٸ<�U�<�4��.��aw=�/;c�<8�[��&=����Z��ؼ��*�$�=���������� ;<�p�8�DR��k�<h�N=����7�Z< ���A�=g�?;�@�<CB[��u�<�N�f'�~UC�=D㌼]�����MI���*=g��;�M=�:K<��#�)b=�b�u6=,=(�"<�]=l@J=c/��P�<R<Zq5����<��,=��6�Q9v<�; =�"���L=�iP��w��§<>���=��~ü��8��뷺$�l�:}�����<��;��}��<�&��(�6F���.E=�X=��ü_nO�Zi�w#;�<f���Ʌ�EXA=��r<+�7�sܨ��w$;���<�p#<�$4�LI�<��=k����鍼�)U=�]6=M9=]w8�b�-��@=�/��~�=�޹<'Z�q֬�(ּ0e1��}�<OQ��䎺B�e�����ů�<̘q=�4����=k����<qp��?L���<ǐ<_� ����	�1=�¼�/"=������;��G=
3��}1<�X�D��<��M��Z,=��a�\�<u�~�9��<*n���?=��&�B��<��
�ݦC=*R:h��<�м�w=�Rc�D8.�i	?=[7j�]y��o�[���O!=6�	;��!0߼�;
=������ټ-=���Q<�~!�~�#<��'=<=��Y���%=������o��́<qR=p��=5�]�Qtۻ�[1��-=l���y�l<#��<�ŀ=rQ�<6�ܺ0�Ƽ��,�_3�@�=��!=6+1�>Y�<P?��+H=1��<T�<��L�pJ��H�\�o��'R�h$=�1=#�p;1�s���<^����q�i;��G�:�pP��N��l`�<<_�P=%�F���<l�o�=/+�_6u=��7=�J=+h>:�e<�x��Kme=��p��a=��n�`Ba=�*���,��t���TB<IV�<Yd[���y<�ru=��4=�ѧ<.2C;�ͼ��7=��c��t)=�==D��<�G?��(7�ԇ:b,=3�Z���v=��κ�l�Q�����ׄT=`tQ=揻���<ƣ= ��<�&j�Z�5<��;�B8���ϼȘ�<�i�/2~���ܻ�`��[��ۺ�`�;<�L/����<�d���7A=�tI�s���`�<�P2���M�w	���<Qo��d��<�
���=��1=_@=��0=�{b�/<� �;Ec��Elc�:�
���
���=T鼚��w���	�x=@g�;�U��|p�� f4���L��=G�F����<q@�x�<�����r��As��g4�������<�?ۼ�$�e�6=O�Y<L"���/=�0g=μ�;��R�<ڰڼS����Ar��|��y#A�)�<��};ao�<P=Q�<Q�J��;N�Ȼd��;~=�<���}u�:)�e<-6O=B�=SE1�}��V���a�=�=)�<Kx5=Ƈ]�R7�<�I=���abj��qy;�o���1���k=4��<2�d��8;�j���;���޼9��<�L=�H��.^�k��Z�<M2!��y�<CB�<}Wu�� =�M��<�z�(���<?��i�X�(�4���i<�<~jX=)";���<��)<a�z=�&ۼ��k=8ZZ=[7���u������`��H�o�;h_;��ȼ��p�_�t���.<Z4=fjs<wJ�>v-��]����#�t�:8ۼqw&�l]<�G�C�J��C�#�b�c�ͻ/aZ���T����1�;��=��O;�D�<%�T={��fN=�\��A=�r��E�X=#Uj<�:h��u�< �x;е��K.��1s%=��B�������=e�绚�@�<t�P���ҿ�=}D�,=i��;�Y<��!;��M���y�&����0=���;#^(��� =7s��L��t2�<��.<��]<eC�)ͼ�t=��=y-7��9�Z}<m��<Cx����:�޿���o��R�<VC�=-.��̄=��s<�ȼ&�<��[=_�3��G5�����{y=�.����H�;���v!K<zZ=�tn���W�7��:2��X*}�*,*��,���7������7�fd���<�B$=��U���9&;��=���;�<E��<ж�<l÷<ԡ��c�v=F�;�#u�ro���B>=ݖ�<��<.f�<G�4���+��->=J	ļU/�<��=�vP=��!<C�=*`��e=��<�`H���P�� O�G��M�����<�H�<؄�;5�ȼ�V<^ﵻ��f=gC�<隌;e�3��_��Z���TƼ��L=�#�=j�&=�W�;�B=s�=ս[=0��N��аd��hռ=�N�I����o=]X�<����q��\<]��z�6=A
��饖��(
�֊+=?�'�":�Y���<]�< jP��e�<��=i���h�<%&�����q= }�=�|g<�A�<��q���1=@s=���<��L��,=aL�:��R=��'�ص�Ҵ�;=z=���<!8�<��L=ž���u�����:TB�;ݎ�3o4=�i
=���<�J����y<�<���<��=�A�O>���c=2_��qc=��<c�p��-;x�#=;�+<dd9�*7=Y�a=�n<b/�;��W��}�CMa��k��{wＥ7�=�y�<ۧ<!\)=�C^��@�<'3�</k��8��<l()�<�v����jA������<�=��<�OB���<<4��9��
�<Ư�<m�<DiT��砼M6}������E={�=����Q�U�q<?G=�B�_`i�!�4=�s=��Y<
L4=Sl��,�f�]���;��;�bM�%�	�;��=3 �<������=,���/S=�8!�U���e��Z��]�^=#+~��y���ʼR�m��물G�<:���Mӣ<�޻.��F*��5q=M�<�����D<S��v�<�`�>��<��<�3r<QS=#(�%g4��%89��<=X�;��=9k:<;I=)��<^�I;g!�<�O��L���`p=l�=���;���a/����<^���@E�m��Uv��))���<=x^=e�\=��缠^S=]�n<Љ�<Ό�<Db��{��<Ho<j��Gނ�VSu;͞�=�<=r�%��'=��F=Mf�<�+u=(u(�)=n9K�񻎙5=�w���$��1=���;wh<#M~��d&=�zy���i=5��<�8C;��.===f��%��|����<jTE��g���I�L+���%�S㏻�=�������+=��3��t=��x=�~���܌���;���:�PDz�|U�<i|���SԻ���<���?�<AZ���<d�����<����S�F��x9�*S<T�+�G�\<
=�42=���Wނ<�x�<� ʼ�_��u�B�vg==�����֤�:�Q<ayq��~,=	E�<$�W.=y�V���<��=�'�<w?���$��@ �Tի<�;+t=�.����=1����S���<�d�+���˼9Kv�����q=�8\=2;�<.�&==A�<�\c�}K3�XAo���;=��G�:��;�X=	Ȉ=/�)�ܟ ����_�;�$=K��<�ĉ=��=�^�;8�l=�t"�K_<�[:='�"=*�<�n7���=OȺ��U=�=�<�T=����X<U�b<��:�7N<�����<pMr�䩼I�8=�h��b�����E=��~��8����<L%\��2`=�
A=�=<�<��=6W>�)����¼'�=Z���ׯ<�c��yq=N��Y��<�#/�vл<�6�=Ն<fm9=��<7͌=�"�<O�<=�2Z���S�SuF�r=l�*���<)?�� :�x�]�Qž;� =��v=��C;��˼sNڼ��<��c�h*E=�pj;~�
=ѷ�;-?߹�A���T�dW=h�1<�=_a�=
�;=��(�%�(ʾ�l�=��3=!=,�<��\��;�B�c����<����s�d��<��w<���<�GG��g���m`��Y��m =��B���s���i�'=7�<u��:�yI�<Q+>����� 2=��>�q����PV�q��
��a�<]`��<��$7=��&=װ��_X���=;��=��<[H)��*��e�t<��t=m/���H�IR�ݩ`=�MJ=f6Z=�Z1<|�<��Q��[=�曼R]<����<#=J�<75��D.=���;�<<X^��e3�<=tT=��i�4�=�֫<H^T=0Q=��<��i�,�N��=�l@���3�<_jq<�Dd�(g4=7�Jr�a�.=�Si=�����o�;N�d�K=nA<��5<�a��(<x��<&�w�6*ݻ\��H�H�BZA�K�Z���&=��=��==y�5�l<��;V]���#��]�A<�R_����8��yN����Rf�1�U�߸Ἱ;=��=�iU�5���P�"V+<w~�Њ8={�<�.=�;<�R��ڍ<4AǼ��=0:�<�v�<X���%\̼��o<�<��HJ�ߢ�<D�ʻˆ�<t�Z�TY����<p�»x5+=������I=*���,=���<`U-�i�~���^=q��&�<1�=��^<SU;��M�S<=(��QT��GT�q�V�e=}��<��<��_=.?�<��C�u��<S5<
R@=5��+��	/;l�<��׼ C�Z��<����B�Ni=��x<q�;=)�=�!!���<����R^>=�Ӛ<���<&���A=Z�k��|r=�$����<���<(q=R�͂7=m0�gXɼ@b�<� �<�=�]�=�d?����X@�;oQ=^�@<�P���<����HJ=/�F=�s���p�<�1��;�<�ԏ<]aS��f�ORF�IF#�9B`�Ø<_����=a+=A�U=��fTҺ[�������w6=�Zͼٝ,=/q2�ox�r�f</O�<�)b=W�ɼ�7�+8<=[�=�w0��^�G�4����n��������b[B�(��O��.=���2Ņ<�+=��D=�9=^�Q<����C�'�[�W�,�<*~=~���b=ƺ؎����q;?,n<ѻs<�;Ѹ=W/�;ů�<n�;��<l�l<��5�j��<!=��R=?K����{;-6=���7$�<�-�Iu==��I�o��=�[L��>}=��B�.߻"�&����a�<��@<�幼L$<KU�<^�:h|�;�;��"<١Ǽ<Z=E0��X�1����;r�=S�Һ	�2:��=`\�V=1���0<�f=�\�OP���<���<��<Ny4�úQ�Y��<���<gM�;j	�<�Ʋ�ѹ��
(������X�j��9+K�<{����@=$Bc���Z=X����:���"*=Ynn�`U�<�oa�8 Z=�����&�j�ǻы4<&3=�b��<�e<����SB�]2��H��vq~<�;k�m���<���;r9�@�#�-4.=���No*=׼*yb<.�(��<��n<Zx=��I?;= &���=U(<�V�:���ѡ��@߼p-P�_=+#s���=���1μ��<:�u=�x����<T+�<
$�F��<��<� ��'�<}C-�����XN�C�n�+tм��T���:r=f=X	�< ��ă�;#l7����<��Z���x=�ܓ<���;$��_Ni<�0��P`*��%��F�7=��������;gX_=&�;��@������O=��w��N=o�X�]�>�Z�<Am;Xm=�B��G<.-K��j�����Y������!&������2�7�ü��<��:z�e��H<.�O=(�f��F�Z�'��	¼��m�>0�<Y0=�P�����)8�;����kV<̦�/C���<!x<\��;�kc=˹<R�<�CѼ��=W��x8;;R�����<!b��X�<P��D<�p���< Ϭ<X�A=_=�H����<kr<�{/�q�<�r�=M�����;�
=	�A��_��6����<?GȼnJ�mLJ��WĻ���^�$=�Qg�!s�j�;4����@=�c=��[��
�y��;B\j=��-=l��<��C���;�N=G��<����(��</Y	=/_̼uD=�3���
��<���<��p���r=E� �bK< <��<Ⱦ���r��	�����I�K�26=2�ܼ�ܼ*ڻ�R��9��k�;d��;��l=Ez[<��&;i���!^����=�]�<o��;�<=Cq=��q=�}�\�l;���<����)�H�X=�"C= �\���*�{�?�0e-=+�^=������"|_<g��ZK�<#��<+���)��VK�</�=��<�x�mТ;���k}���<L�L������<U�����6�g�[=2B�<����U+�ri<���=� 4��7�����
k�;j�X�Y�_� ;F�;�.���ǻ?�b���3=�6ܻvp=����B(P�R�����-=U��<|vC�2|���`�����i�:�U�;�Ү��FL��à��D?�l�8��)T�Ӄ��K]ҼB�)=px=z�<��G��^�< � �j5i<�Kf�P��<��<m閻�S="FX=|H<qs�<F���(=�k<�=��l�����;n-�<z��_?�;��;���<�`�<n�;d�Z�i�d��Rg=ƻH�{<���H=�E;�/iC����<$��������!N=RN=,} �av�u�X=� ���ڼ��9<ᘕ<��(=��<��=�<�� ����N R��>=����!�<b뺋m�<=�=s����1S��AP�?jW:��e�D�=S���I<}}�a_<�0p���;Z�o����:�l��D�<&#�<7`鼍*P=����$(=DI"���T'�*pW=�
�=��c�%=M�(=FD���h�<m(���&��^�:U�/�}=��1;�h߼�蘼����=�.�;����g��YC��==��.������F�KM����S=�:����`=%42=���<]�;�3j=* ���<��)=�==�H0=���;fk��@I��l0<ǄC=�\q;��5<��<�i�<R�==���;��=UB�޲�<I�4��6��1K1�h�X<�=��H�l d<aa����f����<0��u�<�i�<��7��<�`�9KxU<'�ʼ;�O���1��z�T�g=�{=�{�"*y<��=�?0<3�7�0w�<��#=>��:(q0��(ܼ���^�P��`*��B2=k�	�*�y=T	8I��/�=���<�m�<�R��&�;3B���d���<{$e����V
2���K=�`=���=��i�
[���x=5|A=	�iW���,<P��;TbN��3�<�=G�i���N=N�5=�O�>�B<½U��M���<R�X����;��H#C=4�M<վP�z2b����<�ļБ�2&=��ļzA�3&=ƍn=Fd���1�<H���^�M��aݻ�G������j��Y.��o�
�N-8=��E�x�&=};r��i�i��<Tf�<���]�p=n��9o<�F=���<� =�_A��h�=�{x�%QE=8���ˠ��]ؼ�VI��{<z<!�l�<��B��^һ��(:;	��㲼?-Q�J5 ��0�<o�Ļ7�<�K��]�=� =|��+��>��<�+���R<��`��b'�yq�����Ҽ��j���2��һV~_=��ۺ`=��&�_A;��w_����
P�;zs�&;^<}a�DX;(X{�Q(��1TK=5��<�47=.��ڤB������ =�粒����mD��t��H<§���vI<c��U����:ZT\=7�������8�<4��<3�ͺw>�<�֥;�j��Bu=�W�<h=>x;|v�<5��<�H�Gὼ��U8"=�=@�5=j�=��V=�r�<50��!a�ʂ&��,0=�_^�ѓb��?������ ��J{0=&���ۄ�P�b���o��ן<�¸�8+Q=ַ�<$���ŚK= ���Ar��$�R�ǳ¼�t�<��T��O=�=5��ѽ<�ܼ��d��q�����	֫:]T=/��<T#r=~%=C�+=͵�=�ʼ��Y=�{!=��3��eк%��<|�n���p=!�'<��<D��:�-=�w�<��.�h�_W=��!=�9=j=�����⁼>��<�=��;��Si�oˀ<��b�$`��.�<���;D�<���<�@�<2!=p<A$5������	<" ��v��P�<oO=�[=��Q;|��<ߊ�;&ꏽ<��<�u�Z�?=78W=إi��	=b=�����R�N��/=��r���E�4^=����Z<�[��_Q��i<+v�t�l='��<9�m񼅀q<���_�����`[(��ۑ�6��1��<n��ED�G
F���@=c8=�� ��=?���v��2_,=�<ҼX�X��4=_rg���;B;'��@�d3=k�d��=�(i=���<6Ģ<E��>M�<A���><����C���=��=nY��
�j	λq6<)f�<Cٺ-��*O7�-¸<�R��J����� =p3���=��;o�-�{�<c�=��;c���`�?=дO= ��%؂��� =d���"5T��W�<Ѵ�g'<\v'=rA�������X�3�)=������`=~:=I@=䟅=�#�<=6���ֽ��I=�K�<k��=�C�<��2���I=]E*=�ż�~��:=�����h�<�nt��6=�K������;�;u�	�<���P*=X-�<^%Q�N��;�>1����<�U���=�=�_:u�w��V��=˖����U;��FV=7X�<M���l�<�"Q�zM���U=�%Ӻ��"�f��;hhg��N��\y <��<��R����<p0=�dV��.=5��Q�$<sf$=k4=�J��8�| �����b�𼝄B��j�=<|�;=�<ҥ��¸<KػA5� �-��1={u�<c�Z�F�
��̻9I���j�<�*�=,R���Pu=���;�	��<��t��=>J���_�MJ��ߩ;M�<5?�Ww3=r��XX�TN�]��&e�<F'=�V��}<�X�"�`<"��<I��0|<�s��g�!=���<��%=7��<�,�<J�wr�Wd�4�=���Ҝ�����<�!T�Z��N�©�<k+����H=�)�<�x�<����C�*=m4;9���<�>��v]�d����^!��H=ֻR=5<ml<��?�<��+=��z<8@A=l)g� �l�=�=_2�h0=�9������c�������Jr�}�}<ҵ�<��0=3�;@S<�*���ձ<�k��?u<�I"��Ӽ_�f�s�I=��T�x�@r�<���=N	=���<6o�9����y4=�Y=Hּ:�<M+<�g=��.<���m.��<pM7=��	��ӓ<�v�@��Y	���8�C�U��߼R�s;��*�<��H�i�Xc�L=�=��B=Q�ϼz���Eh��v`�ϑ=�6�<�!�;wW��T<���������<���UvI=
4e�*y/�;�1=Z��rB=|*�<�r�7��<�~�<nx�:���d��Y0W�Q�?�%�W�����|�{3�<#;<x:�<l$�<�l=�x=���;� ���¼&�.<q�+���H=Yp��v����d<�'<0�D��	=�Q��2�Q=۷<ƾ�����N=?6�< (k�lW;=N��<�΂;��c=Ȯ3<�@t<������4-=0�c<� ��l[;t�fD=5DW�y�<sN��hp=!A!��K�=��M<YUм��<E�\=�м���<,�G�������*=�=%#�o��=R�ܼ?�P��U���b�;���s��uŻ1�����;W�<�ڻ��]�D��<E=_=��+���<ɺ<��3=�A�o����=�IE�p=��(�5�6�-L�=R?�=C�Nd��|�ڻVQ.=Y2���V�ⶺ��e�/=��}���F����<ċ���D�<I
_=wI��f=n�ϼ󈼍hp�76���
=M���"���n=�k���:_��<brE=܋�;����w �\���J�<\h�<��<�]= ����0�=�W=V�ڼ������<�H%<θB=�$����|;�
z=�2¼_xG=^�x<��<����Y3=�>=�xy=?���PZ</�#=�Rf�jK	=0#��hh�� <3U��թ=_��<�8<a%u;��9�}B���=��_��g�;�2�;D�b��=����+b%=p�=�pHr��>C=�@P=��g�^H�c.��{���L��<�s�<�G=��$���ȼoCQ��y��#r-�2e:��;���;� 滞����U�b�$��/<�X'=�򢼗$:���e="���$�;�5�������!=	�ͼ-��<��=��(��tv�v��;��5<	Ǖ<�� �Ms=��^<CY�<���<�#,���-;λ=�
�<#�<�x7+�н=�����z�<�`A=��|=�.�;�6=�s=�b���i=BS�����_���*=�C =��v�����Y=L�A��.�����; �O��m<�5=���y��rK���=���<��;c�/�+=�r�,z4����<��+�c�;Y�\��R��'X=��+=o��;8��<晊<��-��(=��=��Vl����=Cim�{�=w�<iR3=h��<򹧼B�U�p�t<��Ժg�2��^�=":k�<+�]<�E@<�:ݍ�>vi=�[,��U<#��<���;u��<�1��Q=[9�;��J= ^e��l�w�P��>?���X=o��<R�-�Ve��E�'�<�;&�<=��;;�����j!<bT =ߛ[����6�<�kP����<P��<�����=7/$�͝���g�<[�=f �迎��K<?%#=�p&�l0\����WI:�'�<F�v���s�P�[=�=�E7��e=�Kf=��ʼ��=���=L��<�-��c/�� C�D����3���D<�
=��o=�n�:JkL<m�������yB��j�U@�<X�=f<-���<Ĳ=x��<F&�<��%�6��<����]��<��<��ؼ�?����<�h,=yc0����Z�<J��<���<�X=h�K=�!Q�{�}=�x-=�II��7W�·���x<	�d���4= h��F\<e�^=�vѻ�������顂=�KJ�o����=��b;e�5�5�=ɟw9Q�W=��;sњ��[� WE<��'=K�߼zR=5��̖7</u=���<�����c���&��,"=��<��h�*%�<p������X<�0<��+=�^�<�{�z�5�~J�<��<?=W6�.\�<���<�~�Q=���;S  ��T�<[=
iü�*=g=<�I�<��<XQd<9N��$�<ii� +��x������Ϻ�<��E=K`��Zx�:�x=��<�6�:}���}
=Й�?�&��쉹4���9����j<B!�o���/��c����>��iмκZ���Z�IC��L���>�xH5=�7B,�c�)<��3=C�<@�j��<L��<D#��dE4=�ͮ���=��=Y�j��˧:��6=�������	�[=��G<�Ư��WO���<Xl=�~�<}X�!(,<�����)<���<����4�H?��~?�ڼ�'ջ��,���cQ=�q��-K<��=T��g 弦(�����S=��A<��h��C�;��)�{�ûo�<L}0�^^=���9���=xa^�æ�;�S^�z��<
�q����<Z)=�Ϡ<o��3	�ftf=�݅�.d�;ss�a�?<�ռ<p�<�Vq�@�=�=,�,<P��k˻)n�+�=����Ca��`����<Ip�<����Xi����]Y-�'i=��_�^�<�?/=��<��$=��;���;����&��<�Q�;���"�C=,fT�>)u���<��3:|�G=�79<R��ۼ2��?Cn;5��'����}���;d`=��~;�R�R!����P=/8�B�;=&�S�M��8B��:n�"=�.��2m=YW�<C򦺌�ӻI==N�m�Q��<[��	=^(���L��n^�yM_�3K�5�8��X;<��=ӯ-=>�Q=}@M=S�!=��M="j��s�:�
�<���<��l�V:�ՖV= ��<fM!=�tV���<���<4i�rh�<��;���׼�MJ=�P=e.=y�9�%h1���<A��oZ���F=��==b�6=6G=n��;�=�ᚼ��E��l?��\߼��<x�V=x�=a/�<�?�q\�Q��:��U�x\<]f$��,)��u�M� =ogx<w�E=��k=�lG=��s��Au�j�P=��2=�~=�����<��<=�\=�=�K����<��U=pzJ=���<�殻O!W��~�=ht�3����=os�	z�:�d^=�(y�ws�<9���+=�5
����t��i>����Y��<�/Y��N�����y�̓~�U��<�f�t�<Q��Qp༲�	<��X����*=����2w;����U���¼��	=��<��zA����<Ż��R=@h=��.�鼽�=>�[=b';��؎<<�O=r�ļ�d�<-xO�pf�<��^�3�r<��
�N=�==ہJ=
��<h��<V��<�N�<H�<[DW<�X7����<t�V��eּ�(4=BAj=�:]<k�+=�軼{֭�q8�<Z@�<i@<eS����Ƽ��R= ��;4=?	�<�K<=Te���L1���7=�;���<߰�5֋���]�"��<�=�~/=.Ub<������<�6$�Zx�;FF=ҷD=w�L=�r<�ܼ��<K;P�	��<�2g����<�,<o1c�+k�{ ��l=n��"=�<�<����9�w;ܭ��iI���N:�%�E�I=�X�<��:=G���&�j;B�����:����<&I=*�Ǽ�z��;���:���h�����ƳE���<�W�N����R�<ip��,E����=71*��B=�L��Wv\��Fu=b2�<C�Y=������fT�<SI�<�D0�G0b��d=<��GH��C�����p/=�9�<u�\�&�G��a�C��ѼZ(�<p�<>��<�O��h��cF�< Im<N�<��<� ��廇�2=�Ai<S$q�+߼­=�)a=�<�<��L=��$=$�=�a��}�^���#�� ��_Z�:����K�h=�z���</~��:�%<�Q:#.z=�V�<�&
�s<P=�a=�7=�>Z=k�<�<p��]
��m��r����:� [���K=jy�;�F�n*=+�ۻl5+��==�r�:s߼4��<*!=L7���'`���N�2R�8P�U=�� � ^弁�;(X��aq �cl]<�=��[��<:�<zOѼ%==�I����9�$�/=v=���;A����7~�m�2;���x�<i��<��;1�.���>�M�I��;d��T�=ԙl=�:"=�ڏ�"~�KS��P,��?�������&���2�
Ʊ�Ժ޼�HE=O.�>1��r�o<��J=�*E;O�"=����=�GY�p-�9�_[=`͡��� ��<B���)=��v�1|�;Y�O�)�=�4S=J�ݻ�
���C�.�`�K�Z��=���<�㉻��=Zt;M��$/h���=���N*<kB�<^q�;U�K�<;��J�5C��:��;�<N B���wF</Tr��/��=��ͼ =cK=��\��G� ��<�>����t�f밼�G��J�>=%�=��f=%I/�A�U�K�:8U,=��g�u���D�C�W	=XY=�!;��U=0��<��-=�G`��0�d=�i`�U����<m�#=`�<�´��o!�� �;h.=�v=��d���=T_��)�<ȸN<��9|-ٻ]`�< x��zO=rh�x�E��l�G�3�,zO=(��<"�ݼj�<s�=�!b=%�r�z�I��Wb=���8M��?� �<^0̼{q)�]
=AR}<G�7��0:����|��c�<�^=6�[�Q��<�PJ=�Df=OU��T�"1"9�z��-=Jo2�?��<�5��a+�U���(p輑��<	OE�4���<�<g��=��C&��_�5=Ix<��O�ʏ���e8=F�4��@��@ܼc�G=o�I���8=�X����L=�+c��4���׼l�J<bQϼ9�=nDV��U�;*�< a��^?(<�S5=�P�Q(!=	��Մ<��C�<�f�?S=bF��;��/��H'�u�I�7�e�C=��=_��?�9[C=M=�%=�)�;���<q�q��E�<�|�w�i<
I=t:�m�-L�<S�<E�W<U���S=�%!=�i
=�!d�8��;0_�=v:H�R�ܼ�pp<V�Ǽ��9���6<����j��E���g:9��=�xV����g=�c��-�;�+B� vS��Uk�t��Z�2��Q%=���<���+����v=ݮ��	�����=�x9=F(q��h3�����)�<�b=� =��<�Lw�۟	=�=�`���Y��x>=UUO=!��V%
���=mi=I��2�=Ъz;��b��D=O��<�)�׀"�œ �#o�;¡1=��^����<;�L=��5=$6n���<|��<�=~�м#S�us;�����=)�!<	�6<�-�� v�Yrƻ�?�g��y��=�����Ba���1<���Y��;��GL׼$X-={�Z��oƼMqüia=�)�<�5�<��E�[-�<nh< ���=%�=��<��ѻbx�<j7=���J���oY=>�A��s��&=qJ��H�<�M�;�O�v��<m�F���o��P}�2&a=Dq5=E���4�9ϼ� ?��iQ=��j<�<�B=��=��g<!/����� g(=���:�<=Mz����¼��;�<	��p�;������=ʿ�=
�<��	�+�r<�<|�C��tܺ���4#��zu=�?�Lk;�J= +i�V���ݭ������A;0I��	=�w�����}�<��0=P([��=mK=D#�<$��<d��< ��ػ���<�����a���<�˻0L����=@}����<
	����Q�	}���<�} <��(���:j<f��2v�*x�;ЂM=�� =6��:]1<�C=�T>=�jQ���k;���S�%=��O��Rw<vW�<}`=������<k}P<h_�<��+���"=�*<��׼�[:ld=�~��y�����<��<���: ��<�*=������F��18=tb������ܥ<g��,���V���4<�]j=���6U<_��<� =!É<�&=�(!����r6 �r�f=�I�<�ҵ��<�r}��in=�K����;�n���w�l�M=��<�(ռ�$=���S�$u1��<c=^�Z��` ���b=�'��<�=)R�<�P�����a�;���<,8��8�&��;��T�r����;���<V�<79���T�;❼��<J��<h�m��p!<�)�<��t<-y�<��<Q�<g�<!Tk=*d��y<=F�5=��Z�)�w<]�0=_��<��2�1K��т��]��=�b�X[�<��üA�@��R=4��;����<~��<�OüA@���$�J�\���<�o�<Sݼ�@ ��)����vX=�Fn<�孼q�	����63Ļ�Ơ���|��,g=
ޒ��]�n~�:�^�<hX=I�H=��\=x� <�^��K�����;����o�;��L�Z|e�[WQ<h��7���$.;�j��IǼ�n/������<��-=EGx�{=sOB�^�a=�K=%� �k�h<��y�Ω<{=@����=
=��߼��= �Ӻ�\�<�!.�<y��*�w|I=f{�<�Zj<q~��VjX=�)=����"Y�'��;z�;��P��79��dV���;<�"l=�bD��B=�G1=�R���)�Ee�<��8=H��I	�<�j>�B�=xW�l��;��?�M�=��A�����m6a��`�;ȶ ���^= �8<O�=P#���c��>�����,;�~%<�Ȼ5�;�	���;�*?=n*���	8���Y=��<�(=:�ue��U�ڏ���P�g� �"����9A��Ϻ�c;��=m�<z �<��m;��߻FWl�&]�:�|�<�<`�=��H�b�<!'�V�<�]-���[=ޅc=�I�������:=#��Cg����Z�i<3K\<nLB=:PN=�g���w��Z��q=a;\=@�<��d=���K�w<��y<9:���=��3=��ͼ�O8�1�s�1�;�%u=:�<�蠼�cz�	�Y�ej�Y�g<�B�4��<�K/:?���a���u<��#=��e��Y�;P=;=f�d=h�7=��1��K=��<��
�K��<�� =d3F�����1n=��T=��2:y��=oFK�4<��:%lS=>j�<�蹻dU=^q�t�y;� 7��;=�����ռi��PԼ�or=O=��=�˥<r�(L=�7�<[�_<��;�#=]���<=p;^�$/������ ����Ƽ���w�a�4/���bܼQql�����v���V�<�V?�u���wD=0�	���=�5�Aмt;=��<��:�I!=��5���$=�DS=Ka�=�&V=��ڼ��P�0=5O=jc=B��<��&=�=����E�K����	9���J��A4�Y�J=�t����w��X�@��.��Ӆ��J=t	��S��.��f�;�uL=�0=���<�>�<$�<�~f=j]�<�����8=(���-�<�2(�hZ��Q2��/=�=Y=�is���!��@I=�O�<qS=�邻�Ι<�)����
�������F��j<��Z���y��R=<C�;V�f��y1=��s<}jj=��<6�I���=��;�7����t�f~1<��;�[M<M����<6�"<���F��<�n�9G�Q=X�5=�ǰ�CN�:�G<Z��;�v^=}U��"�#P��f��<tB���<�$+��hf�\D=�	Ǽ��Ѽ0���k=�ߊ<
c�<�c��4�<;_=�ap=L/'=�<=d��^I���m=��~<��q�k�$�yz켺U�<!�(=�<*�F��F���.=i�o=���dʃ�~�:=�g��R%=��<=�� =��U��y)<S�+=3V�<�ZV=�}<�z=���<�<s�:�i<9����_�<&t���?��(�< =��<��<[G+�|.�;)�1�5����'=g�;�q��Yh�`��L�R=r�.U9�7����_]=W!���1;��-=�E�������s�2���P=yχ��I�<L�<8*=2�	��r���x�=!H��h��9�Cg==r�<E/|�AUu=���<��8<s�<Q⼭i�;�����#�4�n<�3(��̇�=q�@�=(�u�5@;r}s������R=��&�?�$!�<ō�<����7R=��*�I�����<�b|�b4X�i %=�8�ˣ+�Q��;.��:y�˼�ժ<�8�l,=����;-�)���^=��=e�<j1=�ub=��|=!x��	 ��L¼�⡼�L=q�u�����H�8�����i��N���<C��Hq=��H���cc<�����ۻ�	^�a2<I�#��gp��S=4m{��K�<y�P=c`ȼdOy���=	R���P=��<B���I�<�"��P��<��=����7$=�\�<t��<n���%L�K�3��E�n=$㊼������<Ky�<�SX�n�=8W�<e�s�S�{��K=؃
��bJ�U�ӻS
i�G+3���)=X#����{<�)t�Xϼ���<Q	=���;JԼ[Lp=�����$�/�W<'���;ܼ�'=g�[=���*�����</-|��l�= u}�̉�;/�<*=���<M��&)B�� �<k�J��x�<�`��g}�8v;=7��<f�����<�><'�<������|=bq(�q�<�1=F<=�b==�S����<��:�]��g�.I=2�	�<=u��<�^-�'H,=�V=�����g�<,w�=T9 =�w=�j\�V`���¼F�"=]����=�!�;b�<�@Q�@IV�Ȱ���]=�W9��u���Q=�1z�RI?��ӛ�����M����F-����	��;WWX<KL=���lh���+=SxJ���;=}݄<�'T=�|:�f�<���<(�@<=���u�;�:м��;*_�.hI<�Y%=<	�_�؅�<�S'��(|�#���_<�X#�@O��T�t���M=��:@�<?b���X��Yp��y��f�<�oۻ����S�<��.�pDa=K,1=۸����`@��nc�N�<�;C;��*�F�}>Y=,o�n��;�0]=��к����\=��<��@=�\� s��Q<;��<��;�d�[�;�9����<�b��}�\=�-`��,#���U��L x��r�</�=r���<-邼�@w�[���!����y�J&�z4];�T=o�'=��;�8!=���<n"�=X����t���}�e�W��=WL9=�]E���=SgR�R�<Ntd<!�k<�4��#<��J:=;�@=(�F<'J�,����Ṽء$��mN����ab�;iId�B8�<YnU�1����׼/�
=��;�w�z����<�D�<=�;d0��Ep���r�toT�fc=��<�q��@�;�h!�:�X�S�޼���;$M��� ;^=O�x��S�;�����+=�A=}q�<{��_�l�.�N��f�)n�<��@��o���<Sp�<d➼��\�f���y�<=�Ig;y	�5����H=˕���s�h�hA;m�����;�n�=�:�1<%��W�����S;�=Z|�<��=/移�����`H=�8��/=��=L:<��R��[���vs���ϼ)�4��S=�==��#=-*�o�;	��<�?k���k�T�мh�@����<\��<B�=�$���߼��;��2=;;iA��$�Y�_*=6.���T#=�Ę�r�=��*=�)�
q	=�^�H ~=$ʑ<S"��n_�]�9���<�@�S�0�J6;=�%=�ƌ��$G<�논3�5��T{<WBʻ�:�<�d�fj@=Y��:���
l;�;;�v];�-�S�;76W�6"�a�; �;�d>�!m��缗#�=�LZ=?�~���T<���<@��=��<���o��<�	J=����Rk]=.���2���͒1=��=�N�v��;{���`�<;WT<@��<�I{���}i�<"'J=	�!=/�M�^�6���`�d2=�c�/�\=Ǘ�k������*=1���.���+"=�L�<�"��ϢF=�㒼�-�Fw���"���<,�<� �`�Ƽ�C�P��<
�B��3����;U���0;�1M=֫2<�=���:�Ĭ:�cy:,��<�i;9�w=�'��[p��튆�q1�}F�<	Ch�v�==�fK=T�6<9��<z��������9�=���;�B��������`��C�j�1�J=�}��'D�N��{*�<�HƼ�s-<[B�I2=��<E7���;ü� ��Cϼ���������j�;�Z�����0���� <�Ӿ�(��<܇T=W==��)=؞�7�<d=r;�<\�@=�5=z�:=92I�|�2��;?����<e��<��==�-=K�'��<{=s�G=D՜�}r-�}�g=�T=5+=�X�e��;��2�����Z;g=�h������W�漼+��d�?=���m��o���+���ٻ&LӼN,�<[��;��=،�=#g=�r==�𑼯�=��W��m��:�	��0�g��=�;�O�;���5�0<���	칉�'�
ll=P;t=�!�@S��������=p�<��J=�ӡ�!�=�������i�<T��:E���� >=�YH�{�,�N����߼�FƼ}�l=� )=kX	��C���-�0�M=i:V��DG=?R����h=��"����of@���.=6�$���M<S�.=��;���q<~ü�=]�K=^d׼t�=he=7�a=1N��	������#���'�Ɵ�8m=,��<9CC�Wb������C"=m�+=��e�I�����,=\li<��1�d�=[VK=g�n�,�ڻš=���<�ĸ<�|�E�V=��9�z�*=�H=�����D;���m:p�!C=�!�<=3
:��ϻ���<K�<mU=鞄=�Q�f: �m��<)񕻯�%<A�*��[����t�1�<�0=�}�;J�(��N�����"=��m�>�H=އ\=�#O;�<�^`���<}=!S�6�z���켏[������Z�*�x#=���=GM�<�s=	L���oS��#l�y'=Δ}<Wk�<�c!<A��:�O;���X=��̼��=��Z��_5&=,��-f�����5؍�Յw=O��\�\Pp�rT?�6��:�4(����޺��?=E��;!������<e<��@=Mϼ$�+<�nG;Cv=N�;Q�����=�o�<��_=�w�<`��<m�z��t/���<�4�<u'��WK���.=��<��.��Eּ��6K�"[R=�Z:��R���� =<�V�Rh=�_�0���C̼�{2�����Af=�<�7���=SG�k�Z=��(<�B���T=���;b���Ϟ�<!�"�j���g�'j�.k=���Rx=z�>���,��;<վ�<"]5��fr�?�<��<���;�Q;���9Y�ʻ)�3�Xr�<����8���?�<�*�<��Ѽ�r<N|C;�>=W��<њ1<��1�y���Kd=}|"����Gڀ:=�=��<�C꼯����eL��G��],�ܜ��!0����K׾<��o=��
���b<q�B�®!=rZ=:��1"=(�g���>ؼQ7=J{�<]:
��6ݼo�<�sd;�Go=��x�@��;b�|�	��<�&\��S�<�7c�"��=dRr=�c;���=���<�UY��\ݼ��-�K=�r.�3qȼ�c��~����(=�#�l�/�</F������ޜF�|kK=�'=p��<�I�;�%:2˂�-Y�:��r�%Z��z��/>��!=\��������p'�|�0��ٳ��@�"���T��q�g���B�A�]=0T�;��<�����!=�����F�^깼\؀<j�^�S��CT=LƳ<�I=�b���=�V����<�$,=�O.=�v�;VD=�h�<��U;�k�=�#�;���<�2���1����:�"�<hG=�#%�]=k��<#�<�E��=o<e�@:�+�=�gO=T��<�]M���O�%d<`z=G$�:��=Q:���D�b_�<��=L<3���:�[�A�{⻼$Ck�y�<d쌼/3:;�愽~���^�_=�����6�אռ*�=b����":�4����<zYI�U��\|���`�@�l�e�`��K�<b�K=�W�<���<��;##i;�)мWpֻ�D<(�O9�,�����)��u=�>{=U*�=m)�;��<^��X�:,�*<v�=�--=�2]=ň��on�<�VE�ʦ���$���g=_d�<N_:=�a��ԁ=2R�<4hH= C�<)=��"�[�?�����G��(P=N= ]=+}<�&0=$#�<EL�<�!���l�Ac�UwI�W.!�U��<F��<\�<��[�$�a��Y� ����ჼp^���P�R��� �D��o<[v�`�v���;=1}���0N=���:]�T:�K2���Y�9֐�p���!�mw��A��<8<l����<:8	��5?=�@���<5��D~W<�fȼ�0V=��5�rx3=54�<� �<J�>��/<��R=���<��#���l���.����<E#�\��</���̨<�.�<�=<���%��;�jj<K�D=ج�=Qa=��\*�i�;桀���)�+�O<i`G�K��:%��<@%?=!��\0=�t =8�><:1���<��Y=^x�ag�;2P`��I{� �<��P�o\Q<A;>=
�<��!=�c�\:�n�=< )<��N=z�5=��9=�y"=�!��9�"ㄻ��r=z��1���.@=�}�<�}=9�[=��!=XR5=�˗<��_=�bV=��P9�EN��=�q��4=�M��0�����I{<��yv�<e���$n4<�ʅ<�N::_I����2���c;�iG=>�=�����"漊�K<)?1=��#���</ �<�l?=��(��pF=D;C������Y_��c=F]�<֕ =��u��~=�?y����������;�<V��<&�� �;rȐ�֮0��4�P/=|G:���m��4��U=Y�<�PG���<N�6���=��ڼ�5=��޼B=�IQ=]����7�֪��bgx=�:w���޼�og=m�¼���da:��U='�[=�n�<G�	�&�_=m���@���d=߷�(���7��f�:6�����k;�5V��0=���<�X�z<��\(<Ze�<��a<` k=�D.��!;=���<�1=m��<��P<MFN���h=�d�����j�=s��<n�`=l[�榼)vO=�U�g~�<
�:�H�<u�A<�u�<�n�<s��;��Ƽ9���<'=<9U=� �:���<ρȼ�0=_�G�������;��5=ȏ�<�ξ���;�ޔ��~�+/�<�,�<�g�<�W=;=L�<g�8=X��<z�@�UI�p?:�OۻC�?������5=��:<��p=�ڼ��������`���S	���a<���'Q=
�1<WLs;�3�<�c=�Q=�O�Gh;�;<3��<�����&=�[=���<O�B=�B{����]r=��L=�2=�ki<�u�<�zӼ�V��MV<�+��>����?=�s�녂=����{/�<_�<��0���<tnѼ�;�ͼÒI=�=bx=�K;I6<�E�<z�V�[%�惡<^$I��t��F<��!�~�<H�I=��<	B��R�=B<�<ޡ�;3-=X��;f�ʻ`�<V�/=�d<H;�< �<.s=�7E�`�S<˓�<zL�g�8=�F!=�M=�7a��i��<�o�V-�~���T����Ҍ�;�f)��Y����<�=f =�G�<�x<:�ü�[K=�W�;x�
��6��1D<�`0=R����M��̹�aM����`��<�,�V���%G;���kG=`:�,�>�$�8�Elf:>����+�<\�g��]�0=���<ӡ�</�ڨL���<�0�<�Z�<���<2��;{����-E���s��B�<k����=D:��C;+�I��c�;��4��b���V�:�d=�G�pd�<]仛lN=-Wg� L�<$���@���
��f;=¼�Q��(�
��<N�;?��<�1�<]�;=��=�n(�~�<x�Y�\�*�m1c�ߪ5=��N��<�R���<;��v<��Q�ĸ7�3���j;}ȼ���x=��;��S�4��<�C4�<\�N<�=@�=��j
��(r=Q����w�&�:�C=�f�VJQ;�=^� μ��%<<7�Z<o�h;s��������e�� =���q,Ҽ�������\G� S��R7=eA= �<�7�;�B=�C��3A� �U���3��H �2��<b=5�Y=��<%]�<��}��q�G�ƻ~/=���;A9K=��	=av�<�
"�; ��"�;�hn<�'�CX1��'μ/��;&�&=�	=?6�U%r������H���ɼ�<=�{���=$=	=&�b=��Ļgd�<���Q��@l�.�;<c����<�^:0�m��QM��=��[[<��<ý ��	�xA��A=��n<��:I5%��0�<ߕ-�<J<�P��z�� ��<^�g��H<i��Z�0�&�}<xC�7L����:��A=[>λ/$8=�Ȳ<�4�<�M#�=0=��=�.���j"<�'�<g��<n0�;&�<�	l:%�]���� =0}=��!�Ȁ>=,a7��O��6���I��LZB�>E=*U�<����� *�x��<N^r�����g�<@!�;P6=J5���r#<96&=��8��冼\�W=ycD=̤�<@�<�YƼ���'�Ѓq�Ҫ��L�>�S=�{m�;��<?7<8C��uz���"���\<�z�<�y�<)�=>�=8����%D=rq=p@�jS�=�����/L�<lf�x`<�覼y�=��%=G�R=5�=*��<��J�+��c�<6�<'5'��=�� �C��$=Q=�tƼM��<vV=���<��K�,�*�V��9�)=u(b���=]��<�M��w��(B��h�><�>����<�N=m*O�3�G��R�8d�:�5}:��F�W�=���;}b	<����v=�TU��`��3�9>R%��OS;�ި���=�S���H=�Z=K
=o��;� ���7�9�ܻC����3�t�ۼ*p<�b=�h;��f=��&�ٙ�;_�a�'�N�D%�<��;=���=c�Z�b.�<�pz<|��90���Q0K�Y:��=v^=K�B��9=l�~<0�D���V���l�����;�'�#�hxw�<W�28��ļ��1i�-l=ߵ3���;?�t��;�t�򸷻�D���<먝��K�<�1�F\4���n�	�케;�< =�j�/��b��ʶ#�����k;
�6��m�H��;���<ԒX�T�<�x�<SsX�A��bxu�UQ�<�kP�{6<�E���<���<�<$��Y'=A�;s
�:��»�Q�<���<Ә*<�C(����=&8�X�m<n:=����s{�<�x��9F<���j�<�z�;�U=������=�� ���r�켿�'��z=�F�<kqZ�p�`=���<̋�<	���.gg==jA=a�b=c�x=w�;>2�����=5�ڻ��=63U=�H��U=�i�<�@����;�X��b�߫�<v"��=���u=�<����f�83=�@���Z=�y��;{<Yk���Ϙ���}����E'�<�fT< �<�9��Z�3%�Q�;a���j�3�A�<V�����9��I=0�8=�k�"�	�E=c�6=�cU��Du���B��0a=z�Y�z�����w?�;�Ae�)�P=Ĕ��\;�<s>:=�(���:��}��	T�����U���Bl<�K�<��;S�A�H�;i4��u�@��=�L;��<� o=��S={�=F$�I�;Iw\=3���)�<W�m<(�<�&	�]߼�}2=-�¼"Q$=�e<�)=�{/=�A�s�W�:u%=6rv����<�Ҵ�8��Ƅ�<��R;�O=��<
o"=�M'=�zC�a�n���޺-e�ו�<��
=��>=�F�2����>�[5�	��w,����:I��!"=,�=�59=�ͼt�-��=��� <T`����#=S�ϼ�=�����t�=�H='yM=��z�A���l=7��=X2<%4I<C� ���\=N�<=�,I�������<�/���4��E̺j�<���7�2�=A1=�O���
5�t͓��#�<a77=��&��K2����:\��<���<*�(��?K�9��<?A��o��DΠ<Vj���F�OK���D�$)�-	7=��:!���%V=��;�]��Ԧ���<b�+�*�Z�x� =ٹX=�7	=i�Y�+l�c�=@�޺�!=��<@�<	������<�B� j�<��~��fe=~X3���μz��%;T=R>�wl��8.='��=i����ߠ<xVo=�~=z�<�4	<Y����B�'dd<ɤ~���O���W=!N.=��<l�<6�=)�z���U=,N'�ؖ���հ�$D�eB<��������Y�/���	=���:��Ӽu�B��˻�hz���<�}�=*�Z�G�=������B+�U�G=c6�ּeW=���
�;��C��g��X��!&=[./=�r�D�<]^5�+�-=h��!�����<�<�5���#^=V�s=��=�|<3���:L=j�v��޼6=W����V�.�<�N=��_��A7=���<u�=ڠ=�s8���ػa~����<��=F=u�n�V�F�R�G�~�1��<��|�Y���M��e�z<���;�ȼA�=Ӑ��M=�Ӌ<�?�/�6=S#�<�+�<�E=x2��Zo����k9�"����M�Z�S��d�,k�=+AN�|�<��L�+�=V��<��s<�+�<�ټ!�ȼ�1!=��^=�2<����M� ��Y=�Ա<���/3�������ػ�'=�=�����UǼ��<|�=<�#��B��a��<(<%���;�T�@=:�<���<�`^<4M� �Z�:��T%=t�
<%qA��g�l�'���;�oļ�ܡ�F���ND=�Xo��#(=Ȕ$�V����|�1�:4�I�H�6��7<�zM<�<ź"=[�=�g=�h�����<9W>�M�-���˾��5��_�C=�<�![=m�]������o�ڊK�B�B=�N:(<<���`�x=�I��t��<���<uMb�qO=�<1'V=81c��u=�5<��;=;��<2qe����mHR<��[=�v=�0�< m�:P��<�,_���E<���8�=�G�<�Aμ�6S=���1??�R"
�M�ݼ�n==]-q��Z �,���+����R:S��I�'=��t=l�=D�uA�<T�Z=�P�<S� ��繼�0u��N�;�ײ�1컏�!�[j�<<�<W��<�Р�R���}<�'o<�)H=L⋼�¼U���f�<���;��]=�;�C����=�?%�
Ǽ2f>=�h@=�c)<����I^u<<ۗ<.��< �������4�Ӟl=�����P�<j!U��A�;L�-��R/=���<P���4s�
�[<�V��\��;I7`=#�źus'=�￼V��=��˼��#<�)���+=�q�<�i����<=l�>��;ʈ��V'=�Oa�U�l�j=�@fغ$�?��nt����<�J���<ʃ�;qkk���<�V <��wAd�>Q^;)h��%�:#"�:0< =:9>�O(=�_�;����)I�:����^|R;�7�<�k�<��4=O����h��xB�Rq<E���q[=�N��w������f�"[B�i�7�0�=r>=Z��<�\�
�<ڄ��qe�K��;�th=[����p�;Tƺ���bO�M�-<��L�:?};q�N=,�����
�rz��#�^p<Jt�NMT<D�=݌C=􇔼�M =�g�1kZ<��}<�4-<�$*�رY=�=7f=���<P4=��
�I껪�;�*<a��<Fd�<7]_���k�=�K�!p=vD=�y��J(=-耼{����<Mc+��>�<�K=[=̶��"=���<Qa<�b���ͺ�	�;��� �?+���h��N;�ٯ��'��5�/��-���8-=0�:�qe=�]��R���n�\�	�\(�$am�3ļO��<Z=*�=P$мs�2=Q{=�N<4����<qP���<�OI;�ݪ�7�C���R: i}��a�:?����*�<��[=�x��y�ڥ1<�[��K4B��6�<�=Rڼ������ɼ � =����=ȣ���!����z���;�<a���q�V�`"t:�j�<:ڳ��JM��ӵ��:=�4�<��<��1�������f=��E�v�v9/<:j==�B.���K<J�7�Lhw=%8I=9D�=A[�<�h\���7=�a=_�L<t=��C=�4��Z�<l�W��<AX=�`��F��x=��W���R��_��<�7�8t�A\=�� W��/�:����=1�!�;U�t��_H=%�(�r��d=P/&<0m�<io��5<޾�:#&[= �Լ��:;$y;��	��?V�#�c��%H="l���H<��{=W5=�U<%n;=˔`��[I=��=l:�;�_�<U,q=��=��*�ǀ�<��=k�a=��f���&<�1j��Q��Ly�C�q���F������E2��cʼ��=�8��h麃�=�mU;��<�~<��e�p*%= =���<a8<��-=9:���T$��
�=�l.���p��\k<�E�.��7�1��XP<j_��`=s�=]�$�� �[/�+�/=NuU���:��;,q��b =��9I���s�I�O��&Kؼ�/�<i*�<%�Ǽ(`ټ,�%���R=��<��
=+"�j��<�><.J;��(�er�0�@�S�2=q�Q= �ԼUb�b�S���=�� <b�=G��<��K�7�!�܃��
a�yp�%<��up\�G��<GM=z<_�vU����2�5�r��rn�<ugW�N`���E�=���-=� ���w<hl����z�d��X�<v6�<Qu=��=�x=���<�.���.r<�2���!��;� =�D=����D���ᙸ<h�@�T�1��5�	
U��xK=X�����<�ڱ��ɀ�� ��T�J=p�<��<?����!`=�����I�4S	�-�K=mE�<V?%<��Ҽs�,=!,��bQ5�q�<�t;��/ؼ�&G�#Y�����R5=�Y= �=�܅;&O�<�<A�Y����<�(<�R
=���_�(�#aμO#��,��;)�<��2=O������4>$��6��8�<EY�:z�)�r
T��_������J=�+]��ۼU^��<Q��<7^%����<�����G�<wU��kW=��Q�:�j�c�=c�����+=բ!�� ��V+e�#F�<�<x��"���0=��=�܋B��0=uN=��<��=���:y�\u�ۊp�M&v=�4=g�T<��=Hm"��K�<-�:�3!T�>��0�;(R�<Le<�l���ޏ:
�z�wP�<h�L=h�ڸ�rռ��<�J[=ɣ$���k=��*��	��A=qb8=�ͅ���T���'<9@@=�0 =�U=�T=�K=Z?���N�(����;T��<a��īO���B=�	�<|#(�׳�=�*�%&��I=ǧ��o�2=Z�8�x8��x���;�<=���Շ;�Z=�%�x˗�> �<�x�<8k���R�E���w�3G�<u�=!h��2����=mc�;��Ƽ�p��V��ƛ=��DEO=��n=��y�$�@�����F&=(���.�e�>����L�ͼ�t�;J;�<y���m�;&<ΰ-=��6����m$����0�����)Ɇ����;��< tH�Z1ػ�lټ9�&�f�����g�#[,��<��=_o����<j3�+��<n�4=�_����o��r`�����U��<�<�<_�c�yɹ<fH=�.K=^x�;e�߼Ax�<�ԟ<LX��wq=�H=�l�;�u6�0��%@=�"�<P= f<)�k�q(�<�AM=�]�;Qh�􃃼�P�<~m=���; =�I%=ݗp�a�}��ݼ��˼G�h��B�;��>��Wb<���<�B�<;�R�X|U=o�<Y�Z=��O��F�(=��<r/�c1=�>m<��	=˟�;M�K��O!<Ɂ�<�o�<���;#i�[@@<:x0�1f`=����T=�s���=��,��|����7�-��\R=��<�NƼ�7�=���qK�"�J���'���<�]�� i���E��<%=�[ǻ~>�<b}�<�{@;���&�����<Ն&�3l�][�<�xL��`7=��<��0=7H*� i�<��(<�����?ۻ�{/<D�_��sI�22��8�<1<!�W��$�[�P<�c;���<�($=lU<��ʻk\򼊴e=�l���,=�R�<{ɧ<�S=B�\<�T���#s�+�������e��<A�)��=�p�DZb��vY=ྩ<1Ă�D�Q����;=�����<^��cH�</&�<
� ��\�=�;k�i=�m�� K���9��`=��=;!#i���@�e|�<Wat�3���5�.E<�$˼SԼ�޼]Ѻ:3��e�<�v�#z �s�<;m�<<��7>=�j�<�=����%�c=0'�o�2�ȓ<y�q�/�ۼ`Ʊ���$��;a=T�K��S��U =R]=G� <�%�<���h<���&�)�/=
�=���=�O=?xB���X<��Q���}<Av3<Y� �`�=w��<��=����
�&�c�>=4�7�(���1)=\h)���?���Q=:W=vi?<�����|=2;%�b=w�7��& ���+�8ǻH���!
�z@=L��-=�Vb�h��<���<��<Ƅ��1�;! �<'Z=�KҼ~e=�d���W�<� ;���s<]���X��;v�3=�x=�ё���>=d�,<�b]=:�+����9*�R=�W2<u�4���4�,~�<+u=��.<�`y=�����:{�~<s��hk�;�,a= М���`=},.=��R=�_�� ����y�</|�<�9r=�w�<��R<�y��p&��:�<#:��	=<�`Q=��G������>�|='j=N�<(7e�f��;m:0=��=�
1�q��<R�=�J<�GA�y��<q�{��L1;Ċ׻M��<��)=�U;=V��(�<�Jh;KӾ���B=7`ټ&Np�9�k�������ȑa���W�a=� ��p�=z�T�>�2{K=D<��_���&��üvC=?�=ġߺ�"'<uK�.:�9'F�<�/�����<-IC�>�l�f�5;��S��9O=GCH�����}<�?���<Lpl��F�2�g��IY��<=��h� �0�{�C�7�a=,�J�t��<�꼺��!n=���<��ﺾ�j=�
<�����4=W� ��èE=ֵ=Z�ԛ&��6���ͽ�d���м.Co=��$��]μ�R�<}���[�U9\=��*<1ݼ�t�r�'<�hj�yǠ<0��<�D=��v=���M�!��=��ۼ5�Ż�[�>#�<"@ϼ�x=���<�N��e=��A����;J��<sC!=I>��D�3=Xo"�,��<����6��w�#���!��>=5���XQ==9���A�:,λz�����xI���w)��b�*��)%=����W=h!B����;��6�,Y���H<� ��a^=Z�^=�;�)��=؞ڼ�=�=�P+=�a-=�KD���$��X�E���Ӡ�h/=�ƌ<''��S�`=t��;�VW��[=���3G������&�_��~������䂻�0 =ƠG�������.6ڼG� �����@=}��;N��t�	��j�'!�0: =�L9���ü{����3� ���?�x=�}=���<�ٻڴ�<�1��S�*�)U�<�G��h�y���b�n7)<�f�;h�=�u9��>ü�J=��Ѽ���<�.=a������s����ܻ����t|���F����<!w�G<��O=v�ȼY��<�"8��܌<me��
ȻK��1C�;'��<�g="�F�1=�R=���B��<�Ł�"z=M'�����<�\�;/D~<�.�U�;9�=a�����;	�C�� ��B�1�;cL<���[�;k:%=$}�<źo=�+��$�x,k<P�,=�ٍ<��b��D����'\M=��Ӽ�}��%!=������4��D��&Q����e��Ж]����Wd=�tB��Z{=�)=V�=ĻE�Z���)PN���3;Y=�@F=&4x<�	7��͋<6+F��;�<(T�<�桼�c��%�*=�CB=��w�@K��󪻢$c��򃼽ސ��܁�jP��LE�:s=A^�<�<=���<��?�]Ta=��=��|=���<�=����N=������������!���HO�:ެa����v)�<���<���q�<RM=f�����_�}�t�g��3=ާ2=4	�vr��,�+}�<],`=����������y=��<k�';�ި<>v<uX㼮
�<�����#����<��<��K��h���9���l���V�Zj�<�H=5�2�M�	=֗N��i?<o�B�[o���J=-���={a���~��W���#=�T;����ټ,��<�gR=�{λ�:=�-=��e��4L� �`ԉ=I���&�<��;�=�\=������=��L<����|��qb�<A�=l��.��G�}���=�_=� ��LO�J���7R= u=�=�;�$�C%.<�P�<[W�<nT���8���<L�=��9:<�D�]���mH<��;ܳ%�,��Ė2=�1g����uJ=�U�û�<�A��@;;��N-�<����?�<+,%���@�bk��f�28j=��;7 :=��D=��t`�;���<M:B�{j%=�
=�=�ܽ��X=&Ue�͞e���M����������=^�=K*;<;�<�[��;�iz��>���;t<�\=e�m�?�໳t<6oϼV�0����;�X=����Ƌ=f=X��<�y<7�<��o�&��<5=��V��iH<�  <H��-u�9���0^i���f=F�ǼMHV<�=8=�=R�<��=�1��Q����V=f�<мZ�G�<�)=N�����<+�ﻝnF=�K����K��w�<�:�\=�պs�=#1�<S?G=Qe�<� �$x;8
�=u7e<?;#���<��=�rF���;���R��w�;�z�<��ټfL8��U=�ޛ�oP���=L��<�#����m Ǽ�~�<z�;�N��zB^���/����;u"�;�u}=wY��+<#>�<�Q0=��=抓<�(Z:��.=�O=�E]�O �;J������6��&=���#M1�[�;&ME=L��<�[���;�J-=����,�&�D��PG=��1�@#�<B$Q�~?��-�	=�s�=K+�[�/�"�Ҽb��Fo;Bl8=vn�����<���<.5r��n��O�������
�rv�<�=� �<b!�<䃶�<\=YO�<2n-=t�̼�ݿ�8�+;�/(�n�Q=�n�Z>'�~>��v:=��9��m=�B�=�j=Z�R�Ӗ=��t��b���G��'%"�Y�=�����u�<����q�<����;=n��<Q3�<p��;���=5����T��!,�46Q=֙D�&x�<O���^�k^<�4�S�J=��`�e.
��g�<���פ	������XW=���=��s<&dԼ��M�y'�!t�;O�3=�KI�>�1���<y-m8�<��D����r`���VE�M�<lz<;4=%(�<!�u=�4�	T&=aE뻺=�����#=�K�<O��^=g=Z��=�8����RGZ�`�"?���a=n��o����V�kʸ<K��<�I���"<�/0���1=����xC��	;�kX=��[�t<�������SJ�磨�]ꑼ�ؼ�,Oܺ����ާ<Q��<$��;�$��O�s��<��t<]�����?���|<;	ûo�:�W߼
����D<���<��]�I�);cL��+=t"�<�SZ=�^7<D1=�Oe�cS��w"���Lw�7��<�@���=C�;W��b<����s=EǑ�d�<Q<��[��ȱ��ƻ]��<��	�v����W<af\=\�~���ļ�V��ܥ<k�D����<��=��;P��;�	=����2=�aE�����N�
�9��j���<�h�q����d=��û�V�<��绠GK=��;-�X<IAN=񢃽`X]=S<�OּR��:�J=�ȼ-A�<��2��	ϼH�l��/[��gv���O=d[�<���<��= � <b_+=�mr=�>n�E�+�� j���b=����,��ʋ�{^׼U�=�2�<,��N�u��%u�\n� �n=��[<X4���Un=�e�;�I==��J�� �<FD�ڑ�����o�w=t�<��4<.��=��P���=�=�S�J��<
C�;$�|�T�?�U�N=�G<�:ּ�{6�Й�<Z��N_��h��<7���[&�ɴd��/�:ul��ټj��;*!#�M]H=ī@��/=���<|�Լz���Z�`��r=�>3<>O=���گ��	�=�`ؼ=%=%���I!=s=� <�N���w<�Y=
i�;��w;���;���<Cq�=���N�=@�����O�P���J=ڇD=���<��=U��<��j=]�:����<�ZG�G����?���<��<ֿ�����<6|�;9��޻���<+9M=��R��9��v�ҕ�#׍���<��<G�"=�ƒ�Z��; 5�;C�w�2
=!���0��"�J������*ƈ=Q����q7='��o�<v�=e�=�=�l/��"�<p��<���<U�b�@��T�'�7u����#=��m�Qe
=�Q����D~7=������!�@�!����O=���<h�
=�1=m�k�2����*<�9�<q-z=��n=V`&=C+�������,_�G�U<�9�:rB
��ǚ����9�5=�� =#�[;r��<:��.��ێ<��=gy
<��O;T	(=�{\=�1�����<˸X=G9 ���q��W=�1=�=�L[=�`����TzμRs�;�m�<��漱!ļ�D"����<⻍��ͺt�S�d'�Q��< K��ҋ���5�:KJ=�v�<v���$�;<=̕B=M'�G�=��n�j�=;K*=B�={*V=��=��c=�Տ�H��<�{=��W��M/��g��?g�I*I�~(�k���=����%=�@K=&ʥ<[E�<���<;�V�;\�<$�V=��F=�+�5�ƼC��<e�<bB8=� ,���<~������b�=�wO��Lμ`�F�0���Q=�SY�sX���I��9<T�ۏ5=��*���m�YP��L�@���﻾�X<z�==+R>=���2���4�<A�a�`�<�(�<$�<�a,��J����;��#;sU<���y�>�O�<_=�?e�g &��}�;�3�;!?��Q�:=H=�$k�`�ڻv�O=whG;,
<���;S�l:�AV������X�HB=�G��Xx:��5�;���;|8(�ֿѼv�&=J(X=�h.=����;�.=��l��T�\ͪ<2��<���ȃ�qY(=��B=�M.;��H�Gm��j>�KS��.����?<F�5��ho�.��Yi��裼�D;�MU�&� ��S��8s��L4��m�<���	=�/=�����<��Ӽ�A=��J=��9Ć[<wRB=K�h�N0b=��G=A��<W�v=�mH�1��<<N=S�<�2������Y��u>�;A����r<��?��r<�&6=P;�EӼu��I��Q�=��e=d�� =Z��;t����E�<��<�.<i�Q<�)�<�@����I=|����+��G���'��]�|�,=oG�1��i�2=?�I=J7=�(F�h8�湂�y�4UI<�<��	;�&�<�U='�=Xd<���;!!��V���<��=x$^<$��϶9�7�J�T��<���<�Q=FsQ=e�\����<Kb<d����/f���"���m����ơq�G��<��/�����a��<�����=��d���뺛 ;vͻ�_�)�<w�(=��Y={�3=�!üG��������<�l"�?=c�0��=��^<Q�[� +S��	��:�G
_:P>�:"=�Xd�����H|{���{= ��<�� =�v��2����<
��<��J�Y����4��BM��[�<�\4�y��{<�z����e]�<{D5�5��=
��1"Z<Y�B��~=1�޼MM���=Uϻb(�<��D<L�|<�e�<#"=�u=�$�O�<PN=��3=�"���J[=
g[=�V==�<Y�;7㕼zY�{�;d|*=�+���<?��;�> ��*<�T ���G�D�V��;�4=1����:�.��{=p���=Ў;�
�=�e=H��<.�S����Ƽ��+=�L�TwF����:�M~<��h��:-=)[%���"=]m���ݒ<8����g=R�h��!����e$��P=F��<B:2�9>[���=ə�<z�T��nD��pz;��f=�<�ά���f���޼�N�~D�<��+=�4=|�b<=;��*��I���=������<z�<�i?��)�=*E�:_o��D��u��3��<3��<�@m��}ѷT����:¼���;���͙Ϻ�X�<qV�</o=�M��:߻Y�F=7g�<�8=:@A���� ��<2Ȇ<�T�h�z�<ܫ:�LlV=x�U=,�{�*Y��x���K��B-/��fU=:����Ԧ���#����1ڴ<D�*�e���ܙ�jF�<��?<�<�S#��ĩ��j�<�z�<�F�<��.=�(=-<�o�^=�<�<�C=��`=�囼��;��=��<�F)��#�m��@r�\�%�w�m�B�*)|���\���O;R@>�����'�u<B�a����aj�]����[�Q�<�Nw�>�;��<I�R�Լ����N�<���<�R*�XA=#�z�;�:���{�m3=v)t:X+<��12<$W�<�)�u��Ŋ�=7��}�>�Dv��f���8�h��<�ӓ<�+��u����<��\�dS`=<���CD=]NB���Ǽ5��;e9�8��!=a\=\�������C���qo����<̀i=*>9�у꼭��n�/��F�<ԍ�<ˎ���Z�)<;�M�I����H���S�X���=!Լk���3�<��>;��]<1]�9}�`<O8�	�>��H�<���&0=�v�����<���o�C==0���;a���W�<��<0�O;$���/='�=	�*�ʁ`=�i�;�,�06=3���`+<U�<��~�}H��~6���<�#�<R���;���-=�=��꼿�i��̞�3�<�pU=,���o<�G�0{��G ���09=N�B����:��<{*�<�Y�<�R�<ok�<	��<kP=_�c=�4�<��<oO=5=$�;��e>�<Nt<�R�~�5��KN��&$�9��&}o=���<7�$�jlF��'��8�<C'Q=\��<�V�V=�-��8��p=Gg�;��<�e5=�Xg��;�	/�N�a=��m=��==S J<�3=����|_=[�;d�e����<�i[=&U
�Čo�ҴO�_�<���ov<m~��hI��@]�w���/a�<@^=�F=�����u��ȏ<�b<[�V=�@=�;����D9=�����a��Y��]��U���P��=$.�"͘�ʣk=s����(����<�Ah:��B�ť�<f;<��,<>s ���K=��yfP=�9<b>j=�RI��ZE=+�?-�<68�<�6�<��+=Fc�<�MQ=o��<��`�#�۶�<� =Œ�=��d����;0ӫ��x��v?��4jz<�Y!=WP=E��(�U$R=�컻�ɻ4=�ܦ;��L��qԼ�j=�z=�3Q���<{��<<Ѽ9Q��
��������=G���=�e�u$�t��<����7z;3�f=��*��I����NW=���׽k;�
�<�� �Q>;<�fɼ�$=p2�<��n<�і<�+=m��<����8p��8*�}Bͼqgx��18=�����r�<�uZ�S=42="5�<�m4�}j=�c=��^;plL���n=�VO�B��lR�<��=#�|<]0v���t�j�=(r�;�P==�����I�=dм<�z���̸����<(��9ĭ��lMr=�n=l�=�\=��<�t˺�|	�g[<�.���!=��<��<l�<�M��s*;�Nz���V=�Zٻ�A�<�؄=P/�|Y=�s= y�;�eҼ���<	�%�	w�<�C:=\�B�\Ɋ=	T�:\=>�>�0X��=�H��͒;��h�; � �C�N��}~���<t;=ʾ���-=Y�@���s=�
=M$4=�9܋N�8`8����y�:�����f�G�;[V�<�/>=E�
=�����ѼF�M=�e=b?W;��=���}J=�
��WE�Q:�L�<^�<E��sa�<b� =k'��޼ �_<0�=0���v�<=,����;΀�<S�,�����3?�"�;�����B��X
=%�"=��=��}����<��;t��<�\M<mC�!?��7���=�6� ��2L;筺�Ԕͼ����|3�;�G=
�@���;�:� @�;��;(Zs<A��<}-<� ɼy��q�K=R��<��9��u�<�=���;�n)��=&Ԍ<�2��Q}s=��<�J�<�j=���<�)��a+�l{���|�΂a��*�:�r��==_��<],�;���ӯ7=�{'�Ǫ=��H���y�Q�J�1=��C=�00�L�;B@Q��*=͟	;�:��.�eM�<�J��c�D;��p=�)<6><F]y;��;O[V�T�T0�;(ڊ<�~����ͼ���bG���x;�23��5����A2�D�v�>.7=�["<Z)0�LE/��:b���<s�I9�-��N�'��<TU�;Ś�h��ꀼ�� $r=io�b鵼V#|={���s���p}<�%<�Z����o=Qё<��<]9"��`s�b�%;E����%=��<v!A��%=�1=��<����&��<�sS���N=[�W�����V<��@=p�F=�8&=�&<rFQ<���<� g={�=��߼_�=@<�<�By�A};<MI������.=RmX<Sc�<e�~����V=�ӻ���<��	�G=dc��^�<HM��3�"&o���;zI����<D1=	k7=g�׼�O*=�Ƥ���e��;�=��5=�P<�>�<�r<��P=ڐ.����<��=�4��l	;�T�>=�i��6�=��c�� �;Ј�����T<�;r��<�<H��H�:�45=�7��U�9�<����A/=�uV�ĭ�<�]k�8�y<$ml���E��C߼�߼��3<Ǖ=��?����<��&�t������;���;��y=���<|�"=�x�=�U=lf3=d�=�k&<m�7�D�[=�����޳<�
��Ij�Mi=��!��?=�S�;[KB�<��:}=ܧ*;�HZ={�=���!�i�+���ρ��^<�5=/�z;'�<���<!�&�S�1=���<�������[=�<&��;��=����+'b=?�=�ʭ<��Լڱ_=y�m��Y���<�U�<ȷ�X�^��=)=*�P=n;���F�wE�;���;��.�	J�<;�D=�fq=ڶr<�?�%����=\@)���Q���
�? �<�K��O��e�9�"V��̧<���K�q>Ǽ�3�; G��F��T� =��Ӽ���$=�O�����*L^<P��;d�p�q�i; %�<*�1��߃����<��=��N=��
��<����N)=V�¼@9����<�V�{��<�(��Xk��L�4�
�}J<W=$B=��U�)��<���s�;=
�J=���<G-<�]��K<��h<P6��~=��� �c� �u=��i����?����;-ȝ<�#�d����'���97���&V��'$�mo=^�D�w̘<~��ܜ�W���b�D�;B;K<��ň;�;��<�o�;Ke���W=����I�<���=n��<V�:<���=�D�f;�<ڼƻ��:�؅��N=JU���;>J���8�΍��#�w���3<�ͼ[f�<�4=��R�i�=��!���\�g�C<���C�<QR=�R�<H�V�]������B��1�6=��w��.Ҽ��<Ȱ2��	?==c���2��8T=�}�xG�ž��J=��;��=�|�<Ki�&c��q�<*k@��1<��;u�=��ۜ|�w��;
L.=b�����<��);ꐜ��n&=|{�U��<�^=�<=m��<4&�;�_x��N��o�;ueA��� ����-Tp����:��i=.Č�DW���e=
D���<�~A��%�T�=���� g���6�#KO�)���T��񭼊k��M_���#=H<��)=����:�(=�io������K=<�ݼ\�s:���9M�x@����ļ6��ӹ�<i @=F�<+���H=u���x���=�J=���������<�1��,u��o�<볁<��<�Vt=M�Q=�B�<��<E�	=�����р=�_"��pQ�8˔��j�<�.�<�m.��>f��)=Ix��J-;�i=��;R���.M=g��<"�M=������I=��=�6q�>B=��E=��޺񶂼�r�u�����S�/��B��^�\=��<��L����y+�<����pI�j�t��#=vᇼ�7�������ӻ�C;��Y�չ�K��<�����9�i:e��<<g��<eȼ��V<˝0�\�=~=�1��S=<�&�<�����#����<3��;��*�K�*��ͼ��=���ve<݁<=�R�l7��7U�CK����D=֮�˗�lA���P=�2����;��'�q��Ɋ�<$d=;�#�V�����(�U��J�<O�)=�j�=5}��g*���W=�j��6��X<�@T=�'��0����5�ޡ��$�<�[��6����,�7���b=�?e=�u�<��~;����4K�٨���W�!눼a:��r�n;�7�T �J�=bE`==�%t=�%;�9=#b'���9x�=Ψ�����;XQ2���]=D=����P��=4=x���n=iI/=X��;h�E=�?��4�<1=;�;W��=����D�<�r=��a<���<����
��'e�rDa<>X}�-��<P�x���伖�5�Җ5=S��<���<OY�7�=♥�eX�<��e=<�������f<�v�3�j<UA=�U���1�<��X�s�i=a��=9S1=��S<}�U���<�K����`v�<��W=�X���d�e"=ʼ�d<A6���A=e"�N�<P�<��[<�b<�]a�;L��j?���9�<*<<&�&=Ͳ�����*7=�+j=1M0�"�˼�R�M����<�7h��]����'�������;����wG��!=�N��kq=�� ��:Ԣ	=P�?=�-=�W��R="u����<`�0<t"=��<��gg=��<L�]��֌<�ʘ�)��<�;һ9^�:D��<�m
=p5���m� f[<U��O���x�p����6���[<�+��/��+6�������'�C�����<w#���������;U=�){���-���<�﷼��0<��R�CuX���L=�1�!��Dv�q�<x�B��zQ=݅�<$��<�����V�%�c=B�#�BJ8�����]q<-��������8����<'�T�R$=B�s�$��=����4�+��fV�OG�<��Ӽۄ���w0;֎R�+"Ի�o���<��=������-׻�r���<V:�<J�,=�_=J�<�z=+`޼sd=�||<
k=��"=AS=J4�;�pi=��X;Qh;<�Ӽx�1��	=I��LS=sg�;�
t��[=�RR<:�+=�u�<B��;��Ȼ�%ڻ��;�R�<?쟼+�X:�'�<�iӼ7�$��G=}��S�|=��<ؼY=���<@�#����]&<��C�J̤�N�8=OA��]�<��-<�C�<u��<)t=���iX=��ؼ�	|=NV�<�z=$6=@H�]�Y<��3�g��<,|��E�n�"0=t{��̕w��n�.�'=)=�J:=����V�3=t�����w��q7��� =��=,�N=�dZ=�F�;��@�\���T��Z
<�Q���,=*a��	fb=��w=�����U=�7��)�<��g=�=M=Q="=���$/�<�k��М<د8�kyC�t_.��ŗ<�E��S��{<:G=棗�O�=EIؼRi=�)�<�gP��G<<ډV�&��<y�� e>=ty�<Wh����<|�|=>�0;�W���3J<2�?=u�=��༄j�;k��;��;��ڼޯK���A=�Z�<�2U<Z+=h��;|�:�dW���7<,� �y&U��,@<�=��3��P=E�e��,��5��4< }P�
,0=�¼��=/Yɼ�=N�'��
=q�Vl=DCb�Yj�<��J��NZ�4ሻ��@=��[��o�<ҙ\=�X=(��~�	��+<(=�B<�]K��[�h��0��<�=��t<4��<�!*=��{<�q��}��<[��<�!=��z�E<�<*`�� =4�j=�M;<�<V��;f�?=��b����<�U��� =$�H��,1��T�:'��;��;]��<��P�h� �kV�<x�V<��k� >e=�B#��� ���#=>��<�Z��&#��=�桼�!=7�S�̠	�����W�<Anm�`����<�~ϼ(����<�v�?ʵ;�-<��<�� <������`<7i�ŭ=��<������n=�?<��=�%�ds�<�O)�n�B��������<�uK=l�=�m#�U{<g<}r4=�N�,��cQ_�6�<�$vB<��L=8%�/c<w�ǼI�J���x<.&�9��<:����V=W;,�}r|=X�C;&»�'I��n�������<
����C��`<�f�<R�=:��&�M����<m�=ؖμ���<��F=�<漌�g��TѼ��;���;�1 ���km������%=y��<�O�<>�(�=�uڼ{�./�<l=�#�^=�^5=��v�<\o9=f�0�Q=z�4�p�;�N���䒻�x7�MCb�^o�Uܴ���;[+Q�|��!zj�T�x=<'���ɼ� =��=e&�<<=S�Ǽ��ʻ.eI<?}ռW�<�R=�h�U�J �z�<ԋ.��J#���Ȼ�d��<3X��ܰ���,�2!�<�?��>t=�v =i�^�E�v�u"N�����ݼ�����9=���%�m;�LV���'�AY�<�`�;߹'�AFO=~ts9�א<!��ĸ ��}�<��Ҽ�XW�>�8�Ԧ��Ui�v¹�B�<���31�<��;��4�.�Q=�I=,�n=�
=����@��.�<�N��/�;��
<�����<�i=��{=�����5��}�<�4������� �r�"=����͎1=���D�_=�Go=���s~��_Q<��C=Ǔ�<((=�]<M�<}���J�=�:��=�_s���}��
��a��Uw�	��<�N<IM�w��>�X<=��?���;������XW=Fg�<C�_���x=9b�<�Z��I��<�c� ��<���<>:<����U<&=������K=A�b�����=ml�<L�˼D�<y��<���<r(���{E��-���=���{��<�=�O��D(�M��<�����=�\�F�>j�<��o<>j���H���`��"���R�;��J��԰<U�&=�=
n��đ<��g=ǥ�@#l�u5��E=��P=�:�<�@=B'8=+��<�N=e��Kx�<Wq׼�� <-k�{�$<
�J<#��<��8�����1�g��)���ͼZ
.=S��<9>����<�I�;�ד���޼*2J��=�u<[]1=Z�=^�2	�=�= �;]x�9~�<%��:��;ѧ��WV=�5�� ��<��<8�4=B���鼖Wz=��:�Q =�＿�@=��<bm,�=F�\󎼘�����<`�=�&߼��c��'Q��|�<�*=&�=/�Q��I&�sIb<kG����<�<��=�\�<�E��bE=j'���M��t�����9Ñ�<h�4�& >��0�<"D5��M=}�;d�{�^=^���ق/��ٸ�y�A=W��<���"w<T���*4�;�1;=Q�R=�.;��0�,�6&t��9^��=�w�v���C�C�B�q��1t;�1� �E;r��g���x�<.�������%';��<���;|G�<��ּ���ښ}<Ռ7���M=GsD��e=ٕ򼲞M����<�đ�wB�<A漃?>=ޛ+���,��H=��<ZQ=+E�<�E���R��G,=(h=?�Y��1#�w�=��k<��|=.��<����Au=J�q<�P�9��;����	�Q��q�.���=�4�<V`��k7=Dl<+(y��<�]ּd����*���<�䇼U�?��=�YR��=�<C�R;��N= �&�|��<�tb�4T(<l ���7���<`e�=nO,=-,�<�]�@���ϕ9�KY�O`�<��o<�/���k�<�?��_�:�Æv���q��UV=w���F���^��Xj<x�O=�2�nFj=��<6��Ew`=X�=̺_=' +�f���C�2�s����{=a�,=;a)=��;=�@=���<\s��B�<��=O�'�L=��9��1���*#6=�<�<Uk[=��׼�Y6=�Ec�`G�A���$�<�4=�h�<�N=e_;<N�(��-}<ǝ����<~>�<���EI=�t��D�<�Rp<�"���= � �W���)�]��=�͓��y=�q��q�`��L�ZF�:���<�2�x�0=�o(�8F=_ډ��R�<òټ4D��s�=��I=c��<�p<�"d�������G�uo	��M[�_]G<���giJ=�A�;y{"={����뼗
L=�_Ǽ��mՒ<�v���g:�=�_R���Ƽ��
;��=
+;}�H������s�ּK���ji� �=q/=¸���`ֻ����=2Ih�;a�ϮI�~O
���<lq�EgO�66&<-q���D�<���=�#=�cY=�h=�k?��)3<u��<�����e���@����s�ż���;<�&����*d*�~X��l�<�f�<0|߼��=&�oY/��F�<�P1����<x���<q4�;a�r<_#���P=~�8��cO=��=�l�<�+=�A�q O� u����ֻ�{�G�:���;=*e��v:+7'�ꎒ�t�=p����|^=���;�|��xN<LM=�L}<��:�AҞ<���=*P������%ӻf�g��j�<�����=^�<>Q]=Q��H�<n��<MX��T>�.�=T�&��nQ�:=p�^�Otm���>=֯U=Ǳ�<�� =�-ǻ����=�9=G�*=^'B�D�<F�ԻGty�лS=��d���`=8��� _T��u���U�Uȓ<6�Q<�f�!���=Pq
��L=�<f�>=5Dj�����E�9�|=X�M�HbO���[������(�<�cü�N/<�-<J��;a�<})� ���O�=B��<�N�:��=�?=�73�NT8=��+����Z�t����><Z.p�i��̵g=#�<6p���1���o�
B=��<�'M��!=E,�<�E<6�E+�9�8ӼǞ�����(�!�2i�oӕ:��F��,Y<�p��h���'q=��=*m�<�� =����j�X=g���<���<�d=�M���\E�{$�;U�d���G=��k<.D�D<����ⶼfu*�6�<�1/�a0�Jx�`��<�e@=
�H�ޓ!��y�9`���7�n�p<��;����|<�=y�<[��=���<R��l#=�.5�|�C��[�3���#q=�:X���}<x�伙�`=�8i<���=�0� ���b=�����<EƏ�`�=�*=���;&~
=e�����"=�%�;7#*��#�Y�;�Х���Y=���<�D=My=]=�	4�]�$=L�=�V=/����m�pG�<`HF����<_#�l�s9�|�e8���A=�u;Nq���%�0Q`�]�=���;����g�<vTg=E�p����<�MһпZ=����E�����>��6�]Y(=��>��c=i��<��]��@k=�2�U����޼�� =���<��=�@�4��]{�:R�#=�.=�ou��5�<5�<v!7=�Z�KG��ɺ׼���<��=�^|=2�=�?;Ng�v��[s<���<[��V/'��6]=���<�s<M=���<i\��Zw�<�8{��QJ�(eL=��5=��/���<=Lr�<�&=^`�<� ��H;!� =�xQ�5�=�=*��V=!k�b=�)F�
 �ؔ =�=��=z�K=��#��`�R� -�;��V<ݼ��=�Wv=-�@�/D�� �����<��'��F�<p��<� ¼W�0����7L��ۣ
�����u;�:Uy��O�<��=`䳼gY��*M;GfR=�I�����@Z=�����Z=1�B=�#;�P�<�.�:�U=��v=��<s��<�eu=Rt�;��<0M�*�=�0f�x�s�t���=p+��ל���m=e�R=���<�J=��E�!
��{�<԰׼�`!=�š�|��<�8�/�[=I <*�޼���G����<B�L��W�<����\�z=k<�`=2�F=�v�<�=��_=��4=N�Ƽ���< x��E��1��;U�s=^�<>��<,�+4\�~&Y��� ��?��4B�
:������g��Tu�&nѼ�:�b��;��	���=Rp=�d�<�����[ؼ���;cp�~jp�
�=�,i�5:�C�P<"7=��/������\�o�T��$=]�b;!�2���μ��j�Ӝ'<Ha�z��;�a�:�_&=��λ,Z�"e =ܫO�5�0��V0=�l?=Ҧ�҉9����r{a���<INм��,�F[S=���̄l��!�;���<�	^= �<��<�9���.�\��<��Q�e�ȼ�u=|�Q=�mj�Ͻo�Jo<s}��;����v=Gc�<��0<��缎�f�V��#��,�t9B�U�p��r&��~�<<.]<��"="��z� =S%ż���7^%�;o��K�=G��Q�=�%(�r�q=M�F�����[м_G�<��w=�0m<��B=�06=�<�<�^<�w=V�4�tG]<j<�<oƻ�a�x�=� =Ɇ��*�\���><�����s�<1�$�@��<����Q�7==9�H����C<2�L;={=q�<@�j=�QL���f=��<_R=�Kռ҂:=�A<A���|�<��;"���z�<ms��{��;7���6=��<{��<�)=�3�(=<�*� b� ��;�z��R��!�<5΍<n᪼�v��C=�DC<����/<_=/�H=',��=ě9�\�<�X���\�Ȳn=�b�;�im;�2@�ʔ�:C�v=��4�E�z=c�`�������T��3i=(vS=9`:��<d�<���O��<��m=o����K�l�����<&Q����6<H�*=!q�<��<Oؐ<h�sb=7�,�r�9�IV�;�?弊's<���;2y=�K-���\�ކ�<��U��u�,��Ը�<jy�H�U�z��<1�<j�<�j�;��.��w=��<$^�����m�"��ǒ<�h�<�C=��=H�d9P!�;[�E��9R�F@d<��ʺ��<h�D='��<�13�d�:�H�Q=�"<=�{=Q��b��74=:�л��ϼ�Yպ���[0=���:B�<�f%<!@�6�l=�큼o'����;N��'ڼ��s�{�=|��<�Э<�v�;���<6���o�-��.=v�b:�u�_ �;>W<=J^<�4<�;J�BV���<����f/= ��:YD<�����0��R����<��J���X�R�<�#�h��0h��<W�"�[�<� �B=<�?v=��߼���<tuJ�
b*=�G���� )?=s3A=W�x��v=�o<%���.�;��;��q�&��e���W,=$��r�W=9����f<�{�����H=-zR=.GE�>q���R�f���������"�D���8=j��;=�s�bJf���L����<-�=��;4�	�0��Pb�
��<<$=�O^= ���&e}��X3=#�n<_��<�C��.��4Y<0�`d�<\{Y<��8<�H_���f�=�ϼ�3G��^i�K�c�P<?=��n=���:�dr�g)�63p��s��W�*<�{N�
����H=�1��a9<&�	�+n��T5=��<0��YG:���M(��) �t�$q�<�\d:��X=�A�<��]�%��;�'Լ`�&��'=ߧ�<��`=4��<�&�<ߓ�<]Hk=�̼K�Y=)%�kQ.�?n�P�=(�����!<�\<!��<�V=Jv�<ԭ*�z��<Xԅ<�+L��M=�^�<�b���;+�����ݩ�z�F��[i<)��<�0<�����;p3�|�l=_Y�;16";����O�Z����<��=߻���]<;�X=O�<��<��}=��&=)�߼�z�8��	�P�+3�}8<�f�5�f��Bͼ�{R;e&0�ɦ！�<�~{=�I��}O�{�q<P��;.�4=���<U��<��n=��<��C;�O�u�U���<��ʹ�O��q�<h䣻��=��6�E�<3�I:bb�;Jf�<���%����Ɗ=�7ռ�9<�+ =��ټ�=d=,���=���;�(�<��9���B=�L�;W���`%<T��:0��>И��E=&s���K��0�/:0[;�T�=���F=];	��0]��^=zT2=p5�<E�������=3���*��r�<_ �J<7�:�w�<�w�<W,=����GUC��LQ��4=w#ļ���}R���9=V�#�<V�T#׼2�s=�U���EF�;=I=d}��$�l=@!��ZE=�<���ųP=6���)=��E=����Cѣ����������v�T�8�ͼ�O=��;q���7� ��=���<���ePA����<C���bK8Y	��p�;�WH=} �0�ҼP���������;$f�ǩ[<����Y������x<0��X2=��V<K{��}��Lu.=b�����GY�cDp��t��������|M�
o;�fs��i/�^=l�=	 �<{=K	�<B~ �=��M<��d�=�W�<��<d�M�U#w<Rb=2�g=hU<�y䊼�g<���μ����L��7�l<1�P����<�7_<�1�<��<�<7"��%3=L)�<l �� ��-�^�Ll=� ͼ�s[��E����I�=
���?9�i4�;;ɼ���<� ;YC��%=V<�<���<�:_���>=}0=G�F=�� �u/x=zV6����<sr�<d�<94(<b�<F��;9�=����1�<&ɛ<��'����<��;Gr�<�s#��*��༌=�x˻�q;;�.�< �d�!{�F��0L;1a�Λ�<5���Mv=i�(=Q��<�,c<QNb=��,=l&L=�02=2+�>,�����<Y=6G<;�����1Z���M=��=�]R�Z _�h��M��� ��K=��;�x)��;U=���SBu;z����LI<�Pv<ZH=`�,='Z<����2�;��<(D��]���\�<�O�u�-�]�E�;��;{� �s�<qXp�p>&��֨;��=�gp;��Y=u㳺}�P;'�N�=���@%����<�)&;kfh���<Į��]%=LF=�ȼ�S=�h��]�@���o<���;��}�B�D� ��|\�ց�<�����/ڼ?&�{�q<^i���f��]麊0l��4;GXM</�;o��]��%�;�3�AJo=��h<�T��+�?�	��Q�;�P��},.�y�N���;��M�-�< K=.�G��|+=DFɼF��C������b�<�X��D3�	e��o����P������;�����<;b9	=�'!=�g+�N�5=~:*�b�W��l:=��Լp�-�t)L��V=�ռ��<�]=��ݻ'�8=��ʼ3�\=���V)J���K=s�=To���ߚ��{ϻ��;}2�<�p=�맻k~+�}���{��V5$�?
!=���<p�M=1����,�2>����<�03�>��<��S�t���&5�5vr��K`�t ��˔�����<ӓ=G���:�G��:��K=F<;=��;Z�L��񅹰�;�m�<��&���4���Ӽ1�j1���N8=��<���;	x<s4[=G�;N�!=�59�׮}�T�����<����()���ֻ��Gm=�h?�n?�<e<�I=�-=�w�W�;5�=��;p4��f;c�%���s=tsʼ�\�V�W;�=�8��4�<nh����p��~9����1=�D�<8>]=Fu�H�z=fs���p=�'�<{	E�	7�;"=:=��=~�{�2>t;*h�<���<��:s����ּ�S�<�w,���2�e<��;��o��D�_��k������7E=�~�;6�^�PW�525�.��m4�<�q=���<h�q<Z�w����<�DL�Y�T�m�1=������D/��׫<��(�_�:� �/�������`]�&#y=J���;Ԗ���]<��8=�@=��$<��=�ZS���==BR= ����0��gp�2�O���ռ��5����X=7�=Cm�z�=��a=H�!�ot���C<��^�6O�:M�%=��ۼ[�X�&Q�"�-;�=G=�޼C�s<��U����i����67=f=\�:�T~=�G���?�<69=�����E��cL��&��d6�ݣ|��<K��2 �=�Ź�r��-\;w�p<� 8�G=)�==�m=9��m���x��=��!=�=�6м}I漫e����<3Et<<?Q=G��J`�<U" �J!�<:��f����<.<��g��=��M=��I=�4=3�Ƽ��D=��(�n�H=�k�<��<�̸<�� =�p)�#�w�Ngۼ���R�?�8<+<�:=ب�<��<��=**=U�<�v�sWe=G�\=�h=�Yg���ܼ����B�Ѽ>�Q�ю/��9E=R� =�t~<��=����l���e<�؋:����O<�T=�ZW��ϥ��9,=K��^�G=��.��#M<A�:;t.r=$��;I��<^����!D="��<'�5��(=u`_�`� ����<˫޼,P'=z\�q3��pK����<�N�GS�(���bi��-����9���.=\�Q��{���X�1KO<2T�<�"=�&A���<�H¼�s����T=�����)��;()�;"f ���=��ݎ}�60�<�<⺿< �\=.#;���D=�O��"q=����cQ.�)�~�`�<+�=�4=���b9��|�L;ɻG��/������˭��R�=Yǻ?b��w<e뼮v�:�<<��ؼ-d�<�^=H�A;�:�VO�-ʼӻ�<�]�uL<K�?=~��<Tϋ<~#���#=���;��#�C��<t��=,�<�f�a"4={�a=�9T=��r���2=R��;A�!=��=�{��N=�:(��m��C�W5,��+)�@0!=vlr�4`�q�;(�F=�9�����<E�=�0=�|�t�D�j�m�ۼ���h��Q<�[�3=�?a<8!=<j�L�j:�v=��#��и�<h�P=���l�7��8= ��*�<A���@�=�KM<�*y����jH<n����=��=!s�<���ZF���:�YL�*9H=V	=��y�A�ߺN�Y='!��e"��(ȼ���5�<��;�(;��"=i�1��)L=����4L<�-�<�,?=�P.�Ζ�<�_�<9�<W�3�с =F�<��O;��������:<<ͼ-�-�����W�<�fI�ʬ�-I$��Y��[Ǽ��
<�i=�9��h|a;n(D=�G�V	7����;�5��Ā<<�@��Ӽ'�5��=vg�;T��<{��<M��;�/#=Ş=I�K�,�~���<�=�;�	�<v=3�<�,=M�ǹY;>�ݝ7�G���U=U.�=p4=I��U�O�}&�<o�'�=AO��\���\�<֢z��<�#db�zDG���B;���{?�<ܵ =�����<��0�
/�uyf<я���k;.�=_�W<9*�G�C=zmѼa�
<]Rm��<�E��r=����5]<[�w�M��\<��p=դ<����!꼻UQ���*���V<�5=\�x���ڻt� =���<ڹ�<��A<�v�J�|<�^1��E�T�v��pT��)=l�g=��c=QL=��X�=���<�0$�~@D=!򪼝	�<.L<�7�<�f<�D���-=K`F�y�R<BD��ROT=V�r=(�)����"�=#��m$0�@A���^��&i�;�Z����T���H=��l������<���<�P^�l����e�:@<�r�;J�I=�>�<�<zB9��f��-��<�^�<��]=�	�<��<��<Q�_<���<���l]���:=;��-E8"o众en��H��{����6�㱻�G*$=qrO�h?��&R����:�:i��^�ų�������T�0<��_;�L;�g�<�ok:�.�<7[�S�8=��+��.&��܁=8���e�<w��<�!����<�u9�([=٠Ļ��<Z�e=-@=`%�烻vB�<V�L��2�<�iN=�����������!�x�=X�8=��<(�b���8�'<L����3=p}�;]�-��zf=�[=n�
=�*=��p<o��fc�<�M=G͜���μm�/=4c=ϫk�,>�[���%'��.��]�<Э=�`6<���?W<�*A�<�%<���}�f��99��%�<{��<���=$P�>�N����:���A;����<r�9=w�ۼ㮼f����q���t�'�P�-���;=��f�4@������E��t�Xf=;J=IH���n��s�<ңU=��`=tw=L���q�;/�=Ba)=�]e�)����K<𛽘��<r�c��K��9�ӌ)=EEA=�m���;��[��+��������<l�_<B�K<ݷ9=��;1�(�	4 ={^���_5:� L�'Ɣ���<<]V�<�� =D�Լ��=�q=�� =��<o2�;n��s�V��k��6u =��j����S[�</�Z��Q�l=PW�<V^���;��=fF����;x�3=�8 ��yϼQL_�>x����<!�����a�Y<�Zh�ǜ�<~�-���~�[x(=O�
����<�1�)y=�޼wGu=?��<'Yw��n=�k�<���3���L*��;|:���-,�5��|���$�>w�<��<0����.���z��r��:h�D�S����i�<l�:�cP����<k� ��Ø����<u�-����@"�Sst���h=0q�&s�<]�ؼ����ܼ���;V=��x��������(=T��q���.��	�V��:t�=Ǳ�;�=]�K!���j=푊=
i�⼮<�{H;��7=�$��
��ϼ򎠺X����c=F�</�׼�:=<�W�<�X�<\�Ƽƅl;��<+Y�1�G��:�<�2��������y=�SX�,�=XO��ǃ���$�\"�<J���U=H6=	�R<���֧f�ԛ*=#�=lC�<H�V��{9��G.�=h=�N�A��=�C=^}G<+��<=Lǐ<L�d=�wL�K�=k:���b� A�sn�˘x���<�$=u#���o�����;�J=ӣ:��,=M��= ���<�Ħ��7�;=���=�?���M����<w\��6[�����aS�;���;��uҿ����.����@��Q��5j=pؼ��]�.\=P d=�x�;�I���=$@����<��&=�I|��^��%Ӹ]-�;�#i��YT<cv�����mWؼ]�;�37<fO�<�P��_ڼ�sh;cX� ������F<����_�t��=]=��ټ����T�<�d=�p?:�~<����"�6=T-\=�8�<�& ��?"��!�<�_�<���;�C=��Ļ_*�	�<=�9#���<��{=ϢH=X��*�w=�I���뼔��P.<c��<$�`=L�#�d`=E�&=��
�Q�:=:�L=��<���<R�5���8>B��틽�ܼX��;�� �]�Z=����=���Q���V��:���E�<�17<^'�<���P<��9�->-����n��:�Hq<oS�����%�t&R�i{���DټVR�<�t�<�&A;���2#=b���Y�༮�� �ȼ��8<}�{�z���4=��Ҽ� R�,: =���=E�i<�@-=��F��@=����X�j� N�<�EH<�,<�W=*�=6�x=�`���=���;ȇ=��;�U$�ٝE���=*�0<�sp��?<��7��e���=t��.~=r �G|�<��=��z;��;��Y<��i�ӻl��kN�����>������: ��;\�E<�;���*�ӭO���<=9M=<�=����4���%�6���e��<\�q<���C�|<;�=��5�ڢ5<4-�<��=ԣ���=C��:�#+�o*=�GB=!
���4�<�z��n]�ZO����'��uJ�~�5=�X=u�J������8Q=�c
�ox0=���_�;*��,ݼ�.�;�>󼮍�<�`�i��=n����~����#8/v�^�=��E��8�����<�|;�	��8{<e+�<-S<���=���<�c=-�����<.T=c}I=����em=�+<��#=@�X<���=DS�<Yz�<��-���6=]��/lg��叽�^={��w���E.�;�@0=�sq���'�k#'�b�y=�y����n<��y=�FN�P�8=m�<=��<�_=ػ�4 �Ξ���T=��G=��;�38="97=�9��6DZ<،c���<��=�Dn=Cc�<���;������3=��X�	�݂8�C����<�M><����dY�Xo�\�������Vg=( =:�˼(����2��{u��3
��<�6=!M<*�<��:��	<���&4�<<$=�{��4�o���<�J��J�J�e���5=H��xZ�W�w�{7��-=(ͼ�KӼ�da����.R�<6��M�=�՜<1�=�&�2��͒"=Q�;w;�R�<���<ϸ�<�).�^�I=��a�D��!v$=�S���pN�䟴<�">��QD������d�d��:���[�ܼL&_����<�i�<�B�¯����L=Y�ٺ;e�q;��¿�<v%м6�<�2�<�B�:�_κaQ\�M�:��R=懝<�0껮��a�\���;�C��{�g�=��;8x�RG=���<=��<l�n�_b�<|4�:ٞ
<�Y=g�9={=��=�n��;B�5��g��2O�y4�<������\ۊ��%�<�tL���<�\�2=y�=\��=,պ<!�<��w�J���bR=V�_<�(�����,v7=�|��JgA���&<AE=�Ʀ;����U(�� =�Tn���ؼHy��WH���(=�td��8*<�<s`J=��=��M<�>B=?�Q���P��� ���F�ӱ���'\���X���<ș=���A�G=�ȼ��t=M漿"Q��⤼6���Q���K���;����{��^��j1:=�Yw�)#L�d�ü�!~�O�W���(=�E�<�3�<�IE����;{��<aO���uo�|w�<��<��g=ȅ�<�1�<E@(��m��(��B�M=S�/==�;F�X���<N[8<),<��%���6V}<�����;c=J<&U�Y3���ȼ���L�I=��h=��D��9|��X�:�k�9J*�ӱ�<0t����r#�]{�;A�B���1=�l�����Ri��xs�<��I�g�=m�׼,���|�<�U;
����R=��5=��ܻ%�`=���͍���c�&� =��C�i+=���Gf.��/A=���g����B�<�Z��m#�<�
λdvh<��m��3=1}����$�"<B���4=���<�o=v�'=E �����<Ţd�^f[�a�=ϰX���<s�<��f=���ߡ�<+�T?=׻:=dt��-K!��c<�v�븈=Z�B=�m�a8�VC�=��Z=��Ӽ� .=�5�l����+=�,�bJ��̂0;I5=N���vA_=��8����<{�B9��C(���y=��H=��=wu~�I?p����;f]���!�(<HF=;��<��!;S����$=񗩼�KN=��Y=�g�<�-[=��<%�Q=���:��W=���7��<k[q=�E��S���3=m�w�ӝ����n�����=e�C=�y�<�hh��+޼�\=3=d�V=�j)=�V����{�<����<�(�;I��
�<1,�;� �;� �X�=��9=�[V=- %<g'�<�m\=�!=��ƻ�)=X�@���o<j6�X=�����I�Ʌf�`�[��<v�a�q=J.=E�e�"��T��&7�����< �����Gp��"'��85�;�W�"�=�n���Y�}���<<=J]�<�@#=V��ze��Q������I���!� �=Z�a��/B=n=�a�nk�<��,=ݖ<A�D=T�0=L�;=F=1TY�q�4=_�d�Fv��^;.D=�W=$9m���0=[����=�7���<)y���;ɓ;5���)r�=37>=f�3=���*׼}�=���;¼�ͽ=�z�_Ȣ<B͠<8�غ�x��5�<��"�>�-=��<�)=ѭ�<~���V-H=�d����<�0��W4=��<tK��H�(<�υ=�XJ�v0��Y<&�:='���>=�5�<%�2����V)��;�����<���=@��:N��<�U=H1
=vU�P;=t�	=�=5jb����U,�+��:�w���m'<\�X=Jw�<OB���$�����2��)=�Nj;V��M�<�黻p�K<Y�]�s�N=�N��FU:Z���~���$��^�<#/�ˋ=Fŭ��$o=�F���&z=�_,� �D=j\Y���=n7�<�໼�{�i�H=��/<F�����:a�<��;gU��)��W�<���<��g�����ώ���,=��"<�_H�9�t��;�=<�@�=��R=��ټ�$�v�4=��=;B�%��;/W ��=��ݼ�����;�A�<�tA:ב�;��1=}�=�<���P��Y�<=�ɑ�_�q<�꼌�s�k�9�ࠪ<X�O�y���ؼ�އ�+*����ĄN�^l�;n_=�V=�����I�J\�<�y7�(��<��S�qa��7�<h	;'׼(��;����c�N��*�@m=���<�a�<Tj:=�.Z=���;j�D=��u=�d�"�x��n =�Ua��Y�;�
��f?����:IY.<�iż�v{<�[h=�p �{�J��e�=�-r�eу��1=��Z=�vҼ��|��<t�X�I�k�<)(��md�gtq=��=�d=)X���ܻ�<<G
f=��8p����f=�'����7�}�.�5���������=��ݠ���O�<6I=�,�<7 �<�'='�<�H�㟆�K�!=gio<�.�<L�>��=e�=b��<��<$v+=LU�<Χ���8<��=@hn�����T=3*�;J"���<c�,=�\~��[�=���(c���=����H�ļ��h=��j��;��!=���<~%�<	o�<ƺ=a���2 =y���C��n0a6�м��o8���E=�(��-v�<���8���D��Ҭ>=X�?��ƻ^.{=�;_��=,8=�!�<dri����<]��ǣ	='?�=K9����w=�n,�7�z=��4=̹
;TU
�|���*��u����6�l0%��"�A�f�Pf�ԏo<�p�<w㱻���K=�ɳ���T<��X�I�y=a����	�f�=�Z�<�^��s+���;�ʸ<0�Z��3�<nz�I��]T_<Y;�;�7,=2�\��o?���̺�;SK<����j�����f5�TG�>m�=+X׺��m� ��<� V=��A=�|��Ue=bV�r�E=�䨼@Я8�&߻��2=��J=z�����V=Y�U���a=R~�<�<n\=�V����?��<�o<��3<̩�<���<��^�} =r]=�� =v�g=�=��=����F�<,��Zg=�c����;�,����|�#��<'C=�C�<�4���>=���< p��V9�8�-�٥��W*�Fb�DC����>m�A{C=���<�.&;"
C�&�����&��'�<p�H=���<x�A=)W3<���r�=b7�=�u1=�&��:I�j=�� =�*�z}���<��";�J�<]B/=��=�ގ<�j��=�0O���	�B��6cE�7�j�a��<q���Hm�;�\<2�<��6=�>���7�~��<~ܼ�y;��0����r������Ԋ���j����s�<eX{<��1<���)���O=%��;�:A<����.=���\JP;U�(�6Y����޼Z�_�ꢚ���X=�%K<��<C)�6�P<V�л�#7=~׺�)Q=x���#�fռ0��������� 5��=�}W�)e<�b��7� <<�<��4g=�������@�:D�����$1=�Sx�I�v<{�6=��m�CѼ��<�}�<��=��]=BiV�4���&��^\���Ud</�4���|��\������Դ��M��bM���<[� =�,=�7S��u=�[)=���YG=���<�6˼��e�=�f�dMK<�ͼ>�;��A�?@�<��C=h�׻��<���<Q�	��<6Ɠ�)�D�"�-���4=?�6����<��ʼ�)^<��=��ͼ�k<��ͼX�<2*=J�T�JN���*��9�(�����[��<ëK�y���H=&+p�Q�H�n�����q��3�<��S�~{�<x�^��#7<M�m= Pݼ��TU���ټ*xQ�/��_��R�U<�㍼�EL=G��:��
���=<��+=NӅ<3��<L�l=ڃ=6k������N@���<��;���\�=nZ`�ޕ�=ޙ}�t�?���=9�e =y`�;��<��=T&�<I-n=��<g�ʻk}��r�󼖞8�I9=%�=��+=�G<����3�"$���<{g<�8�z����h�J=k������<[F^<��c��<��3��=��J����IH=n��=���y�":}���,<L@�=L��HA�<� )<haz=��=_� ��!�#2��}m�u	�<xT�;|Qf��'�=���<�
X<`9�=M.(���#<���E�b���x��*2=�<��L��;���:��<=eHλ��
�]�<�M�<R��;�,C=�U��WcA�T9�R�=4�;=���<�:=�Z�|=��)=�KF�J��=@82<W=��<���>q��x`-���{��?��sH�+,Y=�R�<o��b��ϟ��IF��s�<�W�+���:^ZQ=K���M�F=�#k<�g�=�=�m�=-���	y�<�7	�v���9����;���Cj�<�= ��8/;�<�x�;���Y<s�Z����U="R��e�8���</�ؼ�Wż�bA��=@��x�.�7���o���9=��x=Z�<�_v��E�G=o��t3<m�#�Z� �����Hb=�vb�����8<"=��	�^���C�"=5wZ<;i:=8��z\=%�b=�:<�q_9=F�<�B;�����;��$�*��W����޼çw<���<��B�~��f=��==�Y1=��;��`<�r8����J�<�m(�zJ��m�<��ڼ��<;��(�(�6:�"�rxX����<H�6�Zw<!��<����9ס<Nʻr�*��V�!n�<
H}�99лl̓�Yڼ�m�;�9��=��z<XD��v�����0�=d/�$x�<_���VbB��c�%`J:���<���;�b>=�Ӽ�Up=`�A�Ẏ��-�=Y�;�7,��H��A�=R�<i��<��d�L�?ŀ:R������� e<C"ü(#(�uW';[��`B���/ ټ��l;�X�<@O2��>(==u�;J�����b=�>=�哼��<�r:̳>��ę<d���Pݼ�ە�R��D2�8h9�<�:�xM=.f��du�_	E���<�35=�
<�%_�
��<aW=�4�׮��U�y����}� 9=(|j��ָ����>_�<��"��=8y<!�u<�P`=Ś/�5�J=�!U��n6�k#��	�M��z�b=Җh=��I=9"~������6:=k.x=��$�d �q���6�	=~��`K�=C
�&������Y�1�=��L=ͷ<$#⼈h��ڱ�<'�%�=�8��m�5���(ټM	�._���A��c�=q_�;#=���臼 ����\,;�͑=\�=t�=z� =3�K�d�M���Y�T�\����<yp�<�e��*��@A�<�<��ʼ7������<�2��]����k�+�@@��B"g�%�c��g=���R�<��7<2�+��:��$xs<| @���似
k=D`�<�:��N�<�Q=rޙ:=�9�n�L�P��<��׹��=T��<��<$�v�9I=��u�Iu���I.<��:=��E<d-<���<���H���)=��f��e���]�wۻ�\=�K�<��<3-��ˡ�<p���˴�<G�T<�q%���J=G'h�E�����Baļ���<K�=�R)<��;);�<�]��X�=�=��e����<�Q�<˞+=iw=�q=���=��<Ʌ4�呥���6���2�dA=�[2�ʎB=���m�0�^Ak=�Ĉ<|�_<Vc=��c�	����^C��}=}�<�@�
� �R=H�R<���<%~T<?���CS:�@�g(�<��A��<J<�w<�m�L߭��T�<��k}º~�i<X�<)#�;�QW=��L���<i�	=h<P�@��6��5��/:��S:�J���c���伷S�q��=q����8=N����!�>����m��w=���m���d=<���r���&=Yg!=���=�}:'�ڌ��H����˼y_�;���<k�3=8"���@�<\o3=�!�?q9=�	=�A=��=aOw�I�j�d
�@\=�~v���g���Ż,�V;�����q=k�<���]�`�;E=��/<W�$�� ==��=LV����pK=�8>�Z�O�RTD;5%�;��5;�h <ST=
�=�;=Nl=e�<���و<�6Ҽ��$<�f{<t��<\�c=�D�<�<!��;%c�}�.=|o=�u����I,4=H�;��)=�+;�� �<��<��`�"�/�Ż�:���=ZC^=z�K;�ʼ��^����6���s�q�=��*=�������=��{�6;���<mb<We��
����;����C=T��'=�;s��;��#���=�ŏ�Ae���1:��|����<���B+X�I�,=4�]F���»�ע�\W�<�=�"��S;��R<�o)�!
^<�Q�+S��pu�}Ω�5���5�<J%ϼ�B�;�c=�\�<%]N=s)�<�5�2�@<X8B�rb=���;ƚ��/=E�f=�=ʂR��94�P0d���< �e=��=��,�:DD�U�^=�H�<d�f�GE���=�\X<�@&���)����� 3�0�^<�,�<AJD���<�F�!yB<��<��7����_I����9�=?��<�1��]B��޼�$T�zN�;[s�;\��iQ=�=Bf>��G��Ȇ��;ؼ�M�>��;V���h3�<~C8<*v`;z�<Vܛ���~����;�S������Ӽ�u=ʩD<Q�<;2;_�Ӽ���fS<جK<Ѧ�<0�Ӻ����mǼζ0<���;���;Y�L��m߻����2�.�r���=�����Ng8=�Q`��:������=��(��=��w8�bPq<�<�=�}���v9�O=��<P�e\;��"=;�<�x2=@f�����<�ϸ��W=7�<��0���<�9;��`���R=*�-:U���KO�<V��<q,��a|S��3=����w<L�l��gG=u:��D��(�;��C<� �q0�<b�r=��{<���<��<�b�_�T�1p��e!=~%�CR�<Ĵ�ځ;=<�s��m0�uv��,=?Jk=�iN�hȺ�^�<�ڌ<��+����=�e�%�Z=X׀��r<�;W��|�<������ۯ��hp<x~��W�<��z�UY�;��`�=�����3�#M=o��<��w,><W�=2����I~<F �ԝ�<�P=��м���/n�;ꐴ<�&�>]�<H���`�<��-=s����
���-*F��=NEE�����yw?=L�&�]��<�1��ͳ<�%����պ+�+<�φ���M���1=�=��iI�<�<g��;O��P7
����;1�$��'�d�P�S��S��uű;���;t#=2��w�/��<m��~�P=�%=�4���;��<U�S�*�H�9��<&�<ë	���=5h=Y>���.�Aas�H��;�Y��<�d���
2=%��<B��<�zռ��='7�<$�V���3=w9=*��<�(@==�k���3�b�f��h<=K:���L�k�)�-��)
=��`��iQ��G�8=�ͼ?2зo�<@0=�[ �z�����u਼c
����ZV ���R=p�<�W=��P=�{�E$�1��߮N='�6=��H=�2�3�e=mb�<m!d=̦h����=�[�M�<�E=>��<��мܐ	=��<��<�3=c*;=�ou��Y==�A����="�N=xί��c<��=/ۼW��`0���6M������d���;2�����|���#=��=�)<cp��w�ʼh����O=BP=�_<�Z�<�oV�Y�<�>r=�16���/< �I�hY=�#��w<���B��^=J�*�˷���ػ��"=b~e=c�?�օ������d;õ6<�J�<yk=�=dJ�<j'M<�ja=�8�{K<B����'/��.<��<��[��R�����`]��s)=��I=�6�;������B=�!=��;=�f���`<IZV=L�O�?�&5�=)żps.=��W;н�<����5��a�pp�<�x<�	��F¼�������<u��A�]��<��<n��_�F�u�=�&=��(�Ys:��O=��m^� �4��3���-��LR����<S�<��=���<]�f;~��<Q�l���a<��9<��<�E���9��H=���=X ����
m=���<�F=�.=�	�8�_�U�g;�i=% =F���:]�]���h=�o�<p���|C;^� ��1/��.<^��<	U�<���U$=.�<�,1=q����V��߻��LR=��)�yZh���`=:�ּ��<e�)��L�;Ԁ=c��<*Y@=8�:j�m�6I=�r7=�"o�U[<r,���$��D�<�ֽ����;e��<�7?=�T�<U���4�4P;=(а< ��j�f=��Y�]_�(���3��O0�_,~<�E輾��Jk����W���+�[�o�=���?��<"�=σ=��R=X��	�%�2�b=��A�Zx(<�>=��b�����#;Q�</�,=���#=u��/�=ǆ/�l�ּ�Q,=�?�<\s0�o/�<��J��Ӡ�WS�*PI��Q-�ݨ�<T��<��v=�y�<䴻���>h������9�)'(=�n�\�=M�B�$Ge=��-�a�2����+��pw=O�W=!����U���<0:����������A��<�#�<�qi<���;��Ӽ������=Ϡ�1�2�ˮ��{�;s��<���:d�T��6V��&=x��<_�S=KX�<�4���*<oPn<�ĉ<��N<<�+�8B�<5�<d��=�����o=�+)���ɼf�Q�Qͻ��6<�]�A<��U=A�$�c�H=b<2���@�Q��g�<�JE<�W�dz��[d=��)=*q=���������_�ry=���<>24=�A���r�Ww<�=ب2�>Yj<h�f<��E�͑�=��@��m$�5@�;�G��:�º�=�=l��;��;S�3)�<�i�M.��{�<�VD=*j�<�׼����T������$=�
#�k�h=d�\�5j��NE<��<>�$���1<�D��tLF���<u�3�J�\=�=k��t�q�:l�=�=���}�<��m=�K!=lS�F�<�z�<��J<��	=���<*Z˻�%O=�y@���J�]格�,��(X=�Z(<�	=�(��IX��D�<j�߼�O��F=�|� �Ӽ1�=D{�70;&~�������$=�i$=tf�$<+��<k�`��!�a!Z�/��<]	���=�s�@��y!���NŶ�4�7=���<�n�:u�=�}Ѽ��+=��
�M�*='=��Z�3��{��S2��8��<�Q��CK=��� Z=-�<�\;������Ng=P <�2�*�O<�׼�᣺��F=b�{=���%	[�Ok��K��ϒ��KL{��꘼��<�[<�$���]=�y���r�<5�*<�XF�� �<�I�<��B��.{<�)=,��<�+�� Y^���2=�\d=o-<�8���L��b�J�漑�[==s#8�ǈ;Ȁ�;����C׼,:W�c/�=s����S����=��J��(�<7��Y=p.;=J�E������V�:_a@��Z�<��<5&�<�#D������
=v��<�aJ=(_;j��Q�
�l�$�aa�<k�μK,0=�XҼ���<�Q5���J=׮=L��;����)F�W/C�Eb=�/=f����U=F=d�N=�=��:�(o�黩�>���*�,/����<�_��R>����n=m3D���u;����/=4�%�$�k=��O<�M��<k�<}�=�u�<õ<7�C�.r���a?=@5P�fL�s]j=i�<�B��=�Vk������<��Q={A<�� <�O=���<�x=F��<�ռ�}Z��Z�r��<i�)�v��<�+��{+=�ba��Ń�F���\=���<̳���b<������'=�7�;4hi���e=6�@�R>�B�=�sй+��#蝼��~<�q��G���%Q=��=��$�J9�<�|=�C�<O=$(�*9.����i�t�%��n�B�=�=:�;�*ٺxwd<m���u�<�(�<&��<tpR= RG<��(�%lO=��n=��-����<�}�;�5�aY������ .��:=��K��:��S=)��S@��]$<ݢ����=�鵼僇�#2=���"2�<2��zb.=6�ļm��p�I=�,W=)�D:[u�<Z��k�K<�kL�^¼��`�&��	�2�G<�KD�t�_=!	���Q���^=t�=|�9��{3��=^�S=������<�臻��.=�ji=!#H�^��:BF�;�]ڼ$��< �<#�����|=^�:<�@�5��</�S=��,=� �~:����]$�ɬ��f^W=���GH�<�gټ��4=C4=/�<���<՗w��=I�o�0�~=*�(�v��^��%�ἱ�:������E�$<��<�==1���j�ᶼ�Ƽ<�e�<U�<�qR��S=�*��ֻ��l=�����gd�������K<,�� �[���\=H��}>=�cF<7���p����ڼ��_=�=[=#-*�9T)���Լ�3�SC=~��<�B/�P�!8��)��<�����"�<�5�����+���i<!5a����<�_.���4�{�<�	C��=ú2;Cb=�=%
�;(�<�%[��%	=�<���:�H��ߌb=��<y(J=��U=�J�"�$9�����(=��<jd�����-�=�6�<*_ɼ�,<�t�<��=�L���=�A�<�0�=O�;'"�����׀F<��I��6v<�==B\=�����H��G'=bF�H6��l�<���� ż��N����<�$= �=�XB��R=��=�K=<U�B�Mb'���V�G����<ZW<'GN���u�-R1�P�&<�B=��,= 4=�<�y�����I�8�rn9�i�4"=���<>��;%6�i���u"*=$P�4Ƒ�尻C�U=A�8=&���8D=�8�:�uM�ϐ�<��=hH�s��0�:�w)=��<ES<l��<@pB�iu=]<�z�$1d����:�yw��C�<&:L�u{��<�=zcQ�����ԣ<��*=D�=fU=GV='e꼁q)=�XT��L��2�]��^�<ֿ���N����Ҽ�NZ=����ɦ��`�;��0�	�X���(;�kZ<�;�D�<n߼f�l�7�9=�eh���S�s)<����=�)=��F=�A"=	w6=�Lc<�DY����H}M��Or<�'�<��%=_��>�O=�ya�u�L�;@(�/��<m�<���<���<�Q=��;灓��?b����<�$e��YE�fB��:��K�g�8��]=W�<<� ��� = (x=��<�����#��w��BCL=c^8���<�rR=�4[=�*�XV��A=:��<K�v=*\����<b �;9��겋<��C���,������2=�L�ן7=0�7r��Q��`�<Ċ�<БR�Hߣ��tμKj=K��pbJ=��;�7��<��(=t�'=�1R��=W_?��2�<�s�<%�<��;����^�ļ�ϼ�D=pv[=>��[���T=a�ü��@=q�"=_]���˟&��%q�7M�J*ڼ�Y<�V���f���<J*����<��;GtP�+�m:⛜<�@�<�D�b��&��<�E=��<��������+<�Ń<��<�f<(q =[(�<D=~�=��3<��ؼ�)�<��Ǽ�5��6v=��ւ���g=�2	=6�=i�q=WM�)p�>�=��'��=u=�L=���:��Qb=j�1=d�='��;�@=�8�<hz�<JR=�)��f5=T*�<}fû�'Y�Kw��YY����ټi=��!=6�7<A&ϼ�ꀼ*M!=yE6=m�E��ᵼ#�T���I�T�����l�D��<�v�<J�<oRh=��<��1=#�.�"z
=;e�����5=B��<��=�e%=��\��yD�c�N��=2�����W<9G=�h0=X �<��P<M�z<�Cp=�JN���Y�O�!q��ZL�<s]:���4�L�;�S�<
�Z��q5=��<;��<��w�Z��<�ܼDo=�Y#�KO=b�o=�B=�-^�N������_�<O.>=�?�;D�7<�o��ڣ���f#=��<?�^�1@=F�;KB5�G���&�<�77��3=�;��oZ=���;@�Z=Jz9;'.=4��<p$X=�q�M�����<L]<�:���5=vF�,���qK�FN=b�D=�x=�I=�3B=C=�*>=����M=�iz=Yi<	T/<�{�<��J�����2�=o,�9ҹ��8�z�Ҽ�IT={�=��j���Q=�oa��9�j�r=Vk&=����;��ڐ=Ⱦ�� c�<Lr#=�"4���<U]��r�8 ;	Z<�r=h(�.�;6l��S�<M�$<rm�<�D�<�߶�� n<�j=Oe���(=�=MÝ�
;���)�XDV�R�&�PӾ;!˺��7=��仼�=ӛ?�DX�<�;����%���;\'=;)���v)=J�G<�
�:�F=��G��C����o�=�˻��;�#�<h�"=�=���;�$ּ��˼5v=���,P=_���Y�>>M����<��8���<�bܻ���!��}B	��%��ZD�!���=�<�}�;�������=�P���C�<�*ؼ<;�a?���RS<]i���j=aJ=���;��"��=�'�<@$=S�<�6=!�<�3������< �;=	L=µr=w�<��:=&�V�l
=.�������<*1�d3C<�W�<Oc9�¸�<��;�?)=B1�u�;J8=:]��V��b!=|���Q���=C���0=J0�<�!=�O��[�<�@W=�!r<�T5=9#�t��<X�w�X<����f<w${����;?�A=�N<�۞;��j�K'�ZT~<�$�[P5=м?�E=~S�<�A(=�]����<�m�úN����;�@g;�m;!9=�Z��L<�`I���*=#/=e�ĺb�T�<<߯��GB<��6�CE�������Ƽ�^P=�`�<6QZ�G<.��<����~��چ=Z�����c=b=;��<���=9Rȼ�-�;���O=��=�g=�(F�{��;�s=��l��b%=K���JP�:���J븼0'��}�<�o�< "z<�<K�L<F���G��o(���="�d=�*�Ա6=������=4>O=+�j=B���LM<��*=�.=�,�<zr"=O��<p� =�q'�ıM=��=�T=؎$�q���=%�<J�x�ڢ�<�4�=S���.=���<-x����j=�y�<�׹��˺q��<R�';���<�y8=	n��Ey<�R��hG�O��a[���G<�u�<�t�<ŏ(;qӛ<b�<�����>�<�nϼ�d`=�	=�O=#�X��VB<�;>�����L�PK����  0   0 PK                    " 0 FIN_seed_148_int_414_head_4/data/4FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZp�H?�0=�f?u	">�0�>�E��7��Pm;?�{.���>��-��k/?j��>�V5?�!7?�PK���w@   @   PK                    " 0 FIN_seed_148_int_414_head_4/data/5FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ��'��tɾ�V��7>��k���t>�tH��v�>�>�x���Z�>�?��C?�8?��L>S��>PK��LB@   @   PK                    " 0 FIN_seed_148_int_414_head_4/data/6FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�a;�c�:R�::�<:T1;U�;O2;!�;��z:x�:@_T:���;ФO;��;�8j;q;PK%[�?@   @   PK                    " 0 FIN_seed_148_int_414_head_4/data/7FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ��==�j4��j=�o��/Ab=��;���<v���G����F=�E���؃=F�н}Q��Q~�+�.�v�F�IKI���=��<��������_��=�k��<����4<�����_�+2�;)(��o:x�^HT�u�Q=��]��{�/�;j~м4	f�AU7=��<�̺���=�(�]��ᡴ<�@�=q ��1ü�<\Q�<�&����ֺi��<n��㷑�y��<��t=���9 ��);��Y=څo<�b@�b|9<�<��}��)�=�%�=dX�=d�U� >�!œ<��<�=�\�l�=�L��_���R=��=�Cz����;yW`=Ѷ�����9>H�`a=r9;w���μ�,�='ƕ���3���<���=Ǎ��O����IY=jfz=�\ջ1�<�c��<����*F=�=EJ��Y
<TQe=}��<����D=p�
��)��o���ň�7�)�#�-���=�����R�;�v*=�-z=�b �u^�<�5�<̼ux8��=�f� �:83�=u_!=^o�ӓ0=��=M� =G@�=v=z�=z��=H���k���C��#}=}�=8Ҝ=�i���Rɼ�҃;y�q����^�=ʐ�<AtM<������;=6�;�A������G�<u1��}�G��Ů��R�=EV<��Ӽ�g���]���D�hd;e~�;f���&9��9��ةe�wӠ;Fɵ=�u=M�*���=m��(�<��=�Wd��WV�W��/~��Њ�=�5W=L^_=>��<`��<r�=��V=�����⠼|�(=]-5;���X)�<��p=�J=z�e=�W=@E�Q����<>�� �;���<1)=d��rd&�G�<��;h*w=˫5=�	���y=��+����=6Ӹ��՘<D
W����=�7=�]��~��Y�<`�=�p��|)*=�w=׎}�����}�%=u�.<0��������=7�)=�������a��;k�\��!�<{��=LÏ�9
��%��<�=�<tJ=6�:=��H<H�=�S��1�=��>��gu='�=v�[��g<JH9=rК�{/��`O=x��%�<��}=��J;t	.��=.:`�@�;�Ѓ�;�����=]�=�:�=%�;��:#�"=w�mӗ=U˫<Nl�;=K�ؽ��<�o�="�E��e�<���<*�<�� =0�����=U���aa��7���e=��g�7o��7����'9~���ʼf�q<�c{�[�U<Oz�9��c�X���Yɼ�4�<����,�;4�<�;�OM=G }�����ᗽ�$��6;f˳�^��̪�=�L=�=j����ã<��q:U�='S��Ě�'��=c
=D/ͻ�/�.��3��=w�W��2v90�@�s�~=s���Ǯ,=���<̘`�1�k=���<x���D��='%���ݼ]T�<;���e=�З��9<���t�)	l;��=Z,��K��S==�0�I5�;��������<Eꐽy�$��#����d=u�<�A����<I�<$F�=��=�s���==�w�;a)�<�<<�ӽ��{�AEG=1T��:e�a��<��=w~���+�=�d�<C=K��;Ã���=Zk��Kaz=�#=��<���<��5=�E�-�ݼ7*<(�]=R)��h�7K�=�B�=�.k�
��=-���GռCv=@w�<��}�5�w�Z��<w=:X>��ޓ� ��Fͼ�Xf<����&�� ؛���+=��p=�E��@��+���=%�O=�9*��<UD;�2^<[�u�T7�<���=t =𭒼�"=�==�<�>��<����+<9=o!�Ō���m0=�Hh�v=6ˁ�=4�=���C馽����đ���I=�{(�W�O�d�<%�=��=�=����$�=��O��]=*�=���� =�j��JR�=Hl��+��;$�=�����p�<'y<���	U�t|4=�=���<��=P�8�b
#���һ00�����;�<��<���;���=���g=��P��ы���8=8BH<c"�����<�"�����<�Ü=n�=Gh=0�<�E��!��+3�;��=dܬ��w������{�;��2��!�=U�= Z\��ɻ��=� ��P"=eb�=����t�=��y��$6��7��G�=��׼d 8�Q�K����=#���� �=C�u=,�Q=N�����=�7=�8=��(<��/=9�=B'�=㛒=�L<��=��=H(�X�=,�o��5���A��S������=�o= ��g���x��͗=b��< ���UM=V�{<ˣp�S�<�<o=�k��Ϳ9=�<���!�8瑼bBҼ?<�<b<�q<���p@;<�\�;h��d��=\"�=೒=���==`�7D���8[=" �����7�X���|=k̕�&�?=�N��C�<A�<J�q����15�@�B=��� ą��킽@U뼞<e��黧��<�o@;M~L��!��b�2< d��ʲn���V��ѫ<�͟=��O<{7�i��=��=>Y�<8z;��ݑ�=Hۤ<�gb�冽���n��<���<4�̽���<d�Y���<3w�^5���3=J��=x/=}��=��1���;f�U�Bǩ=�Sa=�Z=�=&f=Y=
�	:���X=�Sv�`h_=�\�.�;�	z�=�0¼hZ������=��=�Lڼ��D�E��.��gF=��y�����=Nj���Ч<Snm�}=����<�/g=L]O�	*#=|��;H�=���/�W��� ��'8=I�l=*[�<�`ڻ�M=0�N=>i~=�ˇ<�N��2��5OV�݅X��#t=��/���~=�޽a����������<��=�<)X=�#�;N낽;,C=���<��B=��=���=�c��b�<g�G=��=ji��4�<j��1��6��;��m=�3���!;;OE=�E����<����.��z�\<��V�CQ=��(=���������f=��M<x�y���b�=���Fe��"��^0��Z�6��.=�b6�0��=.�?=%�B=��b�dFP�:�`=]A�qT���! ��[R<��[�s-�����=�=������ֺ=�7=�S9=�r�'ڼ�4�����U= Z�<4�=-n�=f�d�T=�G=�W�=~
�=�F?;�9��h�y=�w�\���������=I�5��K&=�X���H=2D=�u��Ƚ��4=<�=�r=E!I=�&=8�P<$�5���K�`uP<I���6ن��M� ;aV���G/[���<��ļ��������bZ�cD�Q�m=3`�=�\�_�
=�_��I:=� =��<*"����H�=
U=����##��B_H=]�2��&)��E�<�1�=b@U���5=��¼�/Z<���<̹��0�+=R9 =���=���=����,��m����(��Y=N�a�A��f�=Cd=�<��Y���n�`��-���=�1�=�� �3���N���ýc��\;���|�I=?.=3%��m0���g�=9�l���=�fg����=#�V�kR������*�;/���˜=?�˽|�N=Kf<G�:�Ǹ����
��<:�I<�<׼�6T=m'��w�������<됽���<��C=�2�<���<�t=���<}d���nt<��c=�66�q��#�;&�.<�B�Cم=�!�=�N=q\9=�޼J*�=�K�����;I�a��g̼�G�<~��<��=7+�=<��=�Tp=�[���)�</����ɘ=v㗽��5=rB���푽a���+=��=E�T=��]=�no<�F�;��U=u	�=�p��Y=@W���׮��ԩ=�K<��=�=;�N<K�������k�=[xn�1����0�e�><��<,�=/�<�@��;�<�f��_3�<��=���<��=��y�pi�<󕔽(_�<sa�=CG��~(�e�L����=dvͼ|=o'��=Sw`=��X<��3=_1�����<vu=Im�<7�,<��=.Ay=�μu�.��Oo=�><�n�=�m���=�j=���켅P1=�9�����.��1TZ<�i���w�,�L=h؀=���=r���7�=��,=�����h�X��7�=�N���VM=��<��T�x����<�ژ=4���ݚ�|[�<JM���O��t�v�X��=\�=eU=٥ڼ*�=�'����=#]<�
��=��<`3�=S���������ֻ5�<�4 �2�����i1 =� W=Ƴ�=�}<u���~ �z�}=�ğ��������b�C=��2�Z�<gy�=�|�=�^=�@W=��<��C�hYD=�����;EM�=u�z�ե��rF�<�:e=�,%=�t��:�<6�Z=�Z�.��֨�=�Ի�;=ߟe=G����q���P�=?��<�*&-=4����q���Yg�J���}Y��� �=����׮;ݒ�'����(�=@��<jU�ȣ�������P���p�5�=,5><��<�I0���a��lx8Y���쩻�̶<&�=�e�<o�;dÅ=��Z��@��US0�!�!=V��=©�����;�s����=��	=
뛽�T'=�+<1h���D<Xz9=��׼�LE=#��Mm����&��<e`��L?�<|�=��=�T��n|<kt�;J�L�>�n; �.�Z%1�1�=����dj���s�A^.=T��=:�L�B]9�)ͥ=�_���7�<C�!���Ǽ�UR�>��=@|����޼�-�=r�ʼ�+��<�h��_��l�w=a˼�ʹ�%�I�+� ����¥���=�;���󒽀ػ���Z����E.�<����d�<P3#=�<��������,��*��Q6�9���_����=���HI=3Y}���M=ߞX�6�����=9�=g�j�/=��=s����b=��a��.F=�{<��e=�5�<��<�笽w`���@:=�t������x�S�_�8X/��A���C�а=���<ST*=��G����3Ɍ=L��=]��=/ռ�Y<�H������,g=����_�<��V�<����f�!j�<Z�<��μ�y�;���� �w<tP���(#�~6=>���Ϣ����pO��'���8��R:=�〽��@�����s��T3y�إl<��F�P����2���==�@���W���<�z鄽�|=!K=�=J:�<�X<���4�;zӨ���M��6�=��ȼ<oQ=������j����	ż��5��t�s���>�E=�͝�2ړ=3(�=Ϲ��Ba�<\��'���4����M���p����<A�=���:�u=�F�����(���#Vd���=+ݩ<v��8�����<�� ḼƋI=��἞Ñ��mx�Q��5�K=,��<���:��=G��Ś����G���R;��=���f��_��>�*=l+`��t˼��;c	h�=&;�'Q���,<���;#=.=2������v��=S=�<T�����(��}G�s�`<'��=�U�N�1����=��<�
�����='<�ā<��=lb�=i�3=���<^�<��˽ȍ�2���t>�o�r=#֮���~�����s�A=�<y=��O�f=5�<�2�=rL
��`P=���<oF�<���쫫�k��KQA��۞�kN=�E���,�=���0���6���	�Ѣ:�<�F=����؂=�9�&�u<�b�=np���z�=2��=�t�=�o<��=�p�=�-���]���a���'�'�eާ�c��<�0�<���R#�<$|>=�}�=И�<Mz�:����l��L���&VC=<������|�}�pjU=�����5x=����b`�����է=蚦<᎞=��:߻��`��l;��=S�$<F�e=,7�=O��[ʥ=;�w=~΅�������¥��6�;��o<sU�={����-<Da��s��=��J;�f��0z;��]=����-=���<q�N���b��<�e==n2=�+7<��R���J�7�4=}3��Gm���t�;�.O�t  =Q/��"����}=hPY��=��?��<�:=4�&=���ݴ�cm�<�G�<s���p=��<j�}�j�{�/���|�$=����-�=�+E��>=�;M{<k̓=Q%(= =zWj����;�ֹ�=��<��=؍!=�m���<�}�<��<�ۼ�]o=��=ÎO��f�f�I=h��Cd,</��*�ʼm=���;�<ܼ*?ۼ� c=�ٕ=����T��=� �=�ü=������;_|\=g�&=�߼6�>�gX"��n�=h0��a#����=��=�ʔ�-쑽��n=��=m�><�0���%��/p�����-��=R�P��=3	�=�t�<W�?<��j�����Y��ޢ<t��<��}=����� =0���.=��k�棳�n��;�81��s7��{=(-$=�)=߶C�ai|��!�=��L<�];�FM���=R옼�Z���=�#�=
u�;C��:��ҡ���k���s<���=6<=�,=�ٜ=Q(U=8�[�i�Խe�=�Z�SΏ�<��[�ʻ��=�۩=�1��3>��W�;�b�=�=&z=��\=����\:q=p��<F/��9�=΃�=�6��ږ=FEE�-��<�=7�Q��i�;C}Q���<�n�yR�<�p�����<&&�����=��=�~��5=�F�<�#T;�μ�.����~=�GW<�C�.^=�Z��G膼j�H�53���,���y=���*�=ϫ��Q�<�j�O=�>c���<��4����,�<�NV�˖�^	�</.=$�=7�z=�؛< ��M��u�<����.�<弤�q�(��<Gr=��#<�i=>K��_����x-=p_�<�F=�'�%8�$
�Цi=������<�M=<b����ҽ<��S��DX<:,�=Ec=�U$���E�"w���k���=�}�<��	=$�ѻ��J�<??=�]�=j�h��r�<�t��N��x�t��WY=�ǯ<�����Cn\;V9�;����`�D�2K<���<�#�=������d�����(��=�w�ǻp=^Ձ�f0<�aq=�Z���ަ=0ƶ�p(K=��E=Q���,W�<VM�=��'=&5��Aq�<!� <�*��T5�f)=��	��,�=��<(�=^�*	��I�p��X�$����?{=t�=P�����B=\j�=ѻ���O�=b���m����=ژ�;� �=j2���y�=���8�H<�l���;s=�I9��F=1�F=�8k<��`�4߄=My=�퉽K��<"\�o�w=l;a�9��:�`�'ɇ=)'<�9���=z�=�P"��C?=��=�����YD�%v�<�s�%�-=�ё=�ؼ�rR�4�_=eEZ=8�H�x�R=&�&=1����<
�$��@���K<�oR=fO`<�Ñ��3y�za��ǣ=C��<I9��#b=i����q=o[<��s��S,=c;�=���,U�=��=��x=xa����g=���<j'�+�_=�0=H�<��<������x���4���=ӎ�����9�<��=�z�< >�<�e= V��MHv��M	=�=`?�=#<�KB���]���i�s�p���=5�<W�x=���|hY=<뎼i9��Z�o샽�����Ҽ����|	#��;��g���tZ���;����(��ڷ<a���_=}�<��x���
��_�P�ܼ�.�=��{=�c���ȭ<Dl9�ɤ���i������X��^�)�a���X�I���oμ��:�76�i�����+=�Ώ���
<��<��F<������H�e��ӫ�=ӈ�=R�Ӻ�oh=�?m=?C����f=����c<P1i����~��&���<�?��Y=hA��s8���\�<�fl�4J���"$<��i=P�	��]��m��p3�<ʵ��=qO�<a����q�#VS=V=�3=�/�E�<���$�= ��<�|�\�3��踽2��t�=�O�<�,	=�ļZ��{==F�c=��n��'��`����~=VJ�<'�.�g`L;M�4<�<�=�7��ٲ=�<�7�=W/m�u>���|�=\=z��=<�e=��֨ ��Ώ��+�<��)= �;�<Շ�=��4�vN
<;�U��_�P�=��-�hc^��[9��W���O2����%G�;�b��z��1=]A*���s� �ǃ
��X ��cg<��<&w=)�<T~\�n�ɼ��<LP<�\�<�.< ��=VW���cۻ�ڶ=��n� ~�s��k%�=H��=� �=�x=z�<�<e��=_���~�l=�I��g�]����yX��u�< �j��f><�	�=I�9�=7=��A�d�=*$�=\�=�i�;�Wp=�ܚ����<Hw=��e��¼șu=�x��J5Ǽg�<*��d%��̽@�j����:�=oF��0��<�=ǻ'n�=���S�<8�#�M���Mʻ�וĽN�μ1�<6`|=�8��N��<)p����<}E�����Ż=Ao�<}0���v�zhA=�~�I������+��*���H"�=�˚�Ka=Ua����z<'�g=6YM������ic�������^��<L�<�y��q�)=X7��0�\������n�=в=�@�<q�8=�LN���<����+ڻ@Kp�E!@�<����Uƽ!�d��=�V~<�(1=$N=+Q�CT�=d��=��><��<d�=`��=���=�H�=�Y�;F!�=��=���<�?���q�=�����g=K$f���0=Pc����<X�t���=���FϪ���
��q��E�)������=ȏ��q��<�Ѥ=b_~��h=��=ޏ����#=�,q=uz����3˻��|<ڇC�ڿ�=��5=�犽wTk=�R=��<$��{���.u=��<Ő=�IH�|[$�0e
����<���<�$I�@Y�y˟=�-�����`N���A��ߋ�=�%��`����=Oz&��}=268=e����[��ښ�<�OŽ�;�=��[���=���<�!1=U�z���=��8��a<`{��E��<>c�q�ú�E�V��<���;��
�OѼ/��=J�]�<L@�=.ܽ=��=8\�<R�}��/����=��	=Yj�9��=������!o<=����%��7�@S�<7H �(�ý3�z=�"-����;J��<���XY�/2l���
=�=gvl=P��=	�2=iwN=$� <��=�<<�ݼ?�=�=O�zB(<��=0F�<^��<Eӽ%���n==��J�=�輟Ȑ<�����<	��=�=��4��4�$=�9�8�6��B0��Y��CΤ=�����<�WO=�v��=궼���<G�~=���<7�����;E�u=��=�ӗ=fߍ=ˤ�=<
����Ѽ�U�/�=<w]��4o�\��=X
�=�*ɼ���<�3�=�0=={*9�X=�̴=�h~=�|���Y<=>�=b؁�� �=�����J�E)R�Tք=�Cr<i���zI�=��;7�t��>����2P+<ä���M�;z�O;	��=���f�Ľ�u��.Yo��ˀ=e�-���6�`~@�|����+=r*�;�4�<��N��͛=��ֻ�P�=XX(=�Um= �{=N?Y=�<���d�~�k=̃<�#=҅�<K�V=-/=GHy={M=����_fq��f��K#=�q�E=ը���1����<��\��
����Y��ƽ|�<�\�=����=;�:=^���K�<߷p=� w=_K����<�0�=��=��<�=c#X=�B��@�U�<�=Wݱ;`[�=^�=��׻#��=s)=K01=|��=q:���"�=�Ej�g�wv=5+�=�ۗ�GP=Z�<�<�%��%:9���=��h�E�=MH��(dK=� �˔5��E0=�
=�>�<�ᴽ
����څ��3z��K&�Q,=��e�{	?=0�{<��9��_5���0��Ԭ=��=i�T�/KB����<�^=V�=�>��������6�w����X=�ME�$"��ܳ�o>��(���y���'���<cU=�eƼ�(="�0<�i!=Aa�\�;��=J9��2��=�?��p�7�7a����T=�<�"�J=���'p��O���_��C��::=x����5��ś=�K�=S=�SZ=��o=�Ӏ=z����D2�H��:d}���4<�X�=�L��1�q���8=�����B=*��=!\d=&���	s(�D��<N�r����2�=�]��cm�={�s=��,�#��=��;Kƹ<��;�q���)���f�,�<�E�����%�Ǽ�j����<��;�9=�Wg�(/����~�v�'��=�,�=?��JU�����<ʆ=ym~��H=��=��3���<ǡ�������~�lc=+�ʼP�o�%:\;���
�<O�=����+��b!=��`�s
h;F�N=�j�_<�<�����2º#��<�ⱽ?<�=�� ���<_k?�F�K��v=
�]=�ɽ2r�=�<��W<�$���/F���=�&.���7��<|����� 3�;�Z{<��
=b��}�:q��<rޤ����=]Rn=2�=[8�=Y���#<J�=�g�<�֔=�5<���D<1��=mŗ��&Y��'�^KJ���=W��ɏ������,�3���0�;��s�3��gH���X=��=��a<Qs��T)��2��	v��V��@�^<f�@���輼U��A���������)|6=��=3@=K�¼�\����<<�:=�rq���C;Ԯ���E�����=2zy=�A0=�����R)=�2=\��=�{�<̹a=�l<�y%=(��вK=p�%�ǚ�=a}���%=�Β�7WQ�S�=��p=�?�<�E��矑=.�O=��U=�wE�b���br<�n=H�=i ~=� ���7��GQ�+�J��c�<��P�}����w�=k�u�a苽�w<������;��=�[�4t=�q8�&"
=g��B�����==K۫���=��O��CY�;}�=�s=�J��,�=(?�=�v��$=�8��M[��\��f@�e��;��D������w�Oo��G݊=�Ƽ�c��s��Qg�=,a<�m�;,¶�9$�=�F =M��Eo<K����㼾ԙ=#�=�s��sw��y{������������`���1��y;+G��m6�-�Լ��޼W�<#�#��-=��<%�k<�<;n�=���=?2�=5�=�����;"�=C�<)�=Y��;Wr�=	[�<.m�==t������,�Y㤺;a��)=�G�����=p!�=�4T<�k!��h�
6c���=�炽��=��׹w6D�n⁽����C'���P���=x�������<��~�Í��� ��go��Xc=ܖ�<�Fi�Sm�������<lv;�@��҂���i�<���<(�#�kH�<�{�=�1������>@��[n=����� "��T=J�P�=s�ݼ�5!<�KE=Q�~�=	󪼢�<iǕ<&l��h��f�=�KR��CӼ�L.=��u=#�R�C�=���<��=m��UI�=��~=\]	=E�O��iռ���H	�=�
G=k�#������1��������<�Vs=�6,=�w%=24}���-�6����^E= _&=k�.<>��=K�[���`���=(L=Fz�k?� B�DBB<�m��c�����NQ�<�R�;�<n�H�i&�Ԍ�=>a�=2=q6&���<[�"�H�=~�½_��=~J����ü �=1�=���[E�=�&��e=ź%=w6�<�F��[z�=x����o��iR=7�=��z=��=��,=�X=z9�<6���@Ȉ=�Њ�\ժ=�H���x=)D���}���u\��%(�Zz�=��	:4�=��������&2=�ϻ<���xځ={����H���DY<�V=&��=��f�w=�JD=}��
�Tm��L�8<��W�<'�=Gv����:μ�=eH�=���r\ջ�1K<��?=q;�ļ�͂�馝�����8k�**<\���16"��ޤ=>_-�&���F*��2��=L0=�u�^X=�U�<k���?a޼C�Ǽ�	�=1V�<r��d���d�9�K=Ua�r��;Gc,=X�=>����.�=W��<��==Є��/�-=���PĿ�"q�=n$��O
���E�;�ɽ����_��D��=Ƞ켹�<��<�aB=�}p=qXq�z�=)"���=�6����B�Ua��p�=��t<��ټd�������'.;�#�	�m���;��Z�����s��C��V=b�8�;����6O�D�¼^ࣼ��\�v����)��A=��
�u��<�b��0{��r�ʽ�<l陽v�0��>��u�2Lw��ʂ<��O��b����K��#�Vލ=����)Q= ᒽ�d�=������VJ�=B�<)�S=,�=��]=�:�=RŐ=�պ<YT�
n��6�=D��=2����:�;�K<��""<��g��8�<��;����@ji=JR:��h����1=�z{���<(��*�<�=�œ��E�O=��<`�'=4��=�)~��Do��gs=���$H����=(��<<g�<� �=�=�����1�V� �/=V���7E����=3�=_z�=^��<��OSl=H�#=F�@=���=�,&�^�;={�ɼ-O=��c=�F����6ȉ�0J�<�T�}4���e��F@=Ӎ�<�\���;��r���=:�㼡k������"�1Z������٩l�im���O�<�AS<UV������g;<$=�}\�z�`�&A=-���o=RQ���K�v���M=ko/<F�5�Ik������a6�<�<�<�\Z<K��<�̜=)
��<)=�H=����c�d=��5;wC~=Z�����<�F=P�:��1A=��øNμ��½ZӍ=���=���Q[�<ɐ�<f$��i(�����<�b����]=�1����D;,$L�N5�x�P=1	�<��=�:�<o�<��=���<�=�o���8��̌<�܄��o.��U�<Ǝ�:oi�IfI<�\<WS=ČC=a�=׃�����ʼG-ݼ�]�<n��=�~=�>a<h/P���?�Hf��w0X<���7ѓ=H=� {�mF���2��]��w�����!��F���߼A�p���<q�׼�(�=w�=/픻�v:��A=&l=5Mq�] �=�ǻT�=K^=Gݜ�^���U�V���=7�<t�˽�)u=Dx�z�ɼ�!�=����r�W^m<����%�P�%;B�U=��,=�ކ��ߺ��J1�2팽�H���}`;d�<J�C�X/��Rш;�[=��G���<?5�<�3���	<���s֩=��*=�uG�����a�=}z���7�ou�J7���=�E=���<B�<��-;�W=������������C=lC�<�&t�ӘʼjoW="W����u��1=T�<�z=|��}}���6<�w=}�4<"=<�8�S�%�𚉼-!=�
�<DV�'����Ů��=w=C��<{�
L��s]���N<ͩl�$�=>�ȼA���ޖ��[K�<�1<��e:�0�;a����<�-�����LT��Y����=/6��>�Y�\�O��	μ|�=�
�y}R=�z�<�d�=�z=���
�=pr=���� I=/aj=�y��I=�	���%�<��A�X<g=nY
��8_��8�;x(��m��:�=�<����[��<��m����ԗ<t�3�fT�=����ץ���s=���Vp=��=�7����R=��X=�А��o��Ŧi�w����´;�L��1��%v=�4�v,���vE���|<M,=�� ��<# �=1�<��ĉ�#�=���=ǐ����,=)��T����5=Q�^�4����<��R��ڛ=�V���; �+��h�W=�����^�<y?/={мr�q=��0���=$`�<ۃ�=�5���έ�n��<kp=R�=�(K��2��"!=Oa=F�\�c#i=Da�=�D�i��-�<�g4<�y=Dj���E=U�w��h�����QK�='�����<S�滠u=Cg=��R<p�n��Ru=�\�<^��=\�����=OzB=B��l����@���"�oT�<�ٔ���'�a|�=>\�8�r=9�<�,н������-,���G��O���G�*�@�e�<��q���9=��*�����n.�GgK=_#e=	�==9=�A��{�<���W�=�ɡ=� �@<1=��6�O|��l;��<�ͽ���>�<��	=��=*�=�Zh�~.=]T������(=8#=���<�j�ef�;+������uy= �=IH3�	"��b��;:��<Q�=4�<1����1�^�ü7�򼽜�<�������<�:n�afR<��Y=���B��Ed���S�=�YV=�s7�z����Ă�g^����<���2|�<�yD���r���z��^�=al�<����T����:.</��=1%㻴�<,p�<�(�;��<u�]�g,�<�e\�v==3_.��H���+=�@�/�?=�8R=�ʕ�4O��oa=�4D<�l��g��C�%?=�h��G_3��	�<,�ټ𓣹(�<�f�=Z����9=Q	�=�D�=�ý�퟽a&=�N�)�e=3D-=�##=G=#���wY���<D=	��<��|�݂���F�<�J5;��<�z<�wdüOm>���t<>��=�,/=��<�:�Ĺ���g���Ļ��=P��=\ۛ<er;8������}�<ϣW���= �K=�4ɼ�ȼ<x��T�<ρ
=rK	�l�;l�&����:��<�4�=�l+<�����lj=�;F=~�<�S;
Y5�������u��9��:%��E�H�+(�<� ��d=����~�;^�V���m�< ����3�s=�0�;,���;�`N<�r�=��=~�a=���G������=q�����5=��5=�=��h�8��&����<K��~\�=�B^��%�#~=v�0=� ��s��~��E�U��a�����`}= ǐ��ڤ<Ӥ���kr�t=ā�;�U�=���n��D�t�}ѕ�_��֏<��-��Qż��k<���fmN=���<+��v���\A�=8�{��W�<��~=ߏ=˝���j��*���E=�O��Txe�hg��pV�2��<��<"Ç��n��ߏ?�a	�<�ŭ��?8:������Vn=,�(�އN=+�<`2i�Y�D=a=V�|��X��ۥ�=,т���;َȼ$_$:쑼�^�= ��<p��\P��%��䕽��c��=�az;C�<�-8���!:�C=O�q�5�=�=k<�=T�a��V��*��=xl=�Ȇ#�;4����<�`��o9=kq��Z��<���'���&�,<9�̼z#W<i���H2=m��³*=Mػ.^E=�<x�<�v�=����G��)n���߼�|l���s=#3I��1�=�so=s�=]}c=?4i=�м�N-����<�	������>G= H���Ԥ�U��tu�����;������S���_��2�=�:F<�>0�LPB=-o�9Gd=�����<�ƅ<D�<�y<iP=�w��z\{=���fә<��_;�M<V�K���Q�T�@��ڻ�h����ݻ�`�=�,2��B=��<��.�3�;�pҼ/�>�����N=���N��<V�=xd�<�<=:Tl�wp=f��o�����Y<21=]/�<9�j��"t��,9�aP�0�k;eL<�|%��=B=�w6=5�=-�<�]�����<����Vʼ�lϼ�K���Y�W#}��|P=��t����<
��=�����"� �<�3����^<	o=��~=�|z=,2�zo�<\^�rHм�j��!z�<Xf�=2�=g:Z=�}�=��Y_ͼ���x9��sV=US�;C?�=o��<�����;�7�_�����r?��~.<��=��=��<�5<%'�D��<��=��B=��)�LV���Ԟ=����O�]��W=�s=�=�F6��	E=$ ��k��v7��;�=H�����,��W=����$��W�⼹#\<:J=笣=�3��H+J�K��_=e����<��<�'�tq�����<�B9=Ǔ����<1���d`�يd���H��=3^�6�Q<7�κ	7%��LY=�!����=�8t�
�,���?�׬�<��=k��=���<�p#<�i=�F��z=��[<U�; $�=IӔ=2��g4�=���;�ō�ܳ#��|= �;=���<�x��SF<+�=�v��H}�;Zc�ԩ?=a�8<��9��:ڼ��G�����o�;]�!��J=���]2�����u,�<��K�7���L��<��p=߆=�pn��ͫ�)�/�!	#<ԱQ=��=.L/�쒛<��e=`��=z���ۮ�=G�мh4�=�#���5*�7v��|b=�4���H���h�d՞�0f=A"t��x=���=+�e=e�=Nـ�I��:��<��`=�@='�=0��<
�<&���~O=n��<��&=�(��\�=0;r<~
:��{:��=���֍=Ӿ<5��=
�<KlQ�YX�le[=�����:_\#���x���=s�<�{A��K]�uk<G
>��Ҏ<vP�=/�<f�;.}�����:jЙ�|*���_Q��ֽ<�V�81�-������7<9p!��"�<|��<�=��t=T������<ǁݼ�[=Lm=�{T��*t=���ܻ�<�?��A����r2= = M�<��3�A3��6d2�0��=��<�u=�ُ�o����9�����qr8���Q=D�d<��=���<^�<�Z��h�<8D���;�"��TR�2��BAC<�PP���ʼ�Ew<yh�=� =��3�
��)��vvS�W�=&�=3��;�=<���:)2�=s�I;4bH=}�$�<�=�曽�y0=����؁G���1�CL_����:�s��j�[�4�gU=��1<��l;%v�;(�n==��;��$=�6�<����V=j�·��s=n�5�==��O��o����=I;�;��?R���1�^/,<֭��c/L=i'�`�1���p�
��A��o@�<nvA=����|<�������-�^�P�C<�j�ɞ=��9+����;�t�����5n��/&��@�=j-��_y<�=~1�;iҳ=C#=���N���>�t�=�+����=ud8=c�2=�<>a`=O��<��r=��';�w"=Ph����;��`�<��Е5=/6μJ>���<���H�ԼE�<�"G�L|�=�������<��:Iފ=WE��ż	�y
�:�ɨ<�<�S鞽�"r<>}n�V^`�=g�����==N��ݽ��9�=��<�h��=���=nc��70=!��=u�k=㬗=!Y=8�<�cP��p�<�������:�{�=݇s�LV��C����{�^��=�=�P�=�����:=����������]�=`�{��dD�� �|ܸ=	�<��t��%=J��_�����U_=�k��H%=ĳ����<D�S��9m=��<�_"=`r=��<��M�����1O��|�X<jp=Hf�1�=s�=x��= ���W�@��<��h(�_��^%<�,=�;�R="Rg=�4=8�~�_���<\e=��Z=d,3<	�=�����Q�C.�<Zc������T=�;���;��Y=O=����<��a� ="��T�
��&W�.�����;6�
;�5=��K=��.�H��7h���%�<N�P=R<��<kg�=�bۻ=�����P=��=��뻣/��=}񄽸�!��K�<�t=����I�b���=.�=�=�3�� ,=NU";�g�l�=���=��=�{���*=��=�=��R�s.�=�ƼG,��(=���;~U����=���y<^�O��X����~^>=ӫ�=��=#h?�����=V\��a;S��<{?����<,��w����|6�=f�<î-=7�z=N]=���<uﯽ��=��=�6n=�t�)�]=�I�=�8E;�}�,����[λٺ�=u��HU}��+F�Fi;Qn9=���=H�R����<�"�c�f=�t�=%J0�&�=!�=�f��t�=��=(�w�����4�y�&�;G�=�x�	���n�:�7A=�#g�]�;&Ѧ;����C\�<؅�������m��yd=c�?=c��;�=>^μ�,�=S�t=t�=��s="^�����<H��=%��<Y�����=�G7=c3=c�R;9�K=!�����<���{N�=F=�wݼRy�=� "=f���v!=�ʼ�D�<���+Xw<�M��5�/=D�<�ܟ�;�U��t-="��=�����]�a��<Ҁ;<Wmf=m����=ۥ��bS�q�X<Z�&<�D<r�������di<�<�=�Ƈ<���=�m<���<�=j�$=T*��zn=[)�<@��<f�=c(=|Y�tڡ�rM��6j����[ҋ���={>=�ґ</�k=�d�=�\A=r�<8@=q=�c=v�=�I�=��.����-=�Y\=�*Q=��=�m0�3�;�]�=��<�w���V)�Zlp�^���=G^�=�_=��:�`ƻ5K�= (���aJ=��C�!<m�漖��=Gn��E�=J}/�J� =dL��>p��G̻��#��"1=����b�=��G=j��<�y=���i��&�5������#=��&=&���I�=��=T@��H=. ����=t�v��G��g�z=����)��<r���'���Z"���2�x��:�P\<�=5@�<p�}���=��o�=��<��=�oR=�ѻ������<'�������4�$�pޥ��?���y=��^=+����=�O�? <*�l=~:�=i2��|.�$P���@w� ����uA�C���%��<���Y�b�z%����.��#{<��c<eF�="y����t=i���䶄=�Y+��!=�����ڻ�*�#���:��=�&��1�C=Q�y=��=w���{�����;E\��뱽�����=t�i�>=:ž��y����=�C�;�����=.f�RM�=@�J��)E��%R8���<􇂽�lϼ>�p�Wy�=Ȇ!=.�0���ټNSG�PC��z�=����oI��%����@��"R�Vt�}����Z=��<��b�Y�{��Vq=n.�=�@e���輬=W�_��-!��Q=�GT����6A�<�.<�3�����j�=4��nX��j��^��=�ϻ�-�=Or�=܎�4ԏ=��T=����/<M�<mMY�=��0Q=Z�z�M�A�׵�<Y.=B���]�"=Sҥ< �ܼi�"�P~�P��<��=ku=������B�<e�� ����]<a�N<����`r�"獽�¼3�<&,;�k|�����Z唼u<�����^��)�=d�w=�<.9����<������<@^_=��w��=x*=���<�dD�W�m�\��Ą�ݍ=����\r��s����98�d�==r�w<����v=��<U =;��5�2)�;I��=�\�=y�=�%=��o��
�< ��=^�@��>{��q�<��N��ݎ=��2�E<�z�{�Z��f����k=�����;.<����l={
p=���=�L`=l��<�h����R�Hd�=�p��2)=��z����@�R�o􇼳��<�[=��+��jؼ�3V��w=I�<�H����<�!<�yf=�e�IF*���=5��5:=|��=��;`W>=�ý)���PFƼ���=P��	�K=��<yJc�>��=N�=�"��:T��������L�f���u�=�:<�\�=����W2��J�=<����)缡��=1�i��ǋ���S=C=19<_� �d���е��$K=�\=�$F=ʣ3=���<��`�!邽l����=��
<�=W�=�����S�4�������=��,�E��<�'=G+�;,0�<�G���u=Uk�<D�C=�ֺc�\<�==�=��͵�=�f�=��k=�� =nἵ�.<aV�<�C}�����&Å�B�輶K�<��4=0����<����D7�Ȕx�M�.���=����M�f���ݻ��,<u�I=��=��.��Ӌ<�AE<3QZ�?�"=	�<(^m�������=<��=��=��@=�ɳ<8kD�tZ�
 �Qxh=����l�=A�t�6�=v����̞�n8ݼ�g*=��<���{��<7��q���a <A\�<��:8�~=��+=�=���=^�F�Q�M=�k�����<Z����=ݨ^<�=�`������=U�P=:Ɵ=�q<+ҕ���n�F�;��=ջb�7<r|�T^y�:��<��<7�T��&<�J�=i=�ϲ=�>����f=,�<@�=����-<�<�b�S� O=QL�;�L�"y�=���<9�2=bS���S�������<�3�<%�p=,4+=�_�����;�&�������@-����<��<W����Қ=��?=0"�=��<�/?<�D���@�K=���=+�b�v{i=5�r;�ܴ��I���B�$�ļ�"=@��='��D�=�Y<J/���=Lvf�s�v=��B=��:�Ԥ����=i�a���D=KN=��V�I=���٨��!3��=����W�=c~ͽ���u����;ռ0�0=O�]=e$=�\��*h=f0~�@
]�r��=������@������" �=�����Y�<Lķ��$8|l���Y���r�p�<vպ�&�=�mW=(��=�0O<�L2=Xȼ
|<-��;�<ۜ�BW<<�9�;����
n��"���&<+��=*[q=D�������vQ=ꔥ����cN�����"�<����K�L��R;=����Z��g[=��9=}�=	o�@R��h�<����I%<C��=,���N����=/�q�49�����Դ�<�7߼A�y�.ڒ��8=P�<�V�=�$�������>�+W]�ٺ�����=HA�)Lj�]�{=h��<<�=���<�ؐ=�p=���<�{k=2n=\y=�c��m�<�x==��d�}t���c�=�?_�b��=���=�����_��*Q�����5�='�U=Piݼg�N��/��,�=T��=7�=�o=�~=��<��-=ng�:�B�=�?=�6=��G���<�<���,��ʢ�;�	<=k���Ϡ��8��^<uѻ�Y��� 4=��=��ּ
r&='�=a����<C�V�J��=�20�N�ݺl1=�cj=���M�:=%�r=HW.�u.W=	�����<�g^=��׼�򸽹'%������Me<����[ɼ�����p�'͠=����*==l�n�E����F7<˝?=/�ŕ=���<%������=�"-=9�N=/�!=;?�=K�	=*0��si�<J�$��DG<���<@��w���2=��㼏 ���>�<�=�=ʴ�<&�g���̻�,=�0����<Fd��=V��;��2<�E\<�Z��ڔ%�}=聛�G�>=4�܄ͼm#׼4ϫ;���M\����=�K��VJ��,�=Y�\=ne=A.����=2x�<
��;8.���ԏ=�x�MS�=Ѯ������qi(=����8��j�=���<�m��6_?=\*=�w=�_�=�z9<��I=y�dm=-n�=h�k�l-�FN~=ԺL=鱀;�n�Q�8��3�Ҹ-=I�ؼ����I�a���	�<rg*<|��ޯ�="�:<�!8=��=kʼ���:�"L���,=�x��\��v���O=(�T�L�y=�C����U=Q�Z=�����EP<�c��>L���e;��<_5=�`;��𼳀-��?�Eu=A��=��̮���Ӥ�ǟ�=������U=ޖ���Ug=WԜ��={�h5���	=	��&����ޛ=��<*�]<v� =�<l� =�<1=c�I<L���g���O������݈����kT�=��м�3=t߽<m�<�[`��^���,��Q���핽��O�()�=S�'=��=��<��;i���2����;�O;c��P �=u���z=��= �ǽ����C�2���[=�0C�\]�<�4?�ﱠ�l0��5e)=�;�;A`ѻ�b���_v�}3̼��=�A.���G���<I4g=�8}���u;�4�:��~=-����d�\5�����L#=Qo�<��̼��g=#H>������K�/m��:=�پ=�i�=��ü�R����v���;�k�p��N�cg7=��`=8��7�=����OD�X�m�=@�;��!=��=��֢<��|=P=Ue=�0�/�5;���<E�<�����%�9���)�ּ�?�=�VV=����+�=�:m=����?��=eQ�� _�GȆ�16#�(*���=��E��R^<nrc�ii�=���=
���G�L<o�Q=�+��ځ�=�,=10D��3 =&�伎.x=j�M�=I�����<Ev	=�]=�n��
G��P���:=��ƽ��u=Oμ�w�0&�=:%�;�g<={�k=ұK��A=��6@=�n�ӯo=�?;H����\=Zє=a%�=����h=�{�l�x��P<���<�}S�.�=��a=�o��\��<=q�<�>r�a���rg\=`��ʷ�<_��=~���m�=�8<ɻX���i��&x=p�=�{�<�἞��T��=�㍽�8�=��I����=][D�V�<Ih��"�=�.G��X��LP�\;�ۅ���n�Ԟ�=���<6]�=z*==�ͼ��l�LP^=�2�;���=�3��'=��=�ܘ����U���YЉ�V6O��ހ=�PD=�|/=��5��Ė=���i�X<m�<�m�S4,=~x;/y��MS=�X2�Z�غ���<�����<=�X�0��=lF
��W鹴?���`��"t��Z=�� "��⻽��<=�=\�^<vP�;k� <�`=d^���<ˣ[=� ��س<��j��L� �z���p<��.�4p�=V��<��Ǽ��=��{=�����tP�7�<�����6��u�:6S������Q=�qg=z���;��Ϲ<r��������<k��<���U�l�|�=�s�>c�<�ߙ�i�˼�_㻶�<��=&����F=n�8=�v������t�z�w��=�N0�c��<5"5�s)���S�$񨼝Kw=dwQ�S��8Ʈ<]Q<=e	<�RI<�z^;�=��<?z��o�<�T��t�P=-μ�{/�5��<j#���T<�,I�AC<�
G<ˁ���3=0It��0)��U*=��=���=���\ļݢ�=ق���]K��ν�l���w�<�]=	�$�6�=��}=x��	��=�w�=���ª���}�=�c���X �w9�ELk=cZf�2'��s@�� �������lGv�#ޙ�Oy=w�Լ?���»?_j���׼�u=I����ߟ<=��}]=w	�������L�H=2��@���:��=��=�/<.�=�
u���=��|=�zS��2N��n5=�����#�/���#���˺VG����<���>�r=�(�oc��r���a�=�e@�������d��:j���=��=�wR�8k� O}:Af�=�F;Q?�����<^|�<��ݼ��7�~��<E���.��]�m<*R�<�^�9���=?�<$�R=hW�=�7y=��ƻ��=I Q=���=C5�=63m=�v�={%4=��=KV��aFM9�×=�/��)��82�=ޚټ�g����§w=�B��?�⼢�p�*B��`l�<��=n��=��=��'J=�nH=E9������C{< Nk=�C����<� 4������6-��T�=x
�=dI��Kl�hr==WО�'Z���P=���Q�"��PO��|��˿�<�W���`�������np=/]������Q�zHK�q�\��0���Gкeѿ;Q���8�k��ȹ� <f�^=F�� ��<�N1=�)L�>I���	��cm��^�=�-��ݼ���G�Ǽ;*��l�+=�s9<��:=�6�<�5�����BX�<�}�*N=�P�==�E��%�=�{|�u��=��.��W)<k�
=���=���=<�@<����SZ=3=���d�۞�=��8=߹Kr��#c�=�^=�O��v����<�B�L�Dy�Xzr=��9�T\@�ئ^�S������r=���=�Y�=�z�=�L =E=R��=���j��=a�n<3���ڧ==����в�<��<3�=q�=�=�u?��W!;���*�7=A崽x���<e ��B�==4�$=H$ҽ6�<Xh$=*�m=������b<�̗�ծ�=P�r��+�=7���=WC=j?=:�`����<��b=c�<Ͼ}��cV=�ߝ��V�<?=�落0���G�񻠽m~.=+2��?>=G��<)G�=J���g5b=���=�S=y�:=�@���?=����7e��l3F<���=������<c���'��</�"<�x� �����k���Kz����#=��<�J���8=\�$=��?=1�O=�W��(;�Di���2=Zba���`�쐣���9�^ǰ9K|�*!��9=L0=OR����c��n=:}=;��b"��8���f=�í=�ޚ�$2;<��B��u&�|�<���<�׆=,�ۻ�ŋ=84���{<�E���|u�X2�<(<V���<f>]�k�y�Й;�l�?N��O�t=��b�1q����q=~@<ET��W ����=���=�:�y�I���Y�@53=ڧ�������˛�>���D=2�ik�}������BgD��ü�^��b$:��<�
�=��o=ԯ���r�=/VR�I9��"/�=d�����<�F=[�9=��=̨ƺu�g;�r�.n�< Y�=�M<�p�=sۂ�;<S�}��]=��(<V^��PZ˼�Cм��<{0���j:�+������<�v�=h�3�g=�	�<1��B���kj�<�=�x>=�@��=WY�`�q�0�����=t`=(٥=����}L��A�=얲�ND�=D"}<s���Л���t?='���ױ<0[R�j�O=��c���=�z&=|N"�Z-�=NdʼJZ�Q���k�<!;�<S�Ỏ��QS����<̖�&���@�=��0���\=���*��P�;<༛Q�<�˖=��J=�rs={�=#>캚ʯ=��I=0ɐ�ӥ���O�=�a=���<�ܯ�T��<��<����<�7=5�μ��`:L!;	��4{����K�V��ҝ�<u{�<��<�7O�!�n=�G�E�=^�F����v}�=�J=����n=��C��<��<�*A=y��;�f=�|+����%��I=�/��Z�=�M�6��EN=��Y<�˳;/f��5�=�y˻2衽��H<%����2�=y5]=��}���w=>~�-w¼4�/�u܄=nww��'�$l�H7s��\=�5�=V��<{�Y=���0=4����~]=�=��|=g/���K�a�o=�<�x=�ɖ=�k=�w���@<�.'=h'�=��Z.=`H�����x' =@������<��:<CɄ=�Ү<�R<�.���J<}�����<7c̼õ����O���1=cG?<����9*ڼd��L���l�=<�����=��R���"�P��<3����;�[���yUK=��<��l<����!<�5��	v�<�1=Q6�p���`�<荴��,=ٗ��9����=�p�Ծ�:�^]��(<�r=$�������](=��-��4��H2<34�<��L=�R�;������S�=B�|����˃A�~�=xwμJ��<��2�E��k�ǼEo}<��]<7���&@��*;�?_��NP�y0�=.H&�_g(�w�=�#=C�(��ຟ�MPc�G���� v�|=ߊ�ÊH<r��=M�D=�{?<� �=�pS=���<c�L=izN�}�]��ތ�Ϥ���ϊ=rP,���w<�1�]����)=O׵�7�=�o���T<�����2��x6=�χ=���<p����=�Z��8����L���V��n��c��;��=\�d=T4J���c=��,<��<�0�<&�}=�r,���<|U�=R�ʻ���=. �io˼ۜ�<�s�<OAN=�[���j=�<uXL����T	D=hR��%�Y=��{=�N�<B�[=��=@h����5�iJ�����#�<��
=� ���=���;Uy�<���<G��;s�	�1�=^l��w	ڼ��Q���^����_��cX��e��<J�<�����=�s�<x/�<�*=�/l<?Y����E�;����;�ݼ�K3=�J���������P=û��ҫ�&N�=Id�ɿT�D����$E��sF=!ZF<�X2���λ�KI������<���;�`C�~��=��E�Mf|;�='����l��\,-��-���oܺ�9<��</��<�/=� �:"����x/b��+=�	z=B��w����5=�x�=�+��֣==Ê�/b��r�8�0���;�=���=KϼRY>=⑽��$<�U= �<�k���=���2Z¼*�K=��P�ML�=��w=\f5��dt�Gb�<7q�=�8=��=g�=O;^=��U=	�=3=�]=?��=��*�5���������e+��ӓ<�x;A[�;�m��H�#m=3L�����E���}����+=��R��������<L$�|�h��H1=��e=?�S�\79='�l�T��Z�����2�=9����G;�!0�?n=�^�=f����!�#v��/?�ʍ]=H�a��sS�\됼�p�����[�=�(-��<'�=��G���Q<����~O==��=oE�9��{=�L�s�j=NW�;�zl=	�(�kQ���e`��G=��u=�==���<Mpj��w=��-=�	��;�����:z��8�G=���<�j�;�!r���=�A��%��6��=��L����;�8�=-�.;3e��"�����D=_ݽ�	`��4$T�~Px�<~�>1=�,�7؄���/���7�R>��nǂ�8&<��&=�P�=s����� ���O=�R躽Ǘ�B$��?=�h��=f=�!="8-�PF�d���k}3;	6ƽ�����`=�����{]��j�c�~�[!M<�=V�^=]/��I����'�;e	��vl=���<;́�J�{=f�=��=U�j�a�����7p�=Ȫ�=��=6��;�-�{qM���=-�V��j~�<J�<X��<��<�ۼ�pn�7�e��Fq<ߥ���%�\��d���P�e
G=X5=Y��N��<h����+�J����K�t��ß=}�>=A���ɗ<�88=���十��噽�I����	��)���<�=oc��֢-�ҷ�:>�5���A����<��G��S����#����*E�=|���U����w6�ڃ�<�Gv=hG<�ǼҦK=�O���[=��f="'!=�'�=U�~������iR���7�v�p� �v���;=�,�=�z�;[Y
<�,��{�==�O��f�f��xʼ�?2���d<iH"�T?9�,aI=mS�<vo��M�S=��=l���S�4�a�Bk���	��P�� �<�	:#p�:粼���C� ��=���T?�,���漳�/�{�<q�d���;�<�W�=��C�D�8<�,��X@�ߎo=�=�yh�d� =�n�=������4;�V0;�����V�<!�M��K�9�� :%�r�^�I�U�<�x;�K�;��|��%�Ω�<	痽���;[�V�5?���5]=)��<�d�<-A=��ڼ{���/=��{<��=׼�=�)@��v��^���~��<�g��/��<n�=P���f)=||=��=�=���!= �5=�o�<��<Dq��MTu���<[$W����=�e���r<g�;j�H��V;W�ȼӉ3�;%s=�bz=�����:�I=S�=�y�=91�}��<c=.=ւ����K=5��܃=Vn=��w�ȕ��8�c��5��i�n�SO�=�k�=R,�=A���Z_�:ka��{Z�U�;y�==��s='�jn<8��;��9Ӳ<pQ���ٍ=��V<�p=�����?v�Y|x��Xw��=,�=ܬ=&pȼ�l=T+&�tY���q�ϲC��Y��ɼFx�����Kȼ��a�� ڡ=X�}��M�ii�b4��в��f"=�vƼ��a��oO=�}s=�:m���=v�<�I�����㻸�Ң���s}=�_�d�{m��ns�=�s�<h0q=��L=�	����<�N<Y�;��l=���;kFJ���F�d�R��P�ǫ=��=�-n��eM��J�$=��
<�f`�c��;Q��<��i���ǻ0��=���!�����<�73=�A =ֈh=�d6�MgX���9��R=�4���u�Nl�<}�.=��<��o=�=:�<��6�5�!����<�H�<��:�=��;=����A�<���<n�<J_O�p������H=
_�;/A�;���<�`����*;�t�O3��#�p��"���	< ����t=y@�o�����y=��C��3p<F]Ǽ^�y=��O;�P���`=�$�>�J���=f�<$��<�����l=p=�ZL=gIb<p��=��(=e�%=�4���y=���<��Ҽ��<��v����<��[����9F������z��!�:�V�=!�=��<l�������=�jY�ќ �<�
=���<w����*{�Y��;(9ۼ�ڱ<#�����E=6.=bO�Pj�=��үG=�3�=&�W=KeQ�@-^�N�i��==���;k���cV������9��=��������U�K����b=Y�}�#��;���=3�F<���K{<����@���R�<+֮=t�%�@,m��J��Ż�S�s�C�=#�=��*=o�M<~b�= $�=�b��		�J0;����<��g=4I�<;Ѽ�e;���<�Y=P��]�<���=-G��;�=g�;����=�k�����-�y=3��=ZG���=�ʽ�pz��L=��=|�F=,[Y�f�=�N�<T���w����/=�=�u����L=*'[=�m=���<Q[��Gq�e�M=p'�<��l�7})�JF��q�<'�=�?/'�_=�ņ<f���m���2�<�������<Q<��<���c�#=N/=I�=�ŕ�fn=�폽��=�D�]��������;��l=�(�=b�=ð�<�6=��O���L=T�{<N+�<��=�>=�)��'�=�;@��(1='ľ��<�A�u=H�:Yք���]<y'b=ۺܼ#�����#�=B�Dε;��K��pȽ���=�v���vJ="��<�Ш��Վ:`�Y�T�� �<��=b%�9N�=�(��P<�<��n��Q�!@�<1���B=�#�q�ʺ�M=%�������F��\�z=.�<�P=��=n��<���C<��m����G�=��"�3�=,�4=�"�=&��<�:+=�L�<~�P��˗<��s=�)Y=�삼4՟=b�� �,�WE@�攙=s��<]����lĽ3���	������<W}�J�=��A�eO��*?���f=�����c�;tiz���ݻ̍f=:G�r��V���t���+,��\��=�kw=������	Y=朩��;�NI<��P=�)2:3#��#��<�Z^=�E����N=e���=�.���ܼ5$���qp�[��=�j"=
"V=U����V�<��X�$2�97
����=[à=�c?=���-ه=C���.��68<��Ǽ}�=�U����~�Q-�<G'�<���r��+&�?�p�P���WZ�|8ƻ���� ��D�<>X�@.���{d=4�#=��̼Q^�;�Rh�0d�􋳽;��=GrE�P8 =�О=��j��胼o0<Q+���y�
�2=cղ;�Z��m(-�J�=����ऽڒ�:��'�Xue�K�=t׽�~����a��<�q��"��<�yh�9�;=<���qA=qs=�x=�,�<�5W���9���;�x=�c�=� ���=zX�����T�=��=�1�1���?�<!�1�"�(=u�|=c9軣�k����=Li�=w��:]6�l�K��'M=��L��a��x�<�Ȇ;f�ݽM�$=��� �;,_�9Sᇼ��=�d�%'���=J",���i=�����=�= *�=ӑ��R�a�4d�=9�<qbn;J-���O� �X<�1�=�X���<S�K=���W��=����R�'������`��}���b;'V�<,�%=1m'=-�=��"�D�@Y��� ��+<=���<7R%��`=�ϟ�&+<�x���m4u�wM+=��~�'�=������[=aۖ�cuG=3�D=o½L w=hO =.�(���|���.<�� =���X�=ٍ;��=9����<wV�==��=��=n2��֔�<WtнQ�=S`�>Q���6˼�<�GӼ�U�={�]������Ž��d�,_�<y�;�s��
���0:��:=��z�|ډ���<9G=��P=e4����=�
��b�;r2�=���RM��`��<�|�=��=-|t�ن��� c���X�~�U=�OS=#�7=� %=״=* 	<Pq��{=����S�;j�@��J=(.�=�T:��m2=�ć=�uB=hY��tI���z�ꟻ�żCg�=֖=J=%���"=S��Ç޽-�t�X]�<%;;D���.��ѷ꼎F���i}�_ƃ��Zn=֓<Ι¼�>{���f���<��E��O=>-=���<�I`�Gp=����N	�ܟR����=��E��xQ=Η`;�<|�'�{=5�I=ऄ��Ï�������<����Ү�F�=�v�;�vP���φS<�b�<Pw:��������A�vɱ��z=�=���<N��=~\4=U�=7B�Y{<JU=����k*�kĀ�R=��޻���l�"�@8i������=�I���2���</��=i`A=$�(�����\���T=P�=0��<��(���W;`f�<$Y�=R\���X�H�F=[$=�{���ʋ<f8����R=(˲�Z�绫2=l��=4��;!s<��=q�ҽ�P̼.I�� A�<�*���=/�̽5u»���=�2���M=��=�ʼz�=��L=�lR=�C�<���N=9��7�=4�4=uN=���<�w=��j=�=����<�`�S=D�B=
l��pJ�΢��=j��}�{�?Mm�,��<���=�=�ɼ�]M=����a�l����=��н��<�F��pĊ=��s�^��=�(S=+�}=�(�Gx9=
A�H����='<�כ�=Þj=���<F�;�g=!=v�e�������Y&�=j[��(4�=�`��9=��o���=��h|<����~�U�=!j=�ټLF3�WG=�w=�d�:��;=��-�+}9��޼��7�xʑ=۬$=�=<F�d=���;�_���=�S�<�'0��C=B�=�=�Bż G�=��:����$��>��#��=�� �=�.=*]F���r=F�4�]P���'i=~�=A��<��6�ETh���鉨��b=�=���x@�=�����x��O ?�KIj���=�GS=��[=�>����<=��U�=��<܍Y=~k5=,S�=��%�0ü wr�(�<�+�%�?���#=<����{�J�=�T�<)���$78;�W�%���+=�����$d=+��=�W =<� <tNO���\�.s�W'�;?Z�=3�j�/��<��b��\;����<�z�<���w <i�><��=�۟�L�=�J�=8\i=��ʳ����<�z2��왽�6�/{�<$;!�9B=�6��w	��؊=	�9�OV�����<�a�=�>V��B��ۻ~�<J�=�!�M�W���>����Bǽ�	=s��j�P�����E�`���1����r=R�m�!��=.�A�X����ԗ�����w�F=l���C�=1~�=�D=�rS���#��=�;<��,=�ɼ���@V:=*��<�T^����;�}�y=�=ڽKſ=�� <�#ݼ̊m��k[=<n�<�ۘ�����BK���:=�X=h��<��<�0=Q5ڽ���M_$���C�~�=[��<�\A���h�����\�յj=)ْ<)=�<�MyQ���"=��=>#+����=�e�<ʃ�=[���Q���s��W`=�ކ�R���t�����ּ�^="�=vZ������$���F��4=���;K���<�=c��=����'�<=�o <�L�V2n=9	�Fi���&A��ν/04=��_��Ԛ��Cɼ��2�Y��=䇶�Xӯ<$�x�7g=����T=��ּS�z�Yi=h��<Rg����=�μF����}=,m�<r�b�b���F`=����ڮu<(��:E,=���<�o�<8��=-���E��II�-�n�k�:�9�<0��<�.`=g���߽u���y�_�w=�.��&�-�d���W��t�<�F�=L�T���:=hWX=	A�=��=ڂ��ßp=��H<D�<��<��<�O�<+��<�B�w��Fk=�C:�x�<=BƼޥv<��`���̽`N�<�<9��D��K=��=���=��;&����M�=�	X�r�b;;�)���E���<���=�=l׉�&_7�� �=	�;�����ǌ=Q��=B�=�f���=>�|�0�ݼԒp����=t*��o==�ӕ�P��=w�������8�˅��렽���i/���΋=Ї�<�(C<O�q��Ȃ�:#�<7�=�0�=v��<=�=���sR�=��Ҽ�w����s�g��<���=(�=�
=�`R<n=���X�{=;jC=��d�m�<�$s�͆3���r��o�=��<�ꕽv�|="ߙ��g�=���<kl=������#F��A�:����=6���گ=������Cg=�����E��ru=)�켤���>=�7"<Iͬ�n�='-�=�>A��^=�ߎ=�9j����td�<^n�<1�#=�:�"<���(h��>��<����
���Z-6=��鼈�=K�����A�F=ƪ�-����}�!����v�{9*�a�8=�d���=Q�<���<30k����<�'=�&�'~h������)=�+���XG=�EB�ٍ���x�<X�<,U�=�b�<�<�=

�.��ϭ^��LּF���݆�;`i=��w�V��gY=ZE���M=�2}�-~�<��=k۬��<�>i=�=�!���]����G"���>�����<2��=��J=��e<^�=Se@���-Fż =�ҙ���P���6�<^纽��=g�=�J6��]=�|ͼN�=��L<��<* ��:��<�Ɛ=�mu�4�$�!��<�^-=�A ��h�!*�<��9=��9���=����/��Z�
=�������ba�MI�Ы%���#=�.��0ռ ;q�=����vּ�t�������ۼeA�4�=/Q>=z�=3:׼1�?�n%�<#�<�a�<c0��g��=��<�=�.�<�����:=M��<H}�����6�A3<���=���=ș{���=�]Ҽ�0.=����=Դ�i�V=Cf�=,2F���<Ye��lF�C<�ƅ�%�'�;�o�r=dI��}�sh�=�<!�;[輓�<W뉼��7=��û�� ��N�;y�u=C��\33��,���<�=�<�ZT<u<�=�4ɻc��Uy�<i��=e�{�8���d�=W钼� �=��(;��=��0=\
�<�:���h=Ju�<7�m��_�<�e�<F�==�z=��=s��Y���l-=ҝ�������_�=���;Z�6�.c=VJ>��V�<��3=L�=��Q=$1=9ı�r?�p�A�qW��#ن�c*�<�!�ܕh=�BQ�&�w=q���᯽A�߻�.H<{��<Niw�Ѷ�=fk�<�Y��3��j%=%�=�d<��W=&��=��0��h�ߞ����=X�4=k1A���=KqW�ufx=��8�%\=3��5w�c ��?���A��u�;$=x� <�|�=h��<v����\ �%<=���`̼�����g�1�5��K���#z=<>�;�=�Z=ցT=�"���W)��t���;ϑ=R�=i��<����@"=D����=b=�hk���1�����|�;A��<4�M=�'���[<z�����<��4��F���M<���n^�<�bg����6���Epd;�r�*.;��S�0�����<����aH}= /=�1�:�0����n��=tO�;��=�p��2�<"2�=���<�곺+�v��;�H�C��=u5t���L�۸�<�r�<�"��`�G=��c;z�o=`��:�3d=��<֮�$�_�'�O:Q�h=$ė�EW!�9U<[��7 -<oĀ=��=!?y=y5=P�=
J���f=e�D��Æ��#ͻLc���<�=ZؼM�O=��;6u=h�_��(L=�!��4t���:�r$<,ś���:�m���4�!2�:A�-;�B�cnX=m.�;�ȧ��{��,<s=%b=���=ed-=��Z<����Ibμ�:=\V=4�E=�uR�:1/=�6�_A��d��mۚ=tf�/������*�;��=y�{=b�A=g�;3-Z=�⩼����J����f�=k9�=s�<lƖ�6�=@����&= ��=��n=Vo=�����^;�ݩ=!���5���=K��<�Ii=��*��-ǼǬ����=��g=g�2��U�=N)��L��c*=�@=�A��n
������h=S�?=y{�1���䄽��	<ߺ=M�=�8-=�8O�<ǚ=��<
8U=�����<��G��9������4I����<l��X5��;/�==��<��i��/=��=C�E�z�r��P�=����d���f=<	<|'�����<̍q<�M��=u䳼٬������/����><Fe=M�g�*�\��=�Ӈ�kG����ͼ[����vX��6��cJ�̄=;�!��b��3�a���P<ث�<�����˹��m�<0�����4=k�H=��=��E=��<��꒽�c�)!h=Z0�<8���yE�=�3��m(�gp������=�Wm�j<��,<
�=�}��4�y�}g,�_޿�hW��P?Ѽߍ��7<�%���g�=�3�<P�;4���G�g=m@��]��T�=2��2b��2뇽��ۼ���<{��=:ż�� �[P8��1��)�!��|S=w�W$��`�����.���/<̵P�Kђ=�_��N�4�8��9<��=p8��e@����8��O=����q�?�0�҅���=Zy�]H���p�=FO�<׈'<5��= f�=�|=T�8<�i|<�6ϽJau=�A&=C&�<���<��J=�G=�| =��^�g���e=��r=KU�g^&=HZ�=C=*:�,
=7�<{S.���"�h@,=��@<'�<gK�=��D=}�<q>n��Z�+cP��/_�M�I�.�%��4����1��F�<	��BN�C=�l�=պ:=��<����c3�Y�B=���욈��n�<&Hd=Q�����9�{���B�*����=���<����K9x���_=40��]�=RN�<��U=�p$=����z�u��/ͻ�cv=�̀=��B=jӦ��Ԋ���<Շ;⻅=I�:=�	z<����5�=����V�=�d=d 1��IG=�Z��e��F�=�|��V�ѼQ�=g���a<�"��FU��e���=���;]~��L��3߃��}Q���=
'�>o+=�Fj�^��j���k����;<��5��$�<�L�1�^=&re;>=-y���u=ZH@��--���=9=���;�K���=Nv9=KJi������;�z=��ͻ��O<�8�=���=�Ӎ�=�=�$�3*T=�)M=����L���ڵ���=���<�F�(��5�@����=�?ϻ��Q=F*���]3<�/;�m=�^������y4�=����]�Y=��=��==�尿�\Z=����;=1����鼟���-�<��=�eE��\�b귽yӇ���=�����tS=��ѩ=�:�=El�=��=0Nd�P���t(��2�h�������=�<o���v:��=�
���U<���C-���<�<�U�����7�	����<�d��l&⼣�j<Q��;�/�<<�=��b=~�3;�o��e���3���l�=W=#�n��J�=v S�o�0��J#�0��v,<hϻV2���P��Ʊ�<'Rغ�%ݼI�<8��=)�m�q\N;��I=-f���y�'���={ջ$]�<�-���e�<�����WR<���l�<��W=@8��iK�d�V=�G`=�+=в��I�;CIS<F�v=`��F�=�-d�<9���?�V�L=��<8מ�A���	��h��<SW�<!��g�r=�n<�L-<�߮<'�<[
d=A�g=�����V8��ٓ=Ҳ�;�������=0 E���r=�JR�߫�;�=�Ǆ�Tɐ=�6m<<�z�τ=�ǜ=U���K	A<��G�� ����#=a���Ѻ���1����8=�Ҙ��(=d�=h�]=�I_�>�^<�(H=�Cۼ�.�<�s.=�h=�̈́�mm�<����6�RG�w�';Ħ�<�W=�Ƽ�8��-����J�=)1S=i��<U-��YP�;����O9���3	�:9�V=,�<��g<2�=�ׅ=2W<���=��=֏����=���+Kt<�z+��Ba�z�������s��������ZB�=H��3�%������=�o�ng���ܾ=�3I�qS ����b���X����=�w2��7���=�x<���3���VK��
�=�\8��\=��2�Tτ��M:������,�3H*�|�=j��<E
�<�R�=W��=���-����Q��붽'Z=��';�t��`�<N+�����a�K�=c��<	_=Q�=<%]�+7=�L
=�n����<f<2�W����^U�� �.=@�5=���=Mh�:[���&T=�0���L<���<�Z���87=~�;Ԏ���p��7�f�h=��é���ܼ����V������/0�hM�=4��<�5���n�3��=��U=��r=DL1;�/߼b�9��=��'�ռ)Xu�%�|�+�|	�����St��B4��s�<��=;�8���k�ky<��)�GC�_�z<�=$&a=p3]�М=�<���v���CR=�Au=����?��=��<*[=]�P<(�v=��L�yy���1.=s�d=<�%=Bh	<���4=j]��xW���;��Žs�=
h��?�==S4׼����R����X=6eN=��B<OF|�(\=/�Ͻ��<��o=��Q=P�X�j�p=�Fo�3��<��8=�
��G��޺�{=f���x���2=���< �:�T=F��;�[�HAw<+x���(z��_=��V�&���^h=���=��=h%�<.����+H=��.=f�˼�E�=+�������&�ƺ\=h��;�ڒ���˼z/�=���� Yʹmn<^{�
�j3=�d�<�*�(.���b��џ�<�[����'�6�KAW��K�%4��E)=CzE���<ۤ�<Z��=�\%=z�L�]�L��u���k4���<T˄=�Z�t�7�g�=�9����%�xr�=�S ;@���3꙽ʸ=.��<�:�����<i)ϼV�T�����;
�=�� ���=J�0=�޻-N�'C=)�<�ꏽt�=�!����=hڌ��`��k6��:5̒�����;|�����<��:h'=+<��м�jI=+�D=\��=k�<!Mp=!a��%��U�zᙼ��⼏���<�nQ�sN��Ͻ������/=J7O���<*e�U�Ի��z=�=8w��0T�=��=�HI��	=�Q��B*'=����ʯ�Vy���}���F=][c=,�N=�C�=���6�r=!N���R��L�c�����&�A�x}C<�IX=7%B=� ��Ȕ�b>�=���K�<B�J=�����=�C�M�ݼcZ�n�½�Dݼ��<}
}�_L��2w��X�=� ��ڇ=z�{��8=o��S�W�9=M�B��;n��=e�S��2g��f��<�O=,=p�T�����p�4�C= ���4G�=1��pZ��<s�%=�r=ހ���"�=܊�=aϤ=�?�<]/�</&���օ��ύ=�
=,��<J�=
��j=U9=5��=�E�g�n��#6=?�<���=зY�~zu��}���!,��bC�o��9�{�<�-�;�G=�{�<h��ǋ� �=j��<8�]��~�����QE=�!��;B|�=��=���� ��=�]��
��@B�<d�=6�&��L����ܼsVg=�����3=��:=�<�1X��8�Q%.=W��<b�޼�/r����<~�ͣ�6ҷ=�ZX=�o	=><3=���}�<:m{=��<39�=�jS���G�!?K���<f)N=���G��;0���4ټ����\-=��ʲ<Z�ڼa�;�n=.E�<$6�=��ܼ,p*=](Ƽ��=Aͼ m�`�8;��ּ��<K�=��f<)��=�K����N����㿤=�"�=�a�;Yܑ=�{��YW�<H�Dd�=f�8:�s�<�RѼ��@�2���i����<��_=OO/=x��= ��=��=�_�<խZ<�S��^�=�<��`
<BW�<h=�]4=���<ԏ�<
�¾�<,�d�.�W=��%=]V?<�C�=\0ƽ�`�OK
�q�2=g�1=���<���ϑ=�<=G�W�3�=4KA=��=�^�=��r<��w=VMc���=��;=�u�=jY���=_�<=�~��xݏ���<�ׂ=���ꨫ;�a���v=��<��<0D�]��:W�˼���&�P�<�4<���PXo=��v=f�=�[V��������*H
�9Z��$�<��M=]��`�M=6�=�З=<Ұ<߹��V �=�(O=�O�<��=s���QU��;:=NX=��*��l}9�C�/g���==�Ua��%I=�F ����$ �4~n���=Q��$i=#}�;��A<bӶ<��P=.We�W�=��=.փ=�և�fP�^�3;�t�=�����Z^=�Y���}������L�����)�������:�=����o�J<t�x�X���k&	�hA�=�q�=K=��N�ݵ{�!SK<�I��j	�����=���=Y�	�ۉ=~K=K�u��H�=&7�;��\�(~.=�	��w�=�0=0�\<��<�~%��cn�u�<�;���k�]�f=a_���n`=�d]��.==��e=��/�Cب��'�="��6	=eC1=�\}��J�2�7����<��=FX���t2���;�B}�
ӫ���=���=s�����t���IdP�B���\i=��=�ގ����:B�<��!;��<�##��3�<Q"=�=`��<���U�K=b��=�G(������#=��F=�a[=%|�<�n󼓽������jw<�'�1�d��^�<�ߘ=iZ;:���\
�;7�=�n�<��=핼��<�� =imx=Y;ڼ	3�=4e���=���#d�g=���	��9�x=�4[��I=��Լ���ɰ�SL��e*s=��:��=�>���'�(�=����e�uD���N��޴<�N=�@���w�<���:��2=�@��D`��b:t�b=O��=>�1=EN��%"��h�澯=�0�L�=~�G��0�<�@<�ʼ. $�+���;U�=D0�;K���3�y=Z�j�=^&��m��<o���AE�Ѣ4=�9ڈ=l��=(���T�#�X��n<�u�<�����D=�}�;bW<2=��(�J=Ā����k<JR���_�����<2!����޼'/���m�v唽k��@�M��޲�1�Y�}曼\.	��v=$\�=M)��W�7�'^�:�MR=ڥ��S3�<갃=�k�=��м�Y�{�D=�bW�QE�=�Ф=RzU=	��r�ټ����g=}�<{>��z#��͓��)���e�A��=\�<���y��R�U��=1Q]=�V=Ӫ(=�8=���=mlN��	����3�=��k��b��W㏼z銽��M=#u!�����#
z=C��=���=�z=�8�<�L���97==��ՐX=��\�V%�=3A=��<�I��ז�=�͛�I�.���=���<�K<CǓ��X=�E= ��=E��z�]+;��k�\&V����t�=�ۦ=�I6��:��l�֫=rr���C������t۵��$���8E��aۼ|�=�C�<�\������ ��2�����*G=�[�<IUy�r
?=��N�����~뇽k6q��TL���%�>�y<[��������;�濽�y����	=
3��ן�==�(e�؂P=I���sa=՜�<q]p:�>=��=S=�I�������<i�]=�܃��aO=��=А�.�;��������׫�=�Ў=��ؽ��b=X����+M�D�<����az�@���d�K�=<�W����b=�^<=�ֻWP?�C݉� ���Z���$k�R$��'����{�� =�=p����<]=���G=��z:t��b�D=h�-=y3'<�jA�i�l�Ym<�/c=�&��@�=s�'=k\�;�C��ެd�FP�<#B��+
=��5�oh��.��=���=-����$��Q:�V���^=�\}��^K��>�dD�<�	v�0�7����nl��?B��X�<�����ҽ��-=о~�B�v<i��<X�E=M����\=װ=�N�e;⼁@�<S���'=S���!�����<�ީ��>�$�x=� ^��/j��$=wW��|�=�k�<0^w��P�%��<��K�|{�=k�q��D<c*=G�"=\&=f��a*�<�HI�qu�bZ;�z<�&� A���Q=��<�Z�ہ#=0���"�T���j=<�u��I�=��<ʗ=yY�=��<�����`<�=Ē�<�-|�V�=�g=0��=�W��zE�=c�����h�<X'����o=yE���)=�R;���o��I��� ���a;�`��i�< ���YL����A=.n^��.�=U؅�A�<�2�=US�<v/g=z=*�O��o��}�'=3����!�<Ǒ =���5N��d=m�#�愮;��ԝ;�м�] ����<�'L=� =<;.���<*�����<%��=CȄ��@=+7�<ax����5<��<<��o��=��=�ӻ�����[t<	"=���<�Ug��#=C��;�uK���^]��9��/�=K-�;�k�<�*�K�L;�d���n��:NǼ̠�0DN=�G�BG<d�{��c�<k�v�)ȇ<�N�&����<�����I�=֛=d8ὢ�H��6���-<ά^��Xf�gPV�*�98�����<����8�=捽 HU�`����Y=��O=�ˏ=�w	��,��Ogc�V��=�i�<�y�&)�{=a�
����.
=|�<B�|��'=����Ry�w}�<�ّ�7�����#<�@=n�=��b�����^%���8k=�%t=�}N<[tT<¯�=Mۼ���<��U=|ǁ��5o=޺w=�$=a�C�t�g+n=W ��6.B�N�<?sP��/�=s!'<�-���=^�=<T=z��������#��E-��=�*(=N�^=	F���)1���ua��l��
=�����{.��l�0�ļ �&\��hg=15�=�ㅽp]���	��+<e��B����"=�7'���<j��<�PƽWr"�S"$=���}=v�q=�G)����=�R��Q0=�^����q��<��=Np����=��=�O������ ��=�"���,<'�z=9*�=e�\=<�P�_wB=�q|���o��V�<O1��'��qUR=���=���˼��m��`'�n�ż�e��C
6�j>��ς��������S���@X�=NR��@��W�T;�~��|4���g2��o�=.�w�x�?= �0�,����<��0�=̕{��4:�t =�R���L߼�����=E�;�Y�=ٗ>�ƴv��4��2�lj�VV=h�&�����97�a	�:ap�=eM=K��x��T��<^Ax�D�5=᩼X9i=>A��PS=j����Ն��ݼP�t=E�<�vԩ=��6=o+=�C=�1]�ɋ�=�e�<���ۻ����w;�q=H�ڼ�nl�������2������x���=��e�|���P ����;fy=�X|{=��k�Vl��y+=f>C�Rl����a=���=�l�;�9�u�=�3�����=��Ӗ�;vzu�z`��v=�����@����Tؚ�ATV�۩�=�hB=:�A=
1߼���=� <����6��'=���=*�K�S�a=-�=u�/��6g=b�<��N<?2t���.�w�K���m����<Cfn��'�=�D=f�G=�=m_Ҽ��a<$�Q=���;D0�<��=c�f=��`=1�=:e<=��X<b�=E�x��Q<������W��7=ߤ�<��;ܰ� 3=��=�.�=Z�ϻ�8��N�r=g�[�]�4=��t=�!��6�[M��y|�]QT=���=���< �:;LK��|��p���|=����H�=�e8<��4��t=�+��By���fH�q�ۈ�;�#=�Q��b�$��.���@���5=G�$<�ԝ�ڻ��~=,1s=�4s=�3=8Ws�<�<P�g�d��ω���Y����< ��=�
f=��M<���2_J�Q�@����k#=�~̼2K�<e���ˡ������O�<(j���I;AL�<~���1=��=HX&�_�6��Z=�Q_=�"=�?K=3��=�9���M<��+��j��u�=��<w��=�9g��Z�=Wߨ�¼F=ϫ�=y�y��1���<ǲ�9��=- �=��j=�a	=�Dg��B<C����<UkN�g�x�	k_<�h=Ƞ�=�μ�2l�W��<v�F=\�g� `=��'y=��=��=�!b=Rs=P�<�<G��z<!��P�<�휽��� ���/}=Kt�<,8��Ț��m���5O=`����~�<:==3/=�X�z;�d�=�*���3=Ơ���p��x����K=br�c�T�ȥ`=h�T�2]����(�p˺��Q��͖;�bm=�7=��O;�\��;_T=21X�7�
��W��!��)B�@��=����1:=���=n>ʼ�Hm�����F�<��=c)�=�>Ѽ��;%d��
��=pݘ<����C=���<�?v��z�<�,U����Ɇ��Ê���<�&�']4��%�<��)����<�2��񋐼�ܠ=��<��=A��Xn.���-y����+�h���	;�L��[�<j��w�Y;"�<���=���=�S�=8&	<әڻA����Küj�z=��ļ��<�[��;t���3=�=��T�ۡ1=Ձ��\��l�4�?�<���Ѐ �ۀ<��d=��m=n�]�]�L�,����>����������*��（�D8��zƘ����<\�V;N=x��=�+����<����\�S={�!=����oy��><��ϼ=�{�<��=��z��<Ѕ����������3r����4�|�+�&/<a��:k�9��<�)��|����X<p<�ݒ=	�l��=90��4<u�e=QӼW��<�T���->��Y�����Z�9K=c���(�m;mӔ�K<I=?��z^<ez�Z|�<��<�ݻ��G=�<!��y�k�<,Ho��.ɼ�n���q����=�=�b���=7����Ӷ<�V=z��=��1=j4�<��"�T����k�<����s:�=9�<�n�=3E�=_}8=���${��b����۽���/=���;I�=�������>��ütr�9��s���� =�^Q��T)�Vt��[��[�=���>'�=����<&"=�c���"5=�C<��-���U��f{�f[=��W=�p1=��=�a4=�=�ug��8��:��=��N<0��=��;'�w�@�W=�I=E;�=Y��<&����2�']v=]m���<�d�;~ ����;�Ch�N�J�}�[=VP��M�ɼ���=�Oj��{*��^�;_���?��v%�=A$��=Fz��14���	�=-�@=)P ��.%��v�<�c����;nѼ�Y��]=QW�s�t���e=�2�<�����9=�;�=g�<��%��Eؼ�@=70=NCe��j��/�=Lk=� �=d�Z;�uX�d���`�=(�k�=p<7-��T�l�5������=��^�����'V@�f|b<3*T;�p<����KW~=��I���<�j���<��<��=K޼�����=�O%��eS�e
M=�H���<�љ=�����^=$������<�=##I= q�X���t�4=����8ͼ�+R�"��ihN=({�<M1;=5Q�;�f*���;ܣ�<��<�ȡ=ޑ��2+�;wZ��{��O7����� ъ=Ǎs:Z�(=���J����z�Q:ݼ�i�=�Ҡ<����
;�m�=�m�=�/���~�:�9�=�|u��M<�}��[�����=2t>�DΨ�&��<ϼ�=��m�td�}���Ng��
@=���;�
f�����dv=��=��2�������<ǃ�=�ª=��=07k=ƙ <�MX��Xa=�ȶ<h7h=�)����d9\��������'¼�Qs�O����异E={D�=O䵽S�<�1r<��=����=%V<�W�������bR���W<�[�<�0u;���� p6�렙=�C=�.����j��C���=|q ��̓=HԚ;a��<�O �L��=|[�<��5�X��6�N=� =N�F��i�:�>+�v9�;ۼ��i=Lg����<Z�]��'=ٿ=�B@=$��=S�=�%P=W޼�%���=�/;�鰘� �Q=����jH= gB<�Y=2���6F=̔x=�R'�T=]�9���p��?Y�#�0<ob��;d�<�����Z=�A<0�����<�̥=���{N<,��=P����=I> ��u�����=#s�Ӊ�<�Vt=��Y��]?<O�༳�c�`�m�玞=̫�<j/=����a�[=�惽t�w�.K= du�N��Zn�����<��=~i����*���R=��»}?��Ŏ=��=��x���<��Y=�֞=ۼC=��g����=I�=kL �돐��fW=#�#�Լ7�����؂=�,q����aI��IH=�e��d=�d�=��=�}�<�����"�=���>I��4��c+���e�����˥��#;l��<�eW=�q}<��<��(=e�<��x�*��샽)#�=]T���'�	 U�zʻC�<7�>S�l���j{�i��=g?�����=R��<��Z����M =��G=��:x`=A�=観����<{Ԋ�Zş=�Kr�ȋ�=�����=��V�=�����=^�<'�H���X=<���.��{����=/�����S��<9�=2>y�t��=,d߼�w���=���<4^=P���<��4� �=��ټ�Q�����=��<ə_�����쒼.	������h�<<EC�=k����)=ʪ:᮲�����k�S�_�<ht<�:�<�&�=�d��i��iqw=�w�;(
�:#����'���Ub<D+�Ku�����<�/=��t=��=� ���#����<縟�*J=���=J�	����=�|X����;]b�<��"����=�+�������;�v�����=�\~�{���
$��y=d�4�0�ڼ��*=`f��֎�<��
=����;�O�����G���y��Ά<�+
=��[�Ё?���<�9�=
Y7����B>�FG�;�+
=|�8�e�U���5|<��؊m�����˲��z=��.�&
<.K==�����7���P=w��&<��B�~ ��Xf���yj��
=��g<7 �=��;	�;sŌ�l]N=[c��F�+=����Iw=�L<�<<�3b��u��ۑ��& =q`=��v=~��;��=,�뺠�<U0�x�=k�N�4�k��~�=n�<~o�;ů7���?���*� �]=�|Z<�B=��<6�:1E�;G��U@=�Y��9n�<�D<;�=���<��f=�p;�K�=zB�=�+����3�=#�_��P�<�:�;��1��CZ����=�e�=���<��S<cܲ�	Ŋ�N\<;'�=3b�=��м7c�<ǖY���d�ￂ=DX<�|�%D��A$=���<)�=gk���H<4E=/�H��B=��2=$�=j`v=��=r�!<N{q=a�< ����9`=�3r����c����S=�|��o3�c�p�����S=?匽�cY=u�7=R��=��i=�	�R�=<����P����<{S�I���7Z�՛�;g�C���
�EM�=��<�S��@d=��<<��c�����@7�ی��96��N�F=��=�&Ҽ��<eol;���~T���S�<��r�Ue�=�ث=/&��!n�=[A�¢�<��]��	a=P5�<�U�j7�<���<95༤o�;���� �v=b�<���=C�
�y�<��a���"=?GZ��KH�DN�=~ܢ=Z-{=���@�=�T?���s=�}���	l��1\�ȗs���~�SkC�eー�l=���<���������\���u=�t(�W}=��=8C�=�{B=�l�<ٷ=��=���cs��t�=֘��x��<�oѼ�Si��ԧ=�5�;M������<Fy�<��)��W�=L����8/��HQ=t��x ��(���H8=H�����C=��
�<�[E=)�7=�d�<c�d=���eܟ=mC��g 5=�s2=�߻D�=l�J���=��<��ռP	9�=N2=��s����`�;���=���;��<��Q=bỉpQ�h�&=?��� </���>���=5����u�;h�������+�3��3��\8<�v7=;��yd�;��=<��=�{�DO���;��$�@����� μJx�<��}�0=蓠=�0�o��<)2׼��w��H���=Z���s˼B�O=> ���K��v�=��=t������<~�}<蟋�2�U�GH^=�M�;����8�R�<p<	ܒ�o[�N��=�!=��<��Z=��E=^�<�E�=d��Es(=�M<˿�=��Z=>�Z=ߩO�l���ED+��=ۼ(��=XsC�KE=���=B>M���=��2=�\=~��<
�ܺX={��ǧ�����Jr�_���0
�]!n�w���k�=ڐ�<�Ȑ=��B��,�=���<O!�=��<���=,�3�������w=}��=�c�=�y��eܧ�N),=@N2=C��=Xg���6�=g��=&�<[� =���=�F�� �c=��<�GP�����x��I �ap�<.��m�0<)^ӽ��V;4k+=D\J=��e��NK=��:�K���o��^$r�r�ܻ\Z�<���(mp�iܫ�yEܺ܁�qϓ=����B���=�+��ּw�.=B�D���=��=1-C�d��=�{��������$=bi���w�x�=���<���9Ę�7Xh=x�=���<�N�'�/��_��S�=��N�^/=�Hq�!5==_)=���<�)=��=�zۼmii=�-�g����==Q��=�k���R��b�Q��^7=Z�%=u�E=+{���z��l�<��!��=�H��^���=��]���=���=%};X�@=�����=�<�����ƽ�a��}T=s�˼~?6���<�ת<�g�^��!k<;Me�:��<$=~�Q=�H�"*��������>��J���l�<|
0<|�7=���=��C��_��p��\z�=1����A��
X=A�=���=6&�l*�;/��=L׆=��n=�o���B=�XE��=g8��X�ּ�A�=˰v=9ļa��<V�<`�Mz��]=���<�j�<��w��늽�g�=�͍�x�=Ɓ�=
q���<���=�I�!C�����\ռ]�<����1ꏼ=oY�E�a���	�Tɳ=~Ӽl�̼[���S�=(��=cD���X;��\=Ϝ�=�y��2��B�=��$��
=�{�=N�U�T�ļ�s���,=M��=��G�~�`�̀���lj=�M=�YT<6Z=�Y����U�9��=h����m�MJ��Q?Y��˹��(=?��\T�=r����_�2�z=���=�`�Rb�<�Ku��ݓ��|K�E��=�ʆ��GQ�岓=j��<��<t��<L���{T=�;=�J;=}�;&���t�<aò=Y~=շ�t	���c�=�='�k=�����K=�3�=���q��=�9H�������� JZ�Nk�<���:��x�J���m�%��2�Y=*8�����z�=�J[=��g�{��<{ۻ0�μ�L��=b�1=��m=ʡ�<{M]��.�;u��<��޼@�E��8���n��9�=�K��O��=���<�����؁���p��u=K�G=2��[NR=���ɮ��	[=��=�(=AM-<u2�=>Vz=�m�=`�=��(=�/���h����� �����<�s��4�<�n�=�Z��v�;��<c���%����(�<���<Dk=��y�M����C<�����gL�����׭�����=���<��v=AS:=+Z��D�j=UZ��c��<�6D�D���J�<ʍ=]\=�U�&��=�.򼡠T=bt=��w=_�<?C<d�.=򚐻�M
��v=�Y�#@ټ�%����n�W��;���=�'�=}�Y;��(=qЅ<�Be=)�=��
=��<he/=���OS��$*=��w=�qr=��<���=�+=+�=�^E��駽�o]:��I=����Ɔ�_�ㅽ:!�X���<+�<�7n=��{<�[G=4�@�ӫ��r��<���0塚y+�=���j�<Ax=��^=�<a=�>=c�<�.=eD/���N��.�=���24�=�O��=��&p���P{<�{�=�=�q8�e��i��=��<�˩<5+X:'Y>=GR4��K<��,��L<��懽MA�<zv6��F;=^���caW�墓=��2�Zup=?wl=��'<h
=
�h=x�`=���=Y�6=�ûӻ�=�==��5=/���b��� �3=�u�:�1��#������#�;	��~=Q�������=C�<8[�=8��RC<|�<��?=�ե���VͼE������?=��8-Z0=��<�=��?=GP��䔗=H+�<Y�=^�d=J0�<�~��S��=/'�ޟ4=��#=&6�;)=���8=Q'f:��=�Y�<c��s��=�@�{������Gb��/����3M=��0=�"��ާ{��`�<�W��0�c���F��cO�
���G�;~�=󪩼��):��}Xa���M=@��8�I���g=��Z=-N��yϪ��Ų=A��<H_�=J�c���=�|�;F"<*@N<�(#=m�\��3>���/�!�H=G�7={(+<:�<�y=Zk~<#�5=��<��E=S���b�=��9=2|�=�m<�OE�K�9��=�˝;K����P�V�S=�+���o=�t��̜K��05=뺅�����ƊF=�S�b�ɽo�O=���=KvR=ܗ�=Th= ���OM�m�����c��pn���5=��=�^�=��4<��`=M����Ɯ:��=�OV��pL���<��=��<=.�W�9� <��`=�]��y���$�;�:..��=���Ϗ=����י=���=�����f���<��O<׊��/��<$�N=n�Ҽ�s��=�1���l�=��ݼZ�o�#���M�<�k��nג=:�@�$�K=�-]��7`�+����CC�]�_���P��0	<��/���L;Cɏ��iU=���:�I�<��=�*=mL���
=D�T=��n��=�5�=.�E���=�s;�t���\�<�U���Zʼpz=_S�<+��<�m;����O�g�ּt�����ۼ���;$w<E�μ��d��j��k@�=n��R6=6�+��u�=*}f��J=��d�qQ��t�F�`��&j�=�5=�km=�R�=�UL=^^R�����c�<�?�=�@�=8n=�=�6�<�=q�������wN�==�;5=�G0�I#׻WB��r+;�[���=�<ߴ��r =.g���ļ�B�==*��ڥ= Y�<0~I=џ�Wʙ=JZ<�д�z��<b?üN\�=hX���w�����v���y<=T��<G�_��Ġ�s }<ј�<��<���WѼ�҆=�e=LlE=xU2=T�<V%��r,=�h����g=\�*<i�l=���G����;�����/Y����������<����in���2=��=�z}�Ȗ�=���;��=7ʛ�D�}::�=yw#=|YY��X�=���n��8&=��z��������<�<�;ʖ�<����R�c�D��=$繂�<��üF	��?�=�a⻤�]����1�D�=������6�R)f=j��f�<B �<�R=�ц�A͕���=�=��5�:�]$�x>�*t�<|��2-^=�Ol�l������X��ߊ=�)_�x�N��	!=�q_=�N�=9�w=����m^�=Kh=���Lӻ/��^�=��8�݆�<�	Z�5��ݧW��݁�*�Z=ӧ��\�n=�F��l	8�)]�=R=���S�Y��d�<pZ�=�d<mE=:a9��/[=�T=���=>8�<�x<���H=�S1=��;�߶��ܡ�g2�π<ɗ��}�߼ 鶼�,�=de�����8V�:���⑽s{����;�e�=f�=���[�U���̻n����|=��~=�Ei�H�-�%{ؼ�M�=�X�<���=^1<~�<gI���9n<�Z/=�f��h6=H둼���=�+��~=&
��O =�t�=Wđ�gO�'{=奕��=���"�=m�J<,�����=�9��X��=7=��G����<�R�P�6���7�����Ƅ���<Bn=�]���C =ٮ�#��={��{�=#hV=K6��f�<V�I<\�;V�3��ޚ�(^�=FFH=�	=`���9�<<;����fE��~����=�nɼ=v���t�<�q�6�=pʉ8�;C��f=~)�|g�e�<��<�,�G=���WN0��v�=�Z�=ީ�<����Z�~��])=*�m<�>��_F�=�L����_���~<R�%<�b
�ۄ���:�o�cȃ<~�����p��J�=xS=E�6�㑽����Vv=L_���
=߆��>$c����>��d򪼫���_=s���j��[Iּ�G�=���<pq=�Hs�a�y=L��<,6=�8=�Ո=��o���=C��<ͅ-<����X�=��<�%�=*�a��� �2=�d�V��=������=g̿<�Ɲ�� �<��)Ul=������S=�#�d�4=F�ּMtN�b����U�<���=�=�w8B=��W�M��"� ��U����C��>=5ʼ�^�<���S%�< �W���<o�1=��|��<��<>�]=.�w=����h�0E=�W��?����v�ż%2h=�_�?#�=�+����{$u=B�������̼̼l�5�W=�W|=_���/i <�To��p��yKN=l{=#=É������k�X=�V��`��;ڥT=�>޼�0�<T��=D_;#�=��kZ���ͼ|B`���<8�C���V=ᚅ<V�t=�J�����<���<��<IfN����;����x\��0�	�A3=�=�L=b7;��E={D���/�=
2�<����T7�=�"W=�.g=�
��%�ּ�~: �F=J�(��Jk����<�X�<j����H��==	��m�<L��;4��菽`��;>z�<���<`�;�D�����G�Ȁv=�1=T���K��=�DC=���M#8����<y7���r�R�c���<d	�=e���z�=�Q��pd�=e/=�7i=�ă=(e�=g��;��<�u�=>��=Tż!n�<�:�=��R=M=��:��[b���F="�u~S=�|����<��&������;=��<Cw=A��=�D����<H0(��|=�� �E�R�
���<V��<n W=�����A	�а{=��=��=P7'=��\��/F�S�N��ޅ<�/�u�h��f6=k$�<���TɃ=��A��F���{�{e�=�5z���4���_����<yjѼ-���HOD=�� ����<>�;��o���μ& ��k����<��^;��\��>��漿� �:,��C�g<8.���<Z4=��>;��<-\="�=���:�ߊ=�7��2=>r^<����Bq�=>��:C���<�<�"=���<BjԻ"�;�l;3=���=�=�=ZB��`�<=ى�=�����Y�R�=�?==����¢=�2�=�'ڼ�"��:���e�H�û��+=�.=8aU���x�f�H���@�¼<l�$�k̇���$ .=k=��x������G�=B6��:�9y��<��&=`w�m�m=?�O�;=���<� ����v��M) =��˼�X�=��N��0=����}���!L<�e�<����b��s=k1
9�c~<.��������<��< ~�u�˼�&��������6=��u<��<l�M��a!<�j6=x��Vy=����/�J=G(<Ң�=�LC��S�;�QM=�xv=�[�<�=���N�=�}������z���y:����=6��<�rp=���Z��=��=l=�=(�=�m=�Ҽ�(�<❗���<��&=��<+�f=йO=�\������C�=��8Fz=v�F=��ֺ��ʻ�p=�=ǔ�<�!Ƽ���=�=�_��<�W<b'���N�N;h<C	�<��B�CF�=@5=�<�=�u���<Э?<���p=������1�<�C�=H�J�����\�;gKG=ꖗ=��<Fw�=�=?��:�eN<y�f��I�<�༺�o���R=��v�v]X<���=d(�=q]���E�<V|:��wA=i�i��������S3<�<	�<�����<(�4<	�M��ޅ=ef=�j�;��y����T��<E�==E{�<^-��%䞼Hġ<-օ����<���p@���H=�h=�s�=ߵ�<�˚=X�*=��li�M��<J���j����Ӆ�F���=5�d�lC[=�?#=�ý]�z�$\ż�k=|�����<IL�����=і�=��W�HcX=��:�4=t�M<�n���m�=���;��=�4k�@Us���p���L&q�׮�1 ��g��=�cb=�֛=Ӄ	�-��<ύ��H{O=2[	=�	� q�o՗��Z�=/{%=LO��H���%o=�؟=�.V��(�:���<*`e=�.==L����=�#��9���r)=a�=��X���l��>1<> W=�7�����ʬ���T�<�v�=���'º𭭽zU:=1@��zU=���<�gD��˻<^#�=�ʜ=�9�,�<���<��=v�=Z��\c>=�Wm�oܲ=���=��5�A���f��AJ==Wo���6=7�;<���W��;���(/�<�	; �����|�o�d�����a���ޅ�&�����<�:}=fJ�=$,�<��(�"i�:Lj�<�x�< @�=�H=�32��Z=�`��Z��>�q=���<��{���Ok�Uʃ��Ь��|���䯽0b���R�;�&��f9��=1��]3m=��s��Ӊ���<�V�<h��=�/�<Z��=�;=DՅ=k�ɼeE=3l���Z���=��;Jx�=�����,=tҼ����;���0=J�5=/�ٻ���=O�X=�R]�;�<��=�y�Hgw<
	�<��<㕘�+@�=���xr�=�f_��+ ���̼�|G�v�;8�����p<��`��F��O ��]^=��/_�=����d'ؼ��u=,��;�|��O<S=��½e�=kҼ$�=!!j=D���כ=Z@=e�A��갽��_���f��3�=H
��Bm�䐽<���<5��y�����&=m�ʼ�`G=�É=��)�G��=�ui�[�'=}҈���p�#9=�~��2��L'��9���q��^�=� ��<����=]D��.�=R�;�3���A�=��T=e�=�W=܃�<Ju=�q���P=�1=���]��_G��|Z�� =����@8�<s==�f�<�n��%�ծ�=@8<J)�v�m<�c��>2üm*=^<�2�i���Z3��Z+��2�ҩ= Ĉ=�z#=@S����<���1�E=��0������S;_�4=��Z<ո	=5@�=��;<�s@�E`=&�7=��a=/Q�=z6�����C�!=��,��%|�3�h<%�*�:�@<Ҫ���I	�=�h��=j8\=��;��=r�=}��<jn	=�+�<$Ä����<��=��P���~��=�[ļ�b�<q���g�n�Pa[=�aN=���+.�~pK�э=�8v=`��<���<E�t�m�n��=S�A�`C���J<E�=�Pn=s�1<eR�;��m�ʺ���H�ȯ������
������;kE=G�f� �:�S������\��2Ҧ<�3E;�푼���=��;|�;�S��#�=�/<�:=K�a=����ϼݵ�V9=�<]�ü�;�;_x�:���E���0�<��1��[A�a�;�w�½&㦽Q���4F�����D�<E�K�鱧�)�=G�=�u=k	8=��v�=$p���Z<�9��h=�g.=г���|	=Q��<=.�<DF�<���<ó��C����Ë�KS�ۨ��]8��b�0�v���T���V=/�=���:S��JC=8;p=��&=N���o�m�[��=Q[����+=�z�=}{=�n�<�����8}=(f7��ppi=�T�lic=�S�a�2��]��;�<l�@�㣇�������m�͈�<����mcJ�� c<�H=�����e=½z=&g4����=X�=�ż�\&������=	�.=k��Z�<A�Y��f=��= �<6�����;S��<N��=��*����#���s��2:k}.<ƃ&=1rR��Z�=w
o=�[�<s�<)�=�;	�fͣ:���4�<�$��$��:�=�lR<>��a�:t�=�=j��;W�g=YR�=P�\�����)�"�_����<��ܼ2�;I%u�iѻ<�p<z��6R�<���<�S=ѝ={�=U}4��to���8=����J2�<����>_F=�a���Y�<����"��=.�='9����+0�<G��=W\�;;+�<u�U<�ւ�!��A��dK�ֽ<soS��O���{�B����'=]߽ɪt=* ˽���������պ��i=#�����Q<Q)=R�P;��G�m��^I����<�v�>�H���޼�ȥ�t?�=�O���˽L�\�*^=�=��.��],���G�=F��p4X=�-��:���v�ʼkz�={ө<��ƽ��-=(�==XA�r����|=�y��N�[�z.=�=�g�=웽"ź˱��c!�򄽉q�==q���x2�)�T=}p�=3��=�f��2~�=V"��J�2=�'�/�)�k?�:�2)=�?�:�W<��I;ݻ̼�D�=�6���g�[�b��$��e6�=]#м� �9TX=̗|=6ȼ���=d��=����uz�=���=9�����=�ఽ�9��o����#�ljc��:=��=�M$�\'y=��c=oq='�h=!"<=�=V�e�����,=u�<E��<R��o��+���v�<b&�=�j�<b0A���<�z)�������,� So����A8:=��(��ʇ=˗�L$�=Ԓ�ikT�JZ�=�mI�*e��蔽%�=.Ʀ�W'��ÞԼ��<�\���a<z�ǽϐ=#;�=W�鼯ߍ����<���;�,��Q�<m�=�,=�w��s��Sq<MJ=���<R9=|� =4�=��}<�*j;B��=S���(=G�C����I�P=�V�[.��z�[<�����S�n�Y�O�<�Ձ=�s�����th�R�=�t�=��� <5�;f��<	B<��'<��<�ɽ���<*څ�]�$=�m���}=��=���<В��w�f�)���=J��v��~«�%��<�w<&z����)=�6���=a&P�w�E=���킽\#���4�=�ܪ������=2�=޹5=��׼�؁�����o��gw��٢�NM��x=���[�%�1<��0�����K�_�O� �A�b���=0/٣�w���𤒽������=<�;�sd=/G���>������<�#�=�T��U����;2h�<�A=HX�8Yx�	��=�C�;���[i8=g���#�<��l�9&�=u�O�����k��b����=�;�>����9=���%+=�ς��8=�Z��l�=�V�c@�=�AW<����m<j1�=�����h=��3�=��;C�;��T�rD˼�Y�=}��2g�qd����d$=ri���Ԏ=���G^�?&�=l0y��cI�ɢ<�	=���9�I=PZ���$�:���������=Fa�;)���s*�=�\���^��\;�]:=ɡ<s��������x9Ih�=z�����=~�;_SQ�\,�ґ�=�Ž3�)$�n�j=k�=�<=|=i⠻E�^��Wg=�_�<1�s���}<�z�<��R��\�=�����,�=1�6<kQ�n>Ҽ�L�'=O� =�����B�A���=	 ��e�\=*���0���=N���
��f<�=���\���^%=:yJ=k
�=���b�<&YE=����%+%���C=s%Y��㛻���<RM-��ݼ���<�O������Z0���d��>F=� �=j�=�y��O�=�p|���k=�\p=�����0=>�<����s;X���ъ�� =��r�(�K=P��.=�@r�{,�;��ؽ��}�c��<�M�a㊽�I�$����� =zY�hm=�We=y��F��=�k<<V�𼕩�<$ܦ���&��R=8qU<<�<rhr�:�=�8Z�=�n=mr�=ۣ������=��<L��X�;jһ:���������<%��<�8B=���A��Lݦ=�c������K1;��k�w�]�C�[=���=>��:K���8��e�<�H�=�xh�PH!�x3=�b���<Cˍ�X�{=4�S=u��=L�~=�!K�Q��<Ӄ���x2=Y�U=��~=v�[�wZ��~^���I��f*�z3.��z�='�B=�p�<_Z����#�=O����T�<,��9�����<�'�=�]�}�L<^�{=�9=���<=���<�o=iy�e{u=c�e�/�K9���B;�3=��'=�Z�=�a��=�?=�伖]<]I�=(�<�߹C�_h����V��[=��<�,=��^<x$��$x̼��x<k]7<�u��YO.�x&��<��c`=�G$���W� ��;J��':�(���6b=R��=Q��<a@"�����b������gE=�S�<�"T�:�=�޻<�!h��Tؼ>Y=��Q�Չ=1����g��<��-=�(�;K_��+]�6=�P��A�<��}:��n��1����d=�^�;�ٞ=��5���
:x�����<:V�=nM�<	�;�����c� ѵ=���6�1��%�����)�=tr0�H�I��-�=�=�ٻ�Z�:ũ�=sϖ<+=������\M=�= <�jd={�;�m�=��c����=��I=���H�%��qb�ɫ=n�=��F�|+	���M=��= �=2���!=�B��F�Q=T	��$=� ���C�=7p�=~�i����wˏ=v��3�;��=�V:=�Vq=)Q�=A��=B�����h����:�`K=#,g�mL���YW=����ھ�<�Ύ�oY<!q�< t�g�<y��X�;IB�<�ǹ<���<m�;�B����a���|��a#=�Z<���<�A=�#�<�;U=-3i=V�<HPH�Ԛp��#6�"&<Q�=9R�<!���w��<bO"�Ew=�|��uD=��=��W=kG=��=ѷ�<��3=G�Nu����q?t=�h=ݱ�<͔+=Fk��k�������UV=�������=��a=(E=������<S?¼����&$ ��x��ږ�\�;YM�
�S�<��P=���<<����=��=g�9��q�<��)=�d��z 	���v=m�4��ּ��m=Q�=^��:���;T"���R-=]��;��e���=)[����=�_��b�>�{�6�,�˽:t��Aַ=G�Ԓ�����;�}�<A缱�<=B����u=0 �=���<�sR;�b�=���=��<�cy�2��=`�F���e��;���o�:iԼ�Y]�V�=�=���~����˻���yF�=S뛽���,g;U.���/�ް$=$ |=׍k=� �=v==������ѺH@���;���(i�%��i��=��.����y�:=�$�.�;�g�< ���D�<J-[��Bݼ��U=�m"��G���l=;�p=%v�=��<����V[[�VMu=t��<�G=k��<�dV�v��1zY=��9�W	=e���A�@�q�9�e��:,,W���������m��C��$���[�=A�m=,�=oɗ��hI=ח���E�r�_=��c=@�=�e!=m���(s<����������Y6�<�W<k�<-�.�}��=T�N��F�)��$�:�<���<�,�˪��FZ�=�%��7�F����=�f��i�<L�+�w �=�dS�v�=J�[<�2������R�6����j�i�G���f��O��RG=��6=�=0�˼W��<܅U=���H��X)-=�=@�����=����Z�=�C@�Z{��H�=����K�=̄�V�/=���=��h<�gu���W�>��=J�o����D��� <�)L��Q��K�<t>���eT=
̀=��W����<�:<ٲ;�6���=��S=a{�<��<��{���'������?��҉���=_��=��=(Ƌ�Y=�$5�W�X==9��'� =���=/�q�t�#�'�6=Gs�=pf�<�ai�Oԗ��ٞ=��м�B�Ԕ�<w U�+�d<_9G=���<cJ1��<=��=:�=�'����  P�<q��Og=�~�=��=E��<Bj<e�R�{�_�2;��tk��ܻ���i<�)�<�u��<����j<��a=�p��v=
�׺��o����<�.�<y��Y1`=Q/�Σ�����=�
ռJY�=^	,��{��B(����[=q�y�X�W��N�ǄV�)�=�W�=�ż(-�"[=�(S��/鼁A����=?�)<�5j�?׏=�̽��3="s=�=��{<֤���S�g1='dO=��2;��N=��<Mq��j�˼	���P�=;x!��ƀ�����3n�����A�=s���vH=����zB�C ��g:��ŕ<��=���di��-A�;�Ek=D�w=)�=M�3=JG(��Z
=��g=�y���C�=�=�"6��\=�<=��/��dF�^Z;�:�=�T;�L�{R<���h��H	�<�eX=�w����Ѭν�G=��B<��H=M�����=��=�=�=�k�= �C���D=X���!�o�S	�����w�򼰩�<��><���4ر=Eig=����V�us=gy=�S^���ڏ̼*�Y=.1�� ��m�V��mB�P�=k�V���C�&
��Y'�{�4=���=���
k:=�G��S�n=�	��Kw��2��Fi��Zb��z���
{<��=�Z�<��D�gAe��B
�?n��JQ�;�����x�<h:��"=��7���;���:��n��@C?�R�=xV��������>P�=80̽:������g��|�=,M4=�-�(��'�;ў`=	;� ��<���<�c.=Eg=^��=����a�<�o=��޻������<pt1=y̲�;����1=���dL���/����=�=G���5�=�m���T:Ld���=�yN�?�x=W���6�<����ż����9:���5��l��<@o��	=1�����2�<8�D�	���Ѿ�P��<�0=�"\; N����=Z�=�@b�Ez�=�ӻ��l=�V<'��=��:<j<�k��'���f=�g���c��._<��}=�#�<U�=QpH��]����r:�j=�;�%@=(X�S3���0=Q�E�yc=�K�?��<�������=����V��<>G�<|���
��9''=�M���2�!�*=���;�����%�y%=���=�Uh��`���/żAGl��џ��s�<�<�o_�?ʈ�(�3���=^E�e=]��������<W��n=f捽̜ =)�,=� �9�7=x�T�\�V��ګ�L���r��i�F=B-R=c�"�.�D�"\��t�Y�<�0=h5���[�=y����U�=�
��'3���A,��wż�=2R�<�l,�Y���w��Řz=�4��bg��]����<�缞��=#��<�<=[ݪ=eH�ʤҼ�����C��n!<hm<���2��=c=��ѻ�����6�=G8�<�%k����=�G�G=2="���j��1|�k=K[�=n�0= �=�7=�� ;�X[=��޼W:6��������=G.<r0�&=�g�������s;P[C=qu�P���4�ɻ���=	=3<��i���=��=~ذ=�$���=��T=rA�<G��<�!�t�c�h����=c���`�:UC=���<�З�а���9=�D#�}�X=���<uq�<��\=v8<�ջгC�4�M=��F����<G��>-
��rm=����E�R,��Wv=�B-�����L=v_M=�G�<�h�=� =�|m<��=F�u�Սw�K�w�"������<�N�=1���f�]=�BP<iQ�=s��=�y*=Փ?=ڱE=�5�`�=�Jl.��Չ��_!�0�⺗�{=��"��b=�ғk=|G|����=U�|�F輜�H=�g��`?����<z@!�.O=giܼb̻�E=���,�@=@�(=J�=c{=���<�kr=�lO��p�;݀��N�=?z�<~S����g=$�<����𨸼s���]׺�H���~=h�<T�z��Y��m�o=ÄS���=�ν�,!�0�=0L���<7鐽�[�=���}Z�=�zj<JO<�fg=�p��	\�;'��=�Rü�,G<��:=͐�=m�i��[=&����_6=b�@=W�<U�O=��6i��=0L=�y�<���f�N=�	'=`�-=�,W=� Q�h^�=cL=?��]�5=��u=��W=�M�=(�;1N�<1�=��<�@6<P��=Y�_=��N���=]	��I���;=
�<�b�=|(���=�<	=s=p���Y���
=�d��۽�\]=&њ��i�=Ľ�=_^=Y��]�I�\�=y�=�8�<<�R�b.!�bKW=*�j�B�<]��=�=@�１uh=��=ߞϻ,=8f�� ד��������q�8=��A㱼$(�=���=Y2x���i����l�<V�R=i\|=կ�;��=��8=��Z�A�K=�5O�M$=>C����?<*�<�q�;:����=(OT=�HL��9d���t�A5I���=j����򺽰�f���=!�_�N2�<3�T���3=��=�w �x��;y9�<�+'�Q��=�p^=5��<?v<w^�<����g֪���=jg����1=�t_�%V�=�&�Q�=7�o��Y;:�~��T��7�Cӟ��є�5Y��Ȱv=�py=��=�l�=��=�ڸ<��R<vS�"�G�DԆ=�,?��^;{-�:
2��7���=�2��u=��F���J=�[:o��=Kp񼟂��^�z���ջ�|�%¼ŋϼ��FD=*P���2=;��=�>�==�<��
<�"=���w�=ٟZ=I:-=���;ł�<�B�<���q+��rҎ�9�=έ�������ē=i=�<֙,="@N=5|m��b�=qQ��7��������H<'M,=�, �sx���=D�=�4���r��k"�ə=[5��y�=hN=˥;99M=�c7=�*e=�~z��ڝ<���<���=��p=����Q����ی=�L���eJ��2�=�Ƽ<��=:Q��������<��=ܫo=�=M��=�w��Y=�ͨ<�<�L�:�ٔ=����
;���<��=��=�uC=�-�=e�N��=J�=��=�R����<�:�=�H��t�:��9D=��i=qq��I���Q6�=Zk���=�[3�ew�0�=�`�uv.��5�AX=k/=���g=4'�@������}.'�Z�L<�@G�ƀ���r���OD����<��<�|&=�>�?��=���<~�|="d=�'�=f_�����;^P��>��S#�<U��=�z5���i���9��Sh���=���;t'N=r=�� ���0��<4'/<<j�;c֫=�?=I�=Λ�=�ǟ�6��<��S����.�V;�о�mv�f�¼"z����p=ƈ+�/�=�Ԩ��'p��4��<l=���=1���A<=,�'��<�޼zu<t���K;�ܦ<^'�=!$=폻L����9=���;b۞=��=�k�e���=hl�;L��<K��J���+p���\�<?]4=`�=,z�s�=���=\ۖ<'�J=��:�皓=��4��k=������ۯ1=_=ƙ=�3+=��;��#<s�l��M7��H0�
{�=R=f�h�Rt<�O�<�0��6s� YB=���MpK�+n�<sAx�-�<����v�=y���W�=���:I���A�0�P=g�
��`��tҥ;�Ý=���<_�.��9=I-=�)����V=\�[=*S'�a����='s�="L=/��6=��_�<���=�+�='p�=�e����U=n�=��ʻ��̼ܰ<��x=}0�=H��=�J�j�E��ۅ���Ӽ�ʤ��M�=:��=��=���<��<Y什�N=P�I�F=�����<���yN@=ߴ�<b�U=�mM=���<SҼ빽�0=��:�g�
�B��<w�^<��<����e�Ǻʂ�=@yB<�V<�}o��;,=d6*�8"Q<���9�eI=@/�=,6�������)���i�=�_	=�z���Ѥ��'<�4�<�SD�
��<��=8�=3
i�@+]=��,�������R��=.V�=��.���[�=�ϭ=
y�i1�=C(�<U��7��<�]�=|ba�Uk=G]�D��<��<^^V�@�e=4>|�" �=�u��"��<�3뻂��<?
w<_.���#����=���=��[��dk<�ϱ��t�y����暮< ��=hj�<�E����=��+;���C��<@�=_Z��^k=J�W=�ǜ=�"*<�Z=_-�8�8�;:ӻd�z�/���=ʡ�;��༚���D��iY���o=#��=��<�ߌ=OiS�%Q������R<S]���x=�g=҄�=7��=V�=��&=]����t��#���|Ǽ�!�=�n�����V��,���E��;{����;.��=�G�<C��<���9�=�}�=�72=\N=�"2=,꼠�+�6��<���<�U�[�ּ��7���=�?X��=�N�����=�,�<�(q<Yח<>k=����;��^d)=�!��39��Rü�Q=W�;�=�VL�OI�=�ꈽ�e(�������;􉥽a�K=Z�8=��:�:xN�	S-�|��;��Ƙ�;L=���=���<F�|��<�{M=����h=�M���DC��0F�y��]�<*�^=6��=P�<��{<� �ٶ{=��o�=Z����9=�3/<�)�<���<�����
��FȽN�<{i�U4&�>)F<��l=9B�=���򭽚��<�'��<�O#�w�=y�k=r�=ѵ�<�S=�R=8����B�*M=��u�4=��K��>�=�cm=ɚ<�
�_���o<�U�ó�~�\e:<���;����ʇ����V�<[�=�/=��9=u�����=�o��<r=�r==�EK<�)��)V���@����=I`�;��+<���Ӱ�=�TE=͉7��Ż��<� �=�Y�=7��=D�	����&Z�b C��	|��?B=��&=]�9��������/���g�=&͕�Q�U=\�L=����Ŏ= ��V�E=��C��S���	߼y<<uy���+=E�=�ئ<�_=  �`%7=�V=:j=�-q�甅�z��<��G=�/N=�Iv=57ƺjv�����=�Բ<�%2����=O�<�2�kޑ<6�ǻ�p�� e��¶�=<F���o�=��.=ۖ�Lwļ���O-����s=%d?<�C<���?<���<ʻ��h*�<�ն<=��=�U=��}��@=GQ�=�S=\�~�$4����]�g�1�A=��<o\=>:�H��=�<���⊻iQҼ�z=�A�����<���<�3u�~�'<��a=/�;c��Ӎ'��.�<�6k=�6����1=\�m=.��=h"�*��=d�	=��#=pp<�G�<�r= ��<q�<���6:�!<6��}n�=� �� �㼜η=�蓽��6����<;��=ݨ�<-�<�.�=44a�Gf_=1o=���=�,�=�r�=�k�j���=8e�yC��e��խ�I��<��}����=�p���`q;^}m���<��=�tO��r�<ӽ�==��.(!�)K�އv�l��|=-U�=%f��㼢}�m,T=��:=�@�=3 =��Y��x=V",�v��)��\˓=��$<�ۿ<sɽ���=�[���i�=[@,�pr<��o=E �=�+H��p�=��&�"5
�A\��6%�X��`)�^fi=�B=ߢ<�?���SB���|��ث=�,�=��#=�&>�<�=sH<�p����O��J��g�=�=���<8i:��,�(�"�j��<�b��?��9[=r�=
�<%��K:��b�=.嵽ޡ�=�{�<j��?=%���1텽�Ň��{=�ـ<�=���=%0=]�	= �c�5�r="��0k������hټ��;J̟<�ϲ;��e������Y+��!"��i�9��x��<�E��EJ�=)x
=�h;�P[<^��;�Qr=���=}|��P�=$���U#=��Eu�=Qؤ=�����G<㚙<�a��[�H���^=�Gg�,$7��Z`=5��<�t`����+���*d���QȽÎ�<�`�=�<��8��K�=ݹ����=P��<cۍ��Zg<8f��b��с�u��=�!=ヽ�ߢ=-��=Y��<�m�j�(�8�=h�Ƚ��=`~��{k<3�d=.�<y1@�PK1SG�      PK                    " 0 FIN_seed_148_int_414_head_4/data/8FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ���=-���� �N�:�o�>�v]<�d�
�u�����{2>P�t�H�\>�a=��ܟ�=Kbn>&�>�S�>��r>�(�0���R�4����D�v{:���p�M�e�>�2x���8>�Ė���<ԋf�����z >#w�<qMJ�5����������>~�>�3���\�:��鐦=�>ʗ�=��!>��H=m:�.��>��H�>R>E���Q\6���s>2�*=�M>�����7���>�r��z]N�PKZ�[;      PK                    " 0 FIN_seed_148_int_414_head_4/data/9FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�H�9�S��~�k�
=PK"<T      PK                    #  FIN_seed_148_int_414_head_4/versionFB ZZZZZZZZZZZZZZZZZZZZZZZZZZZ3
PKўgU      PK                    2  FIN_seed_148_int_414_head_4/.data/serialization_idFB ZZZZZZZZZZZZZZZZZZZZZZZZZZ1134580559561873121713097790757992241736PKqe�,(   (   PK          a_��  �  $                 FIN_seed_148_int_414_head_4/data.pklPK          �=�      %             M  FIN_seed_148_int_414_head_4/byteorderPK          �z�      "             �  FIN_seed_148_int_414_head_4/data/0PK          �y      "             P  FIN_seed_148_int_414_head_4/data/1PK          (���      "             �&  FIN_seed_148_int_414_head_4/data/2PK          ����  0   0 "             P7  FIN_seed_148_int_414_head_4/data/3PK          ���w@   @   "             �70 FIN_seed_148_int_414_head_4/data/4PK          ��LB@   @   "             �80 FIN_seed_148_int_414_head_4/data/5PK          %[�?@   @   "             P90 FIN_seed_148_int_414_head_4/data/6PK          1SG�      "             :0 FIN_seed_148_int_414_head_4/data/7PK          Z�[;      "             �:1 FIN_seed_148_int_414_head_4/data/8PK          "<T      "             <1 FIN_seed_148_int_414_head_4/data/9PK          ўgU      #             �<1 FIN_seed_148_int_414_head_4/versionPK          qe�,(   (   2             =1 FIN_seed_148_int_414_head_4/.data/serialization_idPK,       -                       v      �=1     PK    .B1        PK      v  �=1   